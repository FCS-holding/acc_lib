------------------------------------------------------------------------
----
---- This file has been generated the 2020/07/30 - 18:15:51.
---- This file can be used with xilinx_sim tools.
---- This file is not synthesizable and does not target any FPGAs.
---- DRM HDK VERSION 4.2.1.0.
---- DRM VERSION 4.2.1.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinx_2016_05", key_method="rsa"
`protect key_block
iiLxHCp3GL0rA9HBzVe33iq4MJ6Hls0RRI62FxcC+YNHLSNO2y+b6Iq6si3R0k0+oPWUCgiCiHAc
6xOx2a3rfVYTmyoIlVU6hkLDblN0P7m+BUFFnjuNuPkmbYRtfrPiC2pEs3Y2tJaMputxVzlz5Aa5
xebzn6fZP9nSSyw/1IYl4TIbWFn24d2abuU6tWvA6EvfADyE6K7PC8q9ga3xPJNQha7argWcxmlw
i+wdI2yh9y5otlzF3y8LtBKbIm6Q2cOJW5NWhUsNCZxmuce3iMtVEsKXNTmRkwAdhSNSy3Q1BvF1
d8y1aSfw/FLg706NeTVpm8+Qy3yT6iyFF//UfQ==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
g8J04JpNRbCxk96h6O6lU0bmqOB1DaGb8uoHO7SbYmgZu6KPKVJCKd/dffJ7C5u9z/kQPX06D8CH
2ExM6yiwae+SoLhgrQaDSnTA//AOy3p2adDKQI+BPl9eAL0PAkBJLPmAdyoiigdfxaodHqeIkwBu
6wcoW3FsArfHM7ONtA1ayHE3m0jpoLPFK4u1y+zYYsELZ26LEOsEzTth1L1BDjJVrWkRLgBfxpPf
Qx4GdQenyHQd13s8tCqI3oX/G+R6Q3SZSJAwgozFh539RTFuiFFF7t00BW0e0cKCBkRQ9Y5t46yp
1omWLW+c3RXNNE79JhdSVLDye6K32i2EJZFAgQ==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2019_02", key_method="rsa"
`protect key_block
lNwIzHLQIspkjDSYJcobsMRBqh8h6T3l7g6gSOGZS8AzzW9RDaHmh4gG56Uywi2WO7WZaGbB9ibR
7IpU7ZEUn6GuP8Ru8+vz02bJz9X0i37A05yUm0153K0KYUnN9dZakE3LYoAOVqd5h3BF38K38ItY
YvHCdEeFgGYWyPeOvkGFlbD4AUlnnODN324OK//r9SHSkwz9ccywgo0Uak9rw/K58IV8ZJNOACOH
dgmL2qDK3H1wIfQbJKApiH6N6IqA6bXVFg25/B3UeY6JAgmy72BwID2okjU+xJ9DbESUeudZFGXI
NDjj/f2UCJz0rmAIpJa86QDIevugybu/sItrxA==

`protect encoding=(enctype="base64", line_length=76, bytes=856192)
`protect data_method="aes128-cbc"
`protect data_block
ZAROfCXswkZUspB0nZyH/in0D+okMmdAABS6AbGmOVV1zeJaVHjFSDYZnQhY6kw2vVVcNivtKElM
1awqAKO98uKWtkGQsK/628ZbPZiknBqAI0T/viyA8lvJ0donEN+khnP1lK7fXriCAaa2TqLfPT1x
b1R+3HJUrSPhnzR97BJFMf3V/3oAo8qWIJeGaoUqXzBFpdfrpuFQ6TDMnHt7uJSt3eEig2Ew3G3v
DhL3sNzCRA8PcpvzsM1ttw/a+jGhc/qZnxG+Tqbl1qhzQ+5hd+EKI0noYDY4JkJeqsO31rtsTLuh
l43IPK+13gdKW0dEUeduuB2b0+PhxY4bHVfrL5Kw9wHFdzGvvSTMR1cVSE+jIj0uLbTjJUNjhKj0
jIkhz/AiwpTsGx8L4/X29LiuSx0PHNrMJs9nNsJlg8yibZ1q+VSOILpHssFOTNecuyT+W+FEldDF
ek2wqhtgnyFN3mO1XheFe4438WuCTuwxIkxyMuxJY9tdBCew5jGi3i5rh9hwLVOYBtoRtYNonZnU
SMkRKseI5E10SZX6gLUtze1EsJVa3SIMdt9fuHcWXObf/n2X8p8Nfd+0Fv8jwSsxuVW5aZq0ILoI
0skNWOSgebIernxb6aiMgWq/+jzRc1Bn/p2nI5USh2u+OMHQdG0f6o2m0bwRz1YV+rmoluIx/Q2p
12uPkULhjp/Vz7+WVmbv5YIA+sFNj0fS/6/DJmeTWI0g5o9zdQQBYUXMnoEs18SuGOBVszA+7OAx
wGa3ypdygwh31TIIfo4njIeB0qz8DxQlgO9RxbDowcea8B8OTq6x0lsaygVsjkjy7eaHpehoozRl
KBkG7PN43pjtY2LwtjV0bpTLLC0k1SrVti0+yX12TbiW/IG6FDAUbgr/cED1r5ZmTno0C7EAnLE5
fG0okhSjkAUB37QBdtJosUsRRziCV9Sqzv43Wjf4PftZLDt0dHKwq568LPYOT81qRdLSqRw33Cp0
brkEhtRzXcuXFp/L7r4orZZF2U9loOzI7BfhJ8RnnL+Rog8nJkB+5Cpp58eMk9kJcJX1c98efnXC
rSYM7tfqSxHRqEcV2JHzB570vGoT74PVabXqcF5SDUENVdfCbEu8+FuIO0eXG3vdfjlCzz8XhPWE
e1ind3k108nde4H7wpvlXDrEPFWkE7xd1+RwOez6h5u8EivWotk1gyIwyOwB61cPtn+nifJc7X3r
n0gSV9XoSX5x4+APtjkzdzyoV3VOtBuQnpNoTarZrlqCQGlElKAAdOf/idW6n7EzMM9kADubkBxO
Evwk3qDbvawq1wJoOpR93fpPk2SwMO+18nzZECy3ig4UNBljZMRcnPz//RGnJUbw/7e1ANe4wezn
iPunSMZEQ4xU/eQ6OQaN7qt9n2cJcfzkcYhMmXzlJIjf+IAoDwekGHuooaILcEtxMjcUWNZ+y43X
EY6ZI8Sv/VN08WbM2ivurD1nfD106jMDm33yldKQd529NCXToEvp+LjaT4VA9ZpzW2X25LknfOjA
DEyTZ3UvW8iEq+SmE+8tINkxnCfvOoI58sOXey1k1pjQ+kZW8PRlZPfRjz+Z+7f34hMctzW95qZM
DX2dvzk/yVnzy9o6l6OeE4qYKGvDkNW7QJ+Hlg89SNqa5KL7Ft4lWa+2xrrS3JllQVGvLKEXgbS5
8pz8/EqZDcW2ov274JF0HpoPqP454E7XtubZRPS18zL2xAHvuUapwKlyMRNpUmzeRVPP2ne1kemK
Gh81KtEVl8pRd5eFIabIYGmXITkwWbjZPhwwtYrq5AhZZL4g81voq8XKhyG5A3J7vuzgBi1rNt5L
Jy8wHclXgkl3nSe0qVSLpL2gY/kmRWFYdG6zJZ+KXVAei8VvgyqOQl4lqKjynpgzK1X5cOCUIZ4K
EqUqbCKR/Etde/pjwK/8D+rw7Ydz7jnDss4WWu95165RZ9tN75+d1Wff3l+9fn9MZ6E1XFcWooAw
VhoBywsbrrzf4e1RoOGyyBrkWo0RaDalSDiWH4y2zYS611yiwbMPHMr1BTQXFhN07L4kJSmgikad
3JdfK0o7v7hGqBfKBIcdCbnUP+BYWbu4h+nj1smMfb6AvHWKzMYqhlxoFK1KwnOvpAfvYZGXHFaP
HDi4cVuXqR0YmTNsopb22Tm+De1Xqolr7/QTq2Hnj7ZwehcOTp+00sJPSaZ2AmNYG1u2IX0VGW//
QXiYMU3dVwbWdADWwLYkQJdRhl2O2YLLyAsvTk8LT4Nv2hRb92LEJA7sKLRRTNtUJHPC0KJ3vJuA
tN4SBLB+3dRNVEwqnjx41X35x2DPiSdDA1+fNgw2XusZKmxm7ttw9P73TN9XRgq6ACxo5KEZLS6k
THCDkFtQ7yUUiWXvJRTKYP9u8MTyOnhrJaODx8ft4wIUwTpIFIinT86hABxLiuzm4/sPn+3kWWWy
Q/RdvI3kAY5/C1L/FZBqchqLM0e9MJVI438+iSjxjQtFu17JtjRPaUO+lvbSVvCcABVjFZFz4DJ4
2l/xQtq2tltmy/fmpnAFKGtthtXZBA7YFzCwE9dY8D/9QyPw2vHSvB1POOz2PKC51hZNkt7LNM3l
g25y7R/PYljLOgtoz8fWKMOXumiL8StyX9rP/ehY74PkzKhni77eyHonSNLn4DkonF8DRXdwVl2v
aVdJuH8aH9qPHrJqz/gnwM43nfWAeIGqwg8CP3TBjLC6ys0c6IE5XWj/5fEE8ibbS2BgbYHBT/TY
KsGP23sxFgNJWJSLcTujT73f0qxmgEvXEcofMBJrdHNDrXqGANsugkPWosrYWrhgTpgMMOijzlOm
BRBliyFl+vzVd4PhgkJRvRN91rKe5QuR4hTzS75FlM+/fBXuVQDnbHHJnEtusBGETYX/WHSlcPc7
ghAO1+jb+tfqToJrtmGQcPFpNWTOIMtB26ps+OizmOH+gzpODO8oXe+e0WXvB6m1UQwKu0qeu2pN
zGuE6i0FRh/KVyZsyHE7ZNGan4TTxmN+siY6XvRIWpnSqLsUnb6ucnto8VGE+h15BQ8Py1tAbc4U
9gzlBjLaHN/IE2Btegwk2W3HULzt4aN3dGaYlI1dzDbZr4GBils0keGCc1BkzemNuykTjXeV0fQd
NNEJJKSn3maaZFQBhHhgl3uTCYB6gkLKLbrLkIpw8WUfqDr3ixEMBXMjygyiI/4IQ11So8jr8eUJ
QQ8jdL4p2l65OrW+1t8xYAlPHPKhAWlqyyWlpy+1jl9OikfudLt0xrzxpYTtKdAPP0pp/z4b/vih
/Vadwm1tOSn7SGR7TM17EcdHIFtGXzwxGqrZ/iNNgrY79SevKXS/L8b5ekaPTp5iLZoML4R2himX
G9Scohs8/xwyIf7VdgFTzXxmSW5cEY4//qYNdYjq/Lo5e/Ju+z9U9StROL9WqPxhlVfGIma8c/NK
gpm+vsQYzPq3scJ06cUWQkNT1ctDt50BupdAUpfQtKkiKsVRVEXawnbvI5vs4rf/pg/0SUrZ1trp
O88KKUEOxKkL7qKVBp9z7IOnmX0Ejo9ykYB91/1LcrwFiD4SQcRzTIxokjRJs29kTBjAsiNNr1sm
qyyYYNXdV8phqSiQ6t1EXsDl0KXOOVAipwIFrgBpNvvXru0s72m3hXhMreq0gfuU0rgkZqW1yJas
j9InKt6KhVHOJ6ciZh+i5gXMafS7xXDjzXD4MIGm7gu53CdHV8qQAn9Zolk1aA2rTEoJ3qM28Alx
mTqRCvj/hvUuOU32/qAhoC8I0+9XBANse4InDBQXjKzgD8Q6zhyKH8hZirlU3U47WXaiB5lqRqm5
BuuJmds67fTsNe1lrKRfvXapIrp/SXG+HLSmmVdIaEfICZWcmhg1ziqJ6Pb1eVx4P0R24oySXjMy
Wdr9N/i4AfkuiEZOjof9GrtCA9OhLoD+HnKxmFuCsaE5q+kkoBIA7sntsHn+Fp7w3kAz+4h3vxNt
xPBkTnv1pN0e7bMcuD0W+jqOC7+ipzrXvEsXxykqUc/i96t45YYI/V5wsc6nJ9YlF1utGBZXMVre
3Zw4wDzRnyaKR4+8JrrBPC6N/CC6Y1gKPwziMnJVOZ43aScU6mXTSBgYALFpoXP9I0VMksv3W1he
2H8nODoEUzLrk/oaP5SaMYtjKCHalaT0eezcHibgJhBWMrdBvG8qfGKppJj0pPkzWgPX6vum8+VP
CJaMg0a8reXxVmIn07uGlOmdcrsq5doDYyiEmr8eyE0tbhZuL8VvNBdOGwHjZL92L6eQ+hpyEt93
9g2X0SEczqg6rZw+wiEY5CBF97xUbA67u4p60mGdParTv875j2FP7UsYKA/9irzL3rOhzz2J70XQ
IQOfdOBfCVRF/pbr9ROFvtvXzyaDrxHb7aV9lEafuvIjf9WZaIOWLQC6YEQjDArBTqlbISiJk6aj
xXtimhSRxiaXYYfUWAuo1rzB4hPHN5XXEZdwkVGQgZCyR/kI8rwgVkShS+Gct0ktk2y81lihHtQ8
w/nGfGXm8FPxuHBqnKLhL62/llsVDh7O63SdXfWSVQAx7ONia564wQIXHLrDxRK7oxNtzJ7TdABE
P4ANxikH6MHEME9uB0RuShMVC8Tsytix7sCblrsUjuXdFaTdF1VZzqNdfh0ipHFDaT59Ed5Am2rN
AmKvXnHKWD8ME7JgQkWNYIHbIqddJEsZDvwrFej0XjzWb5t8mMtVCBJPq8G2pxU9GVOBAafOVsUM
OT4ZxiivtpXKVNq7BesdTGv1VJs1cyTZs9PT31SupcqFf8Pdr7yA+AY3jNyaNPTft8vp/9m1RP68
tMTWyv3kkYbnTmiLEb0o+sRJvcNbkBu7zMBcwqOYWwKLiXP0tlyNAj6gy+rLmWsJ/dG0y6JGmUtw
uWxmwKSI10cq1rMckSY/yK6NQg5ScmZrRXR8yDStC+tPXnFmtvNnZTI2mQEDxKi0jymlAGcUT1LE
bU0RqlslGd4QAu6hNTv3TK4kfNftk3AGGJHMZzfefzW4KoK2l4LMrg2D1pQohGt1Yqy3ZccFYeOs
QQwDt8rzmQ8CBoDsSXFbzUIb9qvyA34x8HW79yl2fu2dJw3fnki7BYIwVRjr3RpediN+HMkJKNlx
4x6eHwFId7EMt8R+bAmXYQ2Rrv0clm20IXMM7Zjc2Y6OZgjsKYo+e6bMfekl6UImsWdaeJ6495Zl
6+tnbYX0svabiMKY1tfSYW/+EKUK+K0FbVvJWafD1NCucyg5VZ19SP12Hcj8t6bZsu9QNzaZ8XcP
zAHDOxKGRZZNRbRDVVk3zVAgSCWy1dBrIA7CH09CWNECDNYdKjmR9FE05OxW5n5lbvIi3jYUzYNe
t2f95MgEcDd200dTavIjJz3pZloXtWw8hyiI6rTUOwPiaJYSrjgn/Ql+sVQpcfKIJcAtFIuUkrTV
f+/gsGk7KGVlRtoile42jA1Ua8TzBIsZ4F85DHbPFaqSKc2noR4fM2Kd6WMeJgAs11ES/5uaBayM
fwZ0TWZnclDYNXXSvxrSTspnigb0IP2o74jku50YZRsYd+BDZSfzzngldZ4DOBqEn5kgzL0cHDZc
caa4PcFf0E06xrGsaK2yLKt5lxzIIFwggr+v2d8SSbIFv6hRPi7QvPBRiJKRb93kyBB3Pz8dVDDh
NIJKs4DLL6ha3GMxIjV3x/q5GQ+OH61tfjIBrxY7IJGg8JfztOfEmiYcEbxKBTM1dX3zn6zrLTDv
6aHrOiZXhUuDaeOAitfB4tApBCG41BBeYMVYbss60r5GrBmOL9kSJpMytj5uw9bWjFRBjC3cRLaH
8Sox5h/raDPx5l+Afo0Idh54c3UIyzaaiZM/iQdkz9GdWQc0aKipj3+cVXrIye5ZvyL4GyNtgUS+
FzHfbwOTPIDB30F2AVYFJUeAHE3rTBWZCqgEZAmZiAnnOc7p6pfW+3xe/lzxezwud++XHGJZ9TkL
+E+nN9/7wsMF78R+OkyEbdnVjcCCDzoocUJXBG8y6h9k4Vv9C8TcWIVNjPud87OaXob7AzaBmaHa
p4thCkoh5xtpAOOn04QcU4GMsqaCyrAQx6hgx8Ki6xFlTZTX4JLYqNzg+Ob2ZTchJkd63YzKh++W
B/BH6O0J5u+Wbo0GZ5ZUHPLjQN+cD/8KQPYhPLyGXdPPoHpUPGgyp3lPqcs28K0DOpkiIOqnKuzr
Bbp110LH6dO1SzXGClFOLMDBYo3dA74m+kGycs1kRheT/hlzpyR+o1R6phGRPWniFhaE3LFQBud1
DMhDKYEYDJq38i72mj+CT2kOOru4jlC2ByLZgtmKDTkiqGwQdR/7kdvz3DzS6bWlK0N1tL3IZEMy
gtT2keILA52kxJBIYbat3qPvrcfEX+kLutGczoQnlVB0o9vYlO81ZWMcFE7BJ1dozL5VckqixxIk
zfWR6NPhQJJUL+Kc/s7aDpQ6SVKiQk6VQ6yZQqaAZND/1DMs2Grp75ekXhXlMdUTYzA1O9FzP7kJ
lWASHF0lXaleaqGje4efvErpEKyV6DO7H8/dPhGPhfGxIkbeK0rEpnu8B1kP35NF7Tl/9SilvlPj
iIXvA9I6/EkbdWdEeMi95muC3rSMOoc33n7jWviA1VOf5sjFXlJ3JMrJHQLUIxpo0KBCY/UDM4KT
2w1n0lGbjA0B4Qb72mNyaEM8/ZKA1koJ76P8FQHyIJiosScPVZs3fvyFM4FsAkls4wJGJJqOSrvA
S+GXZleJeoSNSi4+ML1uSju6BXQxT9DmV7kn+AokLd6Xy+z3okckpPDfkDOTQsnqdMIQFVefAfYi
1L66O04THDmjZrfIcaJkQqWDwFrXiqvNJ0imF4+Xgd6nrVzeyMxrBlENAk0DI9s+IuY5ZW0qUOC2
ot/gsyQe7VxdfF4TOMzrIZTgS7PRE6fRFDiv/M+FBFyEtmm7yfJg9YN1QnXQZ1gYg4zpehWgWq+c
ECXvsM2Y2OqJM2MD6mWdh+f1WHkOxn0BimqePtTBcnS4giyERei1gdmwSbzvlfOhEXVGdm/7rE95
VAR3gDKHeR1bDswvrb/RvYaJMPkGR55nxLpJufJ43NGADTTxINwxXaqn9wzP29KZOlW9YkKLYsCp
GPd+wOFLTO3ej9ai/qcgwRh7ZVtmtrxLY9zbOywdZoQezygDtQZ3OWRDZ5A1jL1WrsHffjLRVIB2
4zHPKmhOEm8XthZRJzXTn8i/aTcNnb9mqniKpwQsGFrSdc/f4aYtH69x9lQQ97ZOg4l9PRIyAi0+
Yo/dsVCH8cUiDK/R4Q9xmbIn8HLPHRvicWumBx/RX0VuoIf/IoXHtx44uHIYV91pNwgaGp7yzVgc
Vox22Z46yZGuBaglWwS+ZAr4rM83/IPR6kQfifnVzDvwGHJalIv9G3fagzkWN+PkdBSZ7dp1OBug
oefEI2bZ7sin6XDRCPNNRfyWt4mt8OmoK5f9bO+URsaPEmOhlDxsKXyZ4jUxD1Lw4VF4ejhEOYmi
IVAlAcSFLlVu7GmrWr1bsmPnBu+ikATIi2K9ft3tOVcaBVkHnlsPUN7hVWJmU/tGi48hDxWjK7Xq
H7D9nwpQmhBpBDHfLety8gvGQus8r6pI5RZ6kxsrLZ4C5E9uoVjdCyFIx+ToYdKuOdBipAtXuKly
5c6dCGjO0hmsWaqWEL2s4khel6Vbj2hD50wCZ197RPAgFnxr2vbTWKvxL9MQFVAZ/qxSOD/LCfU3
t2H+8LvIwAufQgqIfyStpfsnKGJLaILGHxEoY61fdLAVyrtTWiuxxkQa4ARXQtCNdKSUMf2g4tJp
xQUse2ayWrYnuOhPwt9W3RePezmslOL78DuxLEVk/symO3TxeB24MV17m5wMakZDQfQIfUb+pvsR
C3vDV23c04UFXCIOKvp5OjYkmyGfoOfyT73fc974liTlR0aFwLKjko6CdYk1z7QYY2s590lIrC8A
MMLCPCGAcNfM2b/fTlMYGT+fNKBGySK3ljYj1ie/35tZOawOoJ9moz6Db80G9SZQoefoak1yMJpP
gyR8IYV7i5wqtCh1k+pCFK0Ty483PsCBK1Y1iGRzrxhT1iaxtAef873Zw7RhZDpANiKZgQr9ZI04
pIcZOZ2PopOilAysq00Ef7M/01xGFfNoomVQErVVXZ7mO+JAiX5oNAhY905m3jXnFlKzwH9/zcZP
HlJ0xx7YLierQnGX3mqkt5JDnCft9RNS78aRTKc4/jwDmvLHR0ekkQaqm9hg48Ayk+kGDfkf3TTs
Gx2hblYaeIoALnkSZGgFlwlJcPoFayKf7A6LcbdAW7pMAku6CUfsjJkqzWX12mrczjOdRh8g0UVY
jGxlu25Xw1E5PjMAIkbdmzYmoSE1EqBklm1I4iF8brwKe0Rw7N8v911f9l9iM39GmOKStfxKjdSI
COnpqpqK9XL7X0m94cTa5fiAZx8oZ9Kfk18PUTkDT0KT2VPZlvdPIZGKzETI2JSclSSrOgtneowk
3REiaqFOu+nBHsBmY6d4H9R73GOGf41sMLcIPbusa9XK8dW24P8KqxrkOjtkH6G0p1MOgKP3ZBhM
T4j5UK7NAMJzF5WG4RemV9RLs6QIGUavvRC/1V6YoY7Eems6XhSX+KZrIzM9ANBemlOXVJN7JP3q
pKub9cu92kJiQkQf7G34RAmXKq39W9ayHgproo5s5djHec+tpgTY/NBMCLJlWI2QWPlQ0gerU14P
iUw32948alHDnxEN3Ntonm9E8LKewMvHOxj7Rh7DlyJUEPE4bXQzpxYN8WqdXKw7aUZwGBQWJ/jf
HfuzFMi/QaG83L5l95OUCvWsWGse3vFpL/3Bn5YTOdB3YjWjXNmRnX/WpT0Wft0XtSrYoEfAT8KS
rMjDkFOTvWxd+VwwyvCgX0TbZsz4aZVWiikptmV/v01Ev1IqEpT2Zyn1IQOnnLWG+Xx/0XM0yv6D
7pkvn8WYNb1bXOqv1/gqLw+C0tqlRkQstSzdMbKrEGXQPKFAHnKN5vHvidieD+dSlwzJQd35hBaD
N/B3zv9Y6Yb0MY/4q/I3G1uTzxrrzbp7PigQVrtCT7RD3NUWXU4ThaROR9lz/Rrh68U9Cn0W8Huc
PpeHeN/DITyQieewXTVZ5YPLGtMV3b1EvABy0Feq/hu/3uJd3K7ON5f4OBAdJZw2EkOUK2sAKByX
prLfnxqNm3z+tTPHc1/pwP3sfEUDQXww3lzVBXCs/ctrqMdloQLzwRxuOOrUXonwLOsf7g1DQLqC
5XQcl7EdDaR23a3iQ9a0jy/rZmkIY1rusTsb0CECRoV2sRAe+ulCWbWkn/fsbjW1hauWimpvIXVI
OV6oebOrv0xmLrrU7flGJBvMnJhmM61dAUo4MTRrLwI/HYYJUdcQPua+dZMnv8DYY+9GdmEq3VbW
WSoG1nodCgs/LPVLht6QITyY0IR4uapAum7T09/2dP3idyBJZrH4Xq5PFesIFRgdGUkJf86SPxIv
jycrrd1uPW1cpE3EIt6RP5P+246EkEBqsFYNFOUGHeWipt8VuarRzyth32FpD4xWuz1KITgJY1pr
lvN1zZiJeUMhWgCgwhimhl1D7Tye2QaoK63TlbL/lZ8jrr+I5PPAOJyPbmQlmQk7iTj52t+oCxLn
B+93JxZvGexCCsWoPbJCiXH0p4p+1TD9EAEwK1Lb7Kb206fz2SrTXMTiBAnLUprw1P/gn9PWF/1i
RQypZAJxi89gQRAIDKUsoJan6IEApfxiSQfzzGJiQrIcmWiVXQthV+wwyddjsdox8LWApeonF814
bre4rdssQ7ug/VRZYeht/TNIcAXya0OMm8rOIuPCb4mDn8FjANWWt4BfdvI83z8zQDtvxkfedI96
SSad24bIspoHzjtBat/UnIZs6kgvLn0zm3jPVuj+qQ2fIOEzktdnU9i/83ROWiZ3Z6eoEr884b+S
7+xH3SH91y5pgCfYiJWV/2rwkbPr8svF+TsUseE/ndfxOSuGhQLMG/L5tZ7QzRZKRVx21oOGj4n3
LYeGjaE9/rRxpEROHaSyxMusIkE1Np5FnwAlREk6m23LLqSJbWDMmARHVSlV5GyEFexmauhZRLJB
HLKGCU1+KzyEXWCH+u1k0OSfDkomSxJyeJ8cfoveH3s/7O2FvdqAYzmAyCPWp61pIt8lTZ3VwFU4
Bk+PfA9JWMyoKje9WhtUNnSBUlB5jdQ8O+o3s5BmQ4lsm+crNfHnN6gFrIKwMYZbwJZ/xlJPRhCW
oz0XWWhjP5hvuY/PXi8FM4YMJ97aC92VKYL9C0OGuLI2zVhU0OgMsmBGIJ6/akbZT18zYMu3c/3T
/cS3DQiosdkpUD9uONwWSxb0ujkhwlURMoj8CNVEgFYOrE+/ZrKRkQVLfez/tiKv9lUw5ye+KRPl
kQkvBI+Ko/wnQjhZ6nbm9yVfcoa55gBaiA6Tj+qW6Yj0iwlZ6aesWosiB7N4O3OL3SJ5zDdeZ3sL
/1Gln95bgn9C7009WKjYT5Tzuwwy/uJBXUKEBF8/sVwS6ixiEFPZ3KMcLprJ8qd6yLwKC5oMq2EP
Jt2QXHLvHMueGIPNCFUuv7RXUDfdlTGCGVu286SbfPmcbEP7Jd+rvvwl8Jr1Oam6vYkSQxyp9HLd
E34dUKwG+kDQV3kQvK92JEiRCiDa4I2Qq/WrUST2xm+J3bZ7ifUmXSzExhU6SYd6GYJX+AtRgxsG
Dgvee6SDYPhPgZiS/HjaAcSgsjJEWnSRVoTLzoZIt+v+9oLcLUPkS8Ruf+rD9irTWJVTgjYNfrA7
VAkRiQG2T4xOVKM62Cfr0iQXI5go1AQ+7Qm3plklXqIWHsro43x7bzO8XzvJvvCGxYq1TNUDExiX
69nKO1UIn6v6jUbNXIhL98frkAe7wIJH1cGhbs7BqbrM/eaciT4vd2MztnyyKU0lTWFk/JU1GArh
Hr1iIh7CZzuEOqHLqukoXVTWjakAy717Et1QerTTu27sv3UAMbx9QW53EVFaWBl07UroQu+KRPnz
R9Wr7sLEajEL+BtF4Y4Y4IDCq32W5Pwoxdr8uxSUr1yRizHASWu1/tIdZoAtDb9m3DgGisZ+nqUc
m6BHVqp3P03YDMHFF8P9bQDqBgD5wyDYFspAggQWNd/LnRoqYsT4spaZPG9gw2jys+9E6f2o6K9R
St6kqsot3IrSql8iz2dYf0bx40YLa2ysmcE0Z+Hw45IB6bRCTaNkBMQCmSwUbJiLzqRfza9C0PHK
4QWhrekQ2ZTZ/b/jr3O4VERJ1l7kYCCBooJy8RLVhvO8REbLIYKZ0MFCl8qQUdTxpG1IsBwxmaNI
5W+3nJkB7rHLvNZwTe2Y0dDpClGBSov9GOEtYtejGFDoHjIHEVpovDlyXBwJq94YuuNlJM/lUYAS
7XVZBVG5EH4uAxtG69effCf/E5Ox7P7lNCPI46iTT76epg+S6IagHL/Ue1dxxJ7zm82Z7ToVmYE8
2Iy6mtzuK9HW5javmS6zDxTmfxLlFDjMbloVgZCWjF2Gn2/RH1m3PqgWGfiiz8drJbQCxYjT/HmU
fcu8K98L/1mkMkaExaiSWpr9S5sRRcjomhJbA+B3gelh/q2iY0tEGRIaE/gCwveEYy19OayxwdeZ
2gzJmwcq5TcntjmAUuyPhwHWpUS7VrKdz2I/r3D5VEe58qkO0gWpOMLrF1ounqosH7jrCqO25YZs
qbLylefjEYjuNGOep5Uaz2eWNBAAAJvytCCPITgs1NanfH9Dg4FrnKbaeaM2VZ+a4XpnREAQyHqr
zl9Q9TzYLagClL0uJmf2MuySfRmJnKFZmhHQc59iUc3t18iaq3W+TMNIl17dEDjDyzFYuHmH1l9q
GMsQWux7HOpZ/yG2Ig78Nk0CWd5/QFQ3ewRIeLBa6gjIeTRm7MUYWQCqeu1N80p5wQ51ahhV/VGk
Ux8Sh+iiq2AxrEmjk+2S3ASsgRSq13Vn97A40wEaRstDkpCn0i2edcnEwpQsAmtR4XoWDTjyuth3
LGAXrTgvvjNQb9H3lFxxxCQiA9405ieJFE7yCux02HHqLtuqFeEuX0EHBWvSmI+HVOgpwlUSV0AX
MOCTCYmV+PlSf7MDs4mhPurdECuts0ur5MKSqH1UfTDb9j1XqqNPFOu9kjq4KoXIPWHtOV+A1Pkl
mBjFVAvFNeJxCSEOQzfExqkaP4IAhVyQ+k25wTZIox6sP+Iq1WQN2jHxM9cAWTZEtNoHo34jU1Da
9n89iyoltmqhauguM4YA4mz2AKA2A0s5j0sZE3t643Y/sOixExIYl/8+/TumXyS+4HJahVj3URgm
pKvvoSyGCjA/lr/xii0rfHkI4a+2SwHkDULwkf9AyFuUpSio/5Imb/Kf7HaOK+Pv7/FseF8SiwW6
nNOVuuO4HKtxHttk5EeLUQ9jUpgkQjXHugAkcyzRraeBl0fPe3wSlD2ZPkUOWOW5UCbL20mrNscJ
7eu38XWpAOOdviAVz+ZiZmjyGm7Vha+Bg4l+eU0zItiAR1K8+ISYMdmrE2R1XNTV/LCpnFGqHjAY
DB0ybL0hRs5NbUnk9/+HNBmC+Yv08AVnFYDotm8PhvaAdjeV8Qhk6GRnjdTnlIlAypJy7J3MHnNO
zZ+K1kkwucC8zxwH1HZbPCevoza4S36qCj3ZMt3gOMXzj82GkZwJ+Ia90OBz85Goim3uTU7Z98np
uIYmy+I+GMPW7UrEg5l87vS609uWdNbrr/TMWQQDtk5tUV90dQUYSbaRMNujpENSyB7ADGsA5pxp
JDSC3+/iiw4pu6w4m1t4zuZDxjZUNJENaa0x2IXmGOYITF/7B70BhM4X1TkMMm4KpnuSR9jNiz1u
y9t9cWAqVfqPPNDyNGeXN5hdX5F2yEw/YCxCqcwNQZVzOJq0rmS5GiSRs+Q2VT4NUumDMZoL8imc
dth/ggwLeu2j3tTKgjms1HTbbLbgHwxwHrmUgkml2SWj2Tr3nWK/gRJ2azVH3oXBGDGmy9AAKx0G
O9PNy21LfAQQyqEaRX7WQiAvSe2I7nuCSP87NDn06yHh2o8JnUGxpV8cQ4ybW3z65EWemb37zZqM
EmuyKBdMmI9+sxMUHbl8LiYiuXwWba+GRs7CrU5gZrLbXJQ94plWR7KGkXrHg1Zj7HjgxuNJC4l/
zN7eJPpmygzvli4JSoLC161qwhpvJhFGsBURWbUQ+JtKPPTqksQe0P/EsGPCJ91J+5/MY7xynnKR
yaKwoRxNZAVbW/2n55MA+tLM5iwfNSkH5mBu1NMMpRnWivVVsfQeoMdhsHPtTeUwnfJWaZTzrcc+
j49/l+XN1RO+1BLXKQzVHLeU0esmgBUxvnxIu8qJN4uVEnK0Vg3sz6WNAQeSgdfz7E8AsWMkzCK0
IOqkcr51/lifgmYedCL46ze1yb0T65wH0fN3VpxuSNmF+b8X8yOP7xZJvYxGNBD0fSKvsSKIXsct
RFbE/wdJtELE8L0bIV5x2VlSKnS9VTflU72OJRuxqQaQiRJTB39/yPdZ+Stmy5T0V2/NF7nlvE+6
ZxCkEGLqEB9VAMUW2L5DiyVw6RE3Px4VuoHlBmC4AZ83nML0vT0Znw2JwpSnWJrBls01WXCVQGf1
enNvJ9kNwwJL/oaWf9r8LjBqFpo6AFxzLm6JXIIKB8HanUhHjCdK+nAsUVyfnTsRegztL/fJW9vB
P1i7VDTrCrzlbKH2fUQ+M/TpHYwoM39lkLN6Spd8/R+c2n/DZxgRhoyCHK8RdaceX7iSjGaDPEvx
MiaNxpqYdquwiyyHVIaZUGpPJc04eJrY3zpZ3GHtptMU2UvslU1jjjYHbGOO954y0QWoqHjIiENv
EciwJaEqjqp6jpWHeBIUN6E5iNn294tAFkyMZadelC1gTNoYEk6lQcQjHtsGkLACWfPcVHuItYIQ
n3T1e/mM0FGB0BHGP5h/Taxgy9vDg8maWLvp5/rCYbGsCX9j+4hOgciNyIO2JHBhik9r8EUvsA2U
TNRc/cqIDeGR9shi3BTUu9WAeR5U1aM4R3hJecRR0Uwrw3f4ZQxvvNJ5XNfckjED7dO+4ap1fXz+
HHr3QBIsp2NHYWavna8n6rRMTxObqFqZDeQuoZjCG1dXZrtXjwLFpjQto5cXCsoRj08ohalhDKPS
AKpWMTvF/1TzxRvjfQhr/MXn7LiEIrEgBuKdIP98Kt2CALrIS7QrD8f5V/cBcwexYH26igJphDH6
MonLPzDFsU/ifkRx/Il2pmb4AfPafLUccjlCgR1KVRtbJhos3v9kpRUFJGiHOL0plamH/y4pyxoF
QnD2UkcNi2tlLd3pbkYFo6XDGQ6oYSc3DdRiDSc0QLasIJIPsL/bCEQyLxeMDG5eTtAgNTh8ykZT
gPoF7+yb/+X9j5wfGo8Mls9zvEJge/ZvwxzB7c1v/X1s31RDdF313r99fklFR0suN3qZkiefiib0
59CNpleBVs38hoSrKTkKvD+r1v+H66quHMA03nGjUGfo7PctyZJr0cIL2TxRuiJe7t8Y3FUedenc
bcIG3OQNFO01RhDuVSaSMRvuz2Pe+xFHj22JtKweyAWx6eLPSgLeW9mh0z0v7zGgTCkh8Q0t5QhN
X4uGnIqwzbhi605HFT8YqH4MDHQXqMQ7IHi3OSjrmIfnQMvYnJgSPscy6w7QKTmJdJxFU/7hdxic
51+YVefwy1/ZkI4KgHtRqJgTHQJQXuU9fpuG05xsLsnMSlZsRu/GgimaZSyBAq7NXNPWvjbZWoc5
0aUcRBFVXgFtKGgHbwvsbtHcHYEkAmhjG1SnazLPomdXu0YVuAJPNNbZ9+c6LkiRIYCUsXsa9jm7
PVIHmwpZl0XcScJYZhzUi1oSObO4hZTe0DDx7Z2Yetp6z0C/47crI54bWo0OgDKTcnpeJgWJH+Vc
6bIjOWP83hm0qU9paSz+BE+QcHJlN6UW9Tw0YgLlzFfvvvJj+96SrxuHrl+vTp+DEnL+ot4/EVz4
meANRtXXLyt3V6T1g5SKrw32OY+1Fmy8jRsG8K+sG76C12g1X1x3ehIRZ7cyyXbA/LxvK/ECg6Nd
KLm1yhPX2DHcwzB/cTEg+z8TVImyGD1+xixoBY5zQAiO6GLthpPPqqZbs8G6yfXEfhnapdPAN46Q
EgRRRyBfUJdDlqUgTmDLYBbPVLoEMDBmsleWc3x46+wedVv+eEGi5ePDHz/KLGDvMaAY8uvgYHQL
YgGN0zwCePu6d0M7Q+AK6Ftrj60mOBR3SjAKmfBs9ybdrylg96/M45Kg89sLnM/QnKmcXNzWkh2g
M9pvN9GsOykA2Ar65Aduu69cFncmPlWbk9+F8zoL4BKiXxQFZTAMNyK0j90zBO/BrsGehVs9YDiy
FsU4tGLhgF3jPzuZ+wdWbVLxJML8zPtPV2os15dx0l/RDPUTJ5nrRqBrW4gjxUrxwyA3q2/7f+Ck
V18Pj3Vd5UPfLRPrrAvD0r333GCKkH/KcRu2N0bqWMz2X5LAIVMPopH6RR5ghzw9tUz6lcwYm+YM
0CkVpVuLVeY89+zd/rx32WdFkeD1m2eRqN09MWiPgOpOmKm4G+XYFG0JS8W88Zx/lH0/bel4pDAg
vY5M0eFkjDc+68cPHj4l/XSSzoYHoGfQnvhcNRlzv1KUYUwjxs6PzjfipaHv+a5RZc8wHetsUhg/
eWSd5fwr+HG0mPpw6wmahzKo1CRkk0NEqjSc1/j2Lw7rYgemjNOi5fdsaV4Ea80OYQR4jAbjJkFC
2xGHmD5/xsDuoEHAUVmL919C1FN5Gi3Bq4TUe7xGxzh1rJqt+K7wYQJUA5eW0oFRUGDhB+1RRdUZ
HrqLhFbQxuTNgF1COm3jZu0IthmIFkJv1aWg8doWlIhJaOrXxzaVlT8ddVtB9YnS689n+zozBQXy
JhwQ+4ws4wx8894cGjaAnJkcERuI4zA1nD1yFszh8orBvOg6/vZWv937VfWmoyM9WC/Icp1Q+y8q
sgUbK5J6KFOWg3sJYTO0cWV5ojbR9Oq49pSGwAXslw5O+DG+9QR2mKnAbqrPUruUX2DBKLvcgPZu
9+O6V6dU1QcRXSyyW/ptC4BxMqxUxEefdhe4KJJQDkufb77z6AExfH1ySoB04QwBCToM/FFx3tV+
xkyMYHGCBS5Lvqzwpt6oU7k9K6Bgc4MAXVUPFeNBaxbY0vWz0VYOPc4e27XuWExaWLSAdZf8S3gh
hutLA5LvYmRbTtedadv9bSK+z1AOQ9DTZK/OyTby4kGHinDaFQet96nA88O3rZaDKPo9T6B26rEP
1jPI1bE9YSXqwpa5WPKUsWLaLnlPhg4NSVGcxt69FsRlU3xxxaXMzIIu0c4MBhZqJ/lwO4P6q1TG
46jsl5oZz+8bBU9HglvprhR11mjm5hQ+o5+FUarbGsfH4AT+gDAdVCP8oFFb80Lj3jNnMRhWpFga
naDREfAuCERTPiRSgumVd1tSg9vLpAl9BRs+ULXDz33UKV7Aw5uxpvz6b4o4wQUD0bL2xHcVrL32
edeEx4W46qX9SBbAyOhGTIgKHYuKSnrDKN+8S0gJ9I21nGNjx50pjif7RDAqiBTRt1CCwlNuP39/
znFZCF7u4ikgW27MFU/nGKKL4Oy+cn47V2oESuo6Mba4X1cFqS625q+Xn0m2vWGESiOmg+OAgnna
9EuPaLrKADsNVqlPldY0LxIwdef8Rcq6eWX7jVkApNh0Zww2gHttA9eIau63nxozGAjvLZcaDn1M
CftrVTg2r7JNBehi3HPryI+gx/VLwSfncK39ALvDkBd9guKBQZ+4u4ZylCmpPPJkGDO27ZqmyvLS
K3UuYHtxyTdn5Kyz0ob/pnt/pKoDViv3l0hmu+ed4NBpertFj8MJvQncXjW9XdUYDaaJkhyq7PdX
tWjtKy0tiPua9oRZAnb7YpRtRua8TZeIGaRD3R6uJllhKcZPzomb28CzCG8o8jQo0Qw/ZfD4k1Yn
SsP1l+iYuEO3osDsy9bV9hwP4Ds3BFHh6i6/2J+gHtwBnN3m+9lZlXOESWn3h09RDiz/R0x1Mg8w
cD4byQzz0KiJsZDpbZJVxBwzUpGZw9ardHFcxX19/XcFRHw5Mf4BX8gMx1rnZMmUfkHdEB8gBvTR
fmFjFNMKaOGFs/wg2xolZN+YV27J03jzQJ7N9jE4FwMWws67zIObiss0+CAY5bWbeiGxWGUQKhGX
iXedrEfGkuBR5HiJHlhrMPqhkIWqIUA2127/j+vfYurn0YypwoCBJ8OPHVH2LPXIy8jw2Vwljx3K
kc3IVnIyKPab0NqrQIT1T39h4aZQ7T/Suo/44+hMbh7mq20lVVQ3K4Dd1yEniUY4L8U2jzbj3FEr
3X4T2/77WK0bqck9MDIqj0roHStRwp5XD3U12HrTiTLzvNPuos8vv2L8y4dvW008gyC/E6xG4w3r
vFWlFSfqxd5gl3yLi4fI7Gf//OUMVKee6AupVjEzdCXnlEW75LSQs5KJkgh6nitDYPd2LXdBPJFQ
bGcfvdMlQ4QRpAsP5aPeRXeLJGkJduwi/98CXQSRZF2949Tq2XIJhgDHVKtBQsR/nq0g4HjZvdAh
NEXwif01y5oLvJabOqjZZ080ZBKBCkSXCy5mWuHGiKn4ulQ4LCaVQTeTFsYDfv5vKvGaWaxUjTXb
GUHRQhiUqnCiCBDDqumWEt+gRxdCHFPxHcVVRXAJbKGEG3gR7AeYFEBpP1dDsNXx0VMm0qKTTPVH
aX3rR2V5jGWx18fSl6yMtsO4UM5dQ/bYC8T2FqfaRwfGe0gNKR5y16rkPyyF1ngWc/b6H7fNIF5p
TZzAAscDzqjQMfhPktuyxwgyAri7kqjGxH8yyY+hqc9CJvJWxhH7t4DVOeS9N7BbWwcu7G/fp67v
Qt4G6SqeM/zGs2K5WMT+9nTVbx5XZOZALJywC0/bj15P0U7mV+PQfA57Im63YXXeY1F8gRspowWq
Bw4I0m+y3ar80jrL61gViB+DzUuV2Ar3oc3UcLtb8Myb5NQ+Ylo2+pD7S/KxEqpXcjLqIdQtwocO
Zyb9pKrUSIZO4fwQnLnNBJIWCKXVNsQvsXpGP+6OxlZcdQ9ADsk60WS75psmqDx/1WQSco8QCcM2
vUcAmGnkoES9QzjDLQu06uaFEhsg/bhESbVVLNcpZfNrDVFba9UoHDoYpxF8GQZbq8Jz0hd86v2D
LGOZhHR0EHboXHNGOeQ4ogU2QYCpnt5+Es8rKz1Upr8qx9z5y0vAcqoJHq1b/BdcNZ1cnDWyHTQ+
XyRvGFdimesjTcrwBl40Bes9VE1JFtzpqCvXyGOtRxEWM3d/6cRFbJZ7zgL1K/xljxJJbDDF0Owu
OjNNNiLOsPewQEmwCpgcwiTU+3Frvui+v3vQxqGszi3xaf4UvAwHa0HbP0SqcnJpk6Qi/ydG7q8o
bX+AQB9jFxKcZojJmfWL+TS/mUJVPzCFgjEXa1ohd1f8WYadOtU6iV+i7u5nrU6roiwvxKuUx7PH
xyEO74DUXMXAH/xGegtlZJnfPNFajgUU2OIGDHM6Qgu0zZ7vcmZ0J0XDRt9LXnpZ9awNO7VhDakc
/lUSZUCX+vmFCRl2HUmzpDtX9juw6dDpe3QeZMinbjZhwNM2d8zTj1NobEz2xje7fURKzc+j7tEK
u0NDvCIkWeQ+HpNPhrUFy3uNmjPfAal4TE25j1d0gd+a9cg7hPW4L9fGbMN5gSdha3j5qrPRDMoo
+1dRCp7smFrXCdVsw9Y9h10Fcrw81dXIzbLdU71KolBN0FweyTUOMx/drds+JNHuKyXwLF1AYxhl
h0tNhtKes843cQhNP7tbfjP92YzZ9V9fZWAGvxSuEC1e+5k778bogLIHt/DOtJaJiABkTrW2zhaH
R/G0sO+noFEgVXhsleAWvOwR2eTgQuh781e5Ea9tocv1xmVNeWYCrKNTHCvd8ma6SjBWtgvTBRuQ
D10BfXy/zkwAvuGWbjJP2+SW5wSr7SqxQSh2YkEc/9Z+ediLu3tGNym/f/mPJvu5i+cbKZhfWKpN
tO1LEaqicRBqXtP72L2JskB/v1OJMioh43F+Z9lgrtrldHqmmtT2fJuX05PG3TL+naARXKPmMDLL
sMyAtPMx+3/vB5tfAKMmWmsPwO1ETqVEDrz7QipYAwRkAXw+Tr6peGUCwU/Fwx9FbrYToRU2Khwq
JRjTwJChy3IEJe8wVEa1L9vUPJaWlY+/XlTK+ZDkSAYoFZgbjLsyyJNB9OUmNCQxnX/rnE5GMXHD
Y1OZM4pH3lZi6RvOtHPG76+mll1Z3hTTka2uurydGi2dajZZ3+ivF3znV6GTalB8/ZwtpRws/nMx
EvWhn2bOZnBQk0S5MueI84m7weId9sxR9PhYZMc6QykWqgEOsXeKlxeJO+FnJ5z9b1czQnoLIsIq
rVMrvdQmVkTcX4MgtwHoXPF/MEb7d04p3MFP1iIVMHUcMRUI3dHnCkgrPbvOq7TL31UYU+kx+g/c
s9NGG3M9NxjV1M1ue0WFJ0oLnudEY96kpdGGMuXpDFDZV6qI2g1G2xKNX2aW5zgt2XQIR/cvsjC6
uVnbif4Oi41Togp/AZV6rYVeq2+wg/IkxXgv/UDZuiBIwRlGx3cAQBPMx2DOICffS78LMxr1mol2
Bu1wfP7gPoppCtEhN/TdOhHosXvWhMQt/7H/LTw0hhqvP4IKBccaIwjvVzkRFW91fF1TlqffF4sW
S7jZsGOdwKfQM71i4HE5VAUjxi+fBJ4Kv4/t0Bynn0yyja5XE4bSCEwZNQLhXpa5MtPC6zgpCcxb
excsX18oijPuRDGNEG2q4uSxwr4wsd8TP7VfkT1vOcU1qBscRst2Ct/9kKjur4Elk6Vc4SJKeLgH
c95VCjXBgfC7TorwHhpz1aghlOXDYNIsdKcLVS+WTqrX7FLcHizHV1mtP1RA8s5/k1EHUtJ1YEWb
u11lxo70FVJrqSkseJ7JMtAKCpHi7FWEwkwSJpikQoK/AWwVzCNEREsOn07+T8j77J0wZAwWRYiV
vXyu+NvyJbzN0vVUcF5z5sXMNm+cS+qBHx3B31n/ZHzbMpS4J98IsVsBYFXxq6qE7Lr/6rKRt7I9
CnBsqMlU2GHz8cQxBQRF5xGaXqmZK2/ZQd2Ig0aGPbE8kUoop/KaugGe2m3VscKi3WprGRkMtjOJ
TLQ40/LXThhyNvYheM+QGqo2WNGwzD4ZtgNYX3a15CMtn0tUWSi/rlhlF+jieIp6w0xAJz5RMxJA
FCFXyfhjrkLX4lw+7wyZlra/iXPusByzZk36Lr8hRj2Ka8HlFstyPQutk0GZV9oGVnY5YQJ5aCG4
qyFlYdxcIP77oGBrchsD/Jin4pIuyKYTivD0THJ5DXSSMlJW2+o5c4/Zynp4Sb6/PNPUVFpB9sXr
3MSd2Q4Q3Jrnu8Xnu0z9+8hf4jDBiQCGcJ/rPeluG9hFjEGk0wG0ya03zlboJozfJy+zMeyincaP
TnKRUZaPK9XkqQNkFBfdLz4jIOpFK8x1QZ9mSf9PLAxoqBjycxj4swW1heclCNwmUHad2BAasptn
s2RyxNHEExEjUuelI+l/6wln4fDTaXGB+ZDTuEZIieGKiv5reRobE45A+4guo9wZ8kBZpLouugN1
4fJTBv+o4oxrasvj9UZElTDESynPcKZXMqDdzQy16mJnnysJY7UIYOA/zls9bjoQXHC7Dm5dK6vm
8rNUn3ba0u82eYjCW8iEauylb5CWSlxh+FGf/JjBNo7mLgq3ScMUbUCJbtV1Lw7YGFloBJSykSCm
tovPvCpFHT50Yo+I+I0eftmVQSskwRvpwz1TRo60oiWO2CtYf/RrB7Z6nQiwPdDPHPs33bGyTG9l
q18U7a94BvCFJbY3cK3Z26MijsBeSKHTl8hTjYOJ3t7bKhE284vnutflgCH0KGYoqHO1uCpkJc0B
O8JOIFH0QaFtnfndm8wjYtBj8dOAIvlOi3ZBZfYsPpa0A//A8T8nj4k9sS+7X8Zj2VHX12LrZDHa
/rKK2STaScZsTK3g4zJrL6zPhsmWMMfT2vkPn6t6KeG8kxk6+xuNScsPrk6jmoPEdRlsVDeUZRwc
3tRZ/zQ+/zaqzZrfXNgQQvsWUiw0x6XCIu9u9s8oG33a7lfNWI/T84YyE9FYKlhGtBjx1z9z1Twa
fKDOt6PjY0Yo4dfTWTWrOdLjKeU99KwZG4FjNNER8VGwllsiGiPz/R+bD51nmujBwpQyqTMM4qqe
24dPMu4QC4815Dzt2G5slf1Ffj0T7k4vC0T0NVYqRIs/kbG/y0tHlI5+g+Cdxei3SsRyEw/6R0UM
xWoE6kHew3jO8bGWEK9ATWhoEe0grPD/RGkDsguDCwtfE7J3O3oxjU8b9+yl0y0hd8kLPOeiTyG5
GczZNDT+StpqAuezj9edeYPYdidExaidrhtTyF5wzt7nsriqILBP1/1bCm5mBzi8xl8w6rK3eN6Y
WXT+UhHQDAiV6BNUMz90HWSJBYblcb7mJgoDMpsCIYwLUjrHf8VXvN2BwC7nRczUL+QGLYIg85uz
0e4glBYixoB4kQ/lp0pnkQw0GbfZk5lMr4jZyb3VXy9t7Ne6iWbm5KJGZy16JStaTqPHgQ1h+S7A
h+BGG4kXG1mSBUUDZInkDZRW341UVz4loecoBOalvWWsTy8Yz3U3GwTgA6TzfHxG6FJdPERwfFbU
HoKV657e4Qb6/BTnEYHDDXxhlt/oT/sra5GnJy9mW17yL+FE2tX0FcrteOVg7H+/rnQVp0e2kM8Q
eIxmAm5VKhHPZdmqQBtSrYqus43Uy2rX3OY3pN7vjTfHMkt+MR3uDlURkSgIcHmqan+lHviyL1j+
J/mOez7AvKUJvug48xLmafVTR1Vd2185gqLbXCjprrAwG7p98/o8VbQ8RkkBVfGrRuRWKAfAlUc1
O2oEsEoBzvpU8+M8gEqaXxN4jsZqA1lBDiPsK/2B3kXsxnALxIy/RjE2APgPQ0Su0CmSGLadfy89
5DwDiM82BsExnIS1vLjtaRtVFOo8PF6g7LdYRutn6rNGjqA2JGP4BNIT/YRcon78/qRwuS2xaa2I
7cn9P+Civecq9lYxXLgkMlOc00A25JY0JIftzmUA11UfkfnW9jvO/8d7ZSq4ZBoIYD0CYYBIw+G3
ac5IhnZK0qGnghhAx6N7S119GvJOz4Ah4Q4sQQqWdBDo2hTGb8jMdN7BINzNJMMkHwHIcUxLneyk
gBZJs2R0J2HoMDQUfnlyp0kWRaqteL8QNfjtWkPfT/RGgZ++W8adfNETdt187O81ztpdh+OyCSJp
t7NZrApIhrOBiRwWjStCdqkSbB6IKS2TTSC86TSUd1P3DAVc7ByWYbIjbFLnhv40k+FOC/glG8DR
ChNIR/XLgwA9E+Tu4J/nMv8/+wUqrePlUzaoRD3UcLRU62XMcfiMwtIKCjDqDL644vDcsqTlFYg7
MvVlBtjcPMFErDAaIm9WHy5Z6zXjWI/N6wSdMhc+tm3qI55MCBQPfMwiPERnw88aaWVLe1gV3NvY
WY0iN63A6IjoXtVdH/LBSkIuO2ltc6xzmJJxJm71I6dCBGt3LGETEpnzVgUCnh++lUxrNi2VHG50
+Rz/XTT9n+6Glht5u4jw8tpPfl87r5o51EI9nYrqIa4oj9MvQLwVxZnwUzlySrHBlDCRq/nzCtJg
G398nCFQMSNy5VGSrNMp8rAyZWV7o2+crtM8tTwWKne194E8E2ohGMk4d38ymfca6SN1zZ2oweDV
DMiuIRDY5y8bYH1lWRsDdRJQoCHZ7K+bCEuK2iUAhP2K0Bc+k+iO6yUvVWy949i1yTAAaIw+ypZK
F+Z9CwTPskP4OewBC5UiacpRORh8FBafphSjeW3piIMbH3iuQnsYiAVEQwGHaB+VRl3lIyhh3ZRM
2v//DK9Jxl5UP4r2YrYy9Z+S5Y89nJ6uG1AcMgm40K9y7O6MAT3v8yQEU14fFhKAG0vkD7NvwzAN
fDTBdwyG7BMeroc9nr6snvMHM2QonHi5b4uF/xCFz7JL8qx2r26Z8BBrJVd5BPYjbUFFjdtMtMB6
LV/PPi0ttnmo0SGeVMfJcKNcrzsvEYTHMkXF+BBWQGz05cuxwDLS/j23kEPu1zoA9Lhscm3tlXFX
P+ODyAFkAvZLUBzHS5+wtPEV6LCMTdgWt8UKDgPju53rie582FHyCVR2lVcBAwl9qkZbgD4s0Du1
EZaRT4/tgCotgqYbM6HlgHZ1yaTn7oyII9v45+RzQUcjOYJMcIievgrQfNg02BsQGD5NnWwpO6Ey
I95Cnb9vIv4xhwS/hLVVuBeR9u4l4mgxmUNO11vSqK0/9+lIWtCKhELHhXzJF/J8iZiyBrPj/eaQ
bZkJ8tVz6VMeHJrG10SDxlcuc/Vv3v4j0Ng+wcz+t7fv4cD0ofkGhgToV9NrPTEHQ5tBDILcr0Yw
bd6MW153ZyUMqg0/Rhbf3LDli/hYkAA0gXJiHui+0mRyQZ7tRw5yy6wvVDEuwfAOYbhmdf8EH6HK
rwrVag1nHw1IklJOQ8CiznuTq9R+Iufv0wJVz2UEmxc++78ifnREwKxqcCUkRvwBDDLuyz5frKh0
0q01bHBZds21Co26rpdF/RzcSOz6zM4QKsYKrJso8xz+Ctf5jmeUTDPzlcbVBuFU4jzAJIOWd+1R
P1B/l2CE8hVx25JVBbs0XBfvKSiLvGu+LqBlqbJevHOybmRDuYHVzTSQaalUCU4xwQFuOQfqj0rp
OLOvRsycDKjMjJYNTeLpgrSLA/DQ8G7ge+c4qTgPR4Y6zL7cKi/Qx89MULQXwhPVj5pliSSf65/r
D+xK/1xI9r4S/sICcWUfHBr51b6q0Lv1f1Cdf6WHeW/0Fhm8bR1uo8tql478+KNp4SjUKodgB9tm
+Ae8qq2CdmrhLaxwbYskjOnh2fwIVtl3k5RsZwNYlQQWu3S4enu0MpDyy357jP4cfTOm/h8wIudN
dai2stex3ODxQmBUVjVc2gHwLP3GCV6UCmhooz8yc2G9JvdD71RQMkRpCoqPBQmuL6WFqY9UvQtH
+u/7P+tqniMByVjYTkjZig2S80NSj4ZNc5qlVlhnKcm+vem0S6xdJdojlS6ySo1fWKZOfPIo05ye
FwfJWOq01ZlsFYmRWAI7R3IPZFOFCywBReMzI+9Q2Pjpdhnc/yeOPNzPDFuBy7NC7Kd8ue3+1WDg
PsBFN1X/zfd4fxSSZXni7oy9fALWDiBoxYGemDa2REcpCBmxXGEgP7BOyGl4g29J6OUg+Hu2/rZT
5kFjw60s9rx+HCa6qVe+8CUvu39LiAOH+3VUlCgtzHuQoSMGS/BHBworcgcGF/l/pagrTZEe2004
zFBtfNCwhnu/680nqxXsq9eZ0n+HNx5JTosep89h3YamF/OVcD4r/iqevYzoKVJFAvtQtij4d5nd
MISIuwHoHLnlY3O1/6VQ3k/0jNSpEQ+zmXDpMulsInprnJYEFXcQGOZUrtLweCWkWcmNr53zAUA4
t+TZ5LgjE/URxobBUFzHYBjrcFTvPQnrDJUZeD7Se4CuZ5Qhm8WntsJLv0pjeI5ya9+uIbe59/ff
Ivch2Ud24/6jtM9mAfTa4zhr5/6xn8pBrpUFnKrV4BAVmT2oMDIsFbHRrsmYGrOrXZgyJsI2TDPF
LyZffysHnTlcyiRcd/NNXI2zdws4zbdOyp2J9ju2xO/+gXXErOuNlokNy86pUtnbmB9YQyVe2U4p
VWADEgYye2Ra+snqUotjYKxzowHlA9uX/ha63rRR/NS2E4b6EADe1NYVL0XgbWbgqY3pYAYkxK07
NUfva5InpbRArFL9CJ9tv90AWfhuMXEiYkgnGB5vDoJXnhLCzBJBc2IJP/4fHITcCPr/ZNcEobqe
XDOnrMVcSjwafJSrj3ACbP3Na9DTZYnLTVDz1BmdvVniPH6wiriXOznAZtlD2lvy9mMpL+w2/yV9
vMwL1Q25nzvNKaOYTTRqEqdmTbmh9lWNDTUHId9ydYZqAHBfDUKhqayhjq/WChUWpbKnSawoxUxF
9cFvGWfKqY2tcX0E498cOBxW7w5Ma/eWbTgM/9lU1etAyGqM0h3vFYWgfnHocgWbUSO04KXyM+Ah
MgWrPngGd0/W2Hh9SMWsQaqQ395/cxNi53KLRDt4aE5JD5ad5EwJlypBytrRND7mNoAfAP5J/J/7
u2LrcgHybiCdKCY7N89ZqmrugoeQceiSdy5wbBGbKjdHT1JPXZUD06Qw75/TOv9yqFRA8ccJ5JjJ
uuJcw3nFaXWOMZKSbaaBYBlnQOaQDXCkNV8dbSS9ZJv5DkA++4u+on3+6ie9gDmKcoxiHIE6Kxqr
CRYnz3qhZyBtdKG++M6TobnEsGjgMp8i8PxOhMnEa1tJJUWS1pyv6nqDykxptYIaKvHJNSgdghrb
2z4BUMnCWhMVZa9U3TOb8E2eTxcOaLukEkpSlgKCshrYaCGW5R7QpkkkMlu02/2UsE1yWRARMaHw
ZZ30wt9kWDv8vAeeOsECMJXr38b5b7A4azMosjXtx0y7SHYyYcgP/LxRyn9owxUuSruZh1/T33Nf
I7hKwZIW+Xj1+XJWF2Z56Hmsuue6Y31ezvDo1OJMhKLC3eyhe7u4r6djfuohCJ5GHHTVoESmB/jE
2O0BFyg5Roft5xQQAidq54pqsSqN8kIZ2V6B4Vy/lb/8/z3Tm2woFx11ggMF7EbNUySl5S8T38xH
2zkhxxD840KqXLJFJrrC1InlWBdBiYxIpLaNrx3OZn3ZSTkWFVz6S4eQLO0Pt9znKqcuhYxQJjK5
0qZYUA+5/UmJl+afhZhPqfPs7ryNSudN96lY3oOhCwCtxwfQMteGvIIyghJplmcz4rKLE+zTvwCk
iKGZ8sZf2+CoMpFjqGh74+QIr+WWzRjsxSHegMPoMjvHl2WXvA67C0yohORTl0MnrFW0wbUdVmK8
Zdlg/DLKPEBFW+u4MDxQBamYSdAdJPIVAkomOwfI0w2FoBLSYRdoFlRq1wKnlJlfABtoPRS3JZji
YzkdWEPlzzejLwdjWKwROtfz1uElTBgKf8Cj6vNF9jVccSGKTkwRRg3WUvDmGALhu1kI4k0L2/l1
InM7PdVDAEhWOwWbiNUlDQIh0abmENDF3q5sOJ80RNiB8X/3qZctZpOFAgD23Pwv7iqajtDZUYdj
AU2UxM9LwhyQGZhfcrmAUZdp7Q2fx/5NDlo/hKni8LN1x3OMEkvfxwv9GgU+7zITA1hi0KqSJxof
uGq0FqFysfd8njSkl47a1Bfgvrh/fVuv2Ld08Lm9LefyWExUZi/zMVFWjA2MgWGrrqJTHK0L7oIE
IJDBnpXL39Ca9igTeZix+qXrSYd6E2yNTLTywoqMBvLKw9KVTEPoWRzFwEHJ1Ko0Xz9sXzI8lwRu
vBDWGQOvd8R7WHRtwrp9G3auj5WMUk7nwTZCLHPceSO6cyyBRMeMze+hUA/w3QXT0Sogs/H0hBl/
OrYVA6LsWsRYl5o5aciXYLy6R/Jsr8WMT6NVARGpQ56ZmDLNbxyaxN6tNj4ZkpmmlpXEmjAHluDU
MNH7NVbefuCZzRWlb3kzPr7SyLTREJLS5mvBLoKWnICUivYClrI0GqqZ+B4skiyJfRmUm0UrCD5T
v2CO3zdzXCeVg4hWOAnQZQdz3/3JBH/MiEe90HA2LLUM7soid+kCmw6s5sZNo/sws1WjYcP0wN4c
Nm1ssYaAPHXp4iaCpUhWxB+2i5j7J62+bFOQHsrK9hFxv2iSLB/LEIEF+RFMYsDCXROPZHHOnQJL
gd9y5S6Wt9cZSYl1qOK5f9a7oGmeQDSrO8CRMTIcoF+qKQBvD/pFieLeF42JErvti4On8KWRheyj
/KLRH/1gzCaeUZfZ/d8ATX+2gUoypMmYhCvDfTi9UZlGPQuC4YiZzB2gQ5/0efkiG1+bRXhoqImm
fkvoEfuP6I+vdI1A1ld1tw1cg0QJ8pNLTSr3xWutuiQk+rQd9vw11ad7hJy0coB1USCxaw0MqCkf
W7Zwqxn9dlOb6WsYYYHP4xcXUbzCOxnbPTXSZvUUZnF6f7Mf2/oJ+ikCUG4L//6LceMaZH5i8vcI
PTxvyBHP50SwhlZPUMc2KpX1xPQ7SJQu+uIBM1Adw1QIHTU9m/EEheu3DzguWX1UaCdNW7qMeG6u
3Kc0fxY+QxozCm1sIpSPJZFqmb36Ti+dzH8m2mIUX5wZp99hhneR/qyVDtKkS5daWQXX4gCw/jF1
DDH9Xslg3jSFxKIYNAe0jT6vTxYTKlpdkm/+H6/a6zUCbuoIGPZOlZeXELZ2CQHWNIID9yboAF+o
9yZQj9EiDLH0gk6rkYHsjZpb/3xhZlz6hf5QtHYXsOaXX1HavBLVjn7jhHtZkHJHLxJFFsT9oaS8
yhrrNMauRY3wjFSHvxjmVXFtaMVUB4RaaVbtW66hUJHnMlyTz8MhmQtfmbWORtPOlcvtF+a8HR8c
owFGJWQETTxs0tONnmw/fe0JSUnT5RtTYldkZRmduw6EU0F1iuBC8VcrgEaxoIjUmruSlJiRmDXF
SqJPHGVlEhq9Y0a4YOJ8IUnRxvJdt3nCMWpyP4vDtdfW3kzO9rhgOEKbgskjk6RDHAv49006TwyV
N9HQfNsRtMgwCDvtXHAM6MlNLm+PZd7bgcHZ0GfaC9fKxNgrT65X4lc8XRgJGlsQyNeH2kj+qavD
ZdILkWLen5TtX/wlpfjBBU33vAT4F6Mtpx3j/utMvb8tdqnBWlmuOgn4VYWJeeaGR58ynhmkvQ+r
cCsFA1k50rvNUwSj3UaWjD7xQwBpEztbcKfKg/NjzBnciRc+M4tVVc5mVoaoaPVjoIrafimAngOU
GwrMCBZQoGj3xoBn1sHemuhueeiDMaNtrAjGvZoJ3fk+KijccglU2V6vC61dWdlXxzSrg0241Jpv
7wGhChgppvyBRpqsyvVaZvFUQMMjw3n9H73qnQQbcpqQWoFFDwW3xId76qxyx5QL7SiqitNpoAJK
Qs/rkm+t7+URHTF5TsN1cRO92qg/9nREgOnAWnBSJsdOCSUDK8C8Y/hYdSevDCA3tzNGD69k7bE1
ubq9ObN+QaSBCEvSeOcLHwedX0elePiG8APSXvprIBngZQDMsUb2u5Ll/NsRwKXR3avIGn+TVBOm
wUiz0ZSGZLoonM0ncX/Ko1GMZO8RyDytJaBdD1raef6DNM2L3vERbkvdKvRIN3/OYfVfbsdpqWV+
qWeq4CTmqPTsZA0iVm4i1nrTvDwk4ZM7mMoblu2P21xHQ8g09VF36CfZJUdZMdUt6xGOpb80siW/
mXjFVc0yRkd11tsgyH0jsbgPltkXS9LkL2yWI0UxI5+eybmBBzEq9gdpbI3HjiTb/XVBhGgzuKYO
HaPXkh4GY8/0Mdc+iE8mVT8M1vaKgU2m9yqp9kWJo13Wrk54PG/vvwNQAvM8XKhjonbozLHocU8o
O2WZnsUlxNZJeNBlv93g2vi73+iIev8tqZLeEg0/P121+2vkg8xos0MKtJJLZLu8IN7Kc3AhVmPk
kylF60XVAEufTxvSAY05qEgHHEJuo6n71N7Dr/XfAleuPZFD9LFBaUj9fIPI0Wm3jB0+smRgfoJW
XVwCsvvczS3CMSL4/dluPMc1G7Fia/Ps+1vhFyTstY3M7U7FeDxxVVj3yO7uz3OmofGVJhDnS0BV
4c+5JGIyURLHUd0mts/wCstMKqXtC1d0R16NoLe1j5kkDuFLtsZ1Vu9bpxRla/RD1J+ZNpPGxbtV
rFtRLTzb6Mo2t+4UWkWGPjdpt9T+zXRZJdlg0Z+XNeMkxMw+DruKxtyKSZztDQtTjxQtK7VJuKVv
W6zYfJqoWb1BQFX/cuH04mvtEZUOK246DLslIShRrEemb2Nu1MJwmU7J7MHTCLhfjmNEZm8hh+Le
smc0gRhST9hAXzsv5MSJGmKqqx2qEY2ecBj/Bwlb7K+Kza1Xd4r7xJviSgrbbtmc2JrzI4/UKuGp
Q8TwTlmSM1Bp1+iphIbVJHVf9H0YguXf2wjWIANmcysrQe6SCDBg85npgHC4JHRbx5/r+Tz9386t
7otCO5oWFMgKW3MkWEdjUZ5viaq8otKhDHMO88RbR9qH+lzxcvStl70yoZQWJX5+WNM3hZzGpRjY
xLt6pFCZbXRpmARU1iT6BOQrX4hrvWqSyiwLReZ+Zu4Y5At/9WALaxnAE10VA2ptqDWrDKDHPMpu
RX27yR8SVAr70RIUzdcfOJJ6t995p8DPG9GsDIj2PY26SYIimh7N9yMEF1mxE+R9HjeYtFIJAhsh
B5jELsj2Tv5UFw0WmaETWzUDQxO+qnOOjLQOSKPm1XyyDGh28Pxk/kEUy4WNuBCssedh6T3kmduQ
majAm763XsxE0OvRhY0kSikRmh9Wg8yu1f0oWWTlafQ2lobtnkT7UqeMZ8W1byy8tDQMugTqPsP2
8MYqP/uFBNVCsYaBPjufCs9eRtPsRagSvQX18ofo1lPW19EksQnvFg/o66FvJRCNA6K+ckZT5BOA
EgoqKhei7APqVMrWQlJ8m4TTH0xPI5Em/vS4dZONhXHnKtVOsFUA47MpMLrcBIw6Nq3cPuD/0DUg
hVgAhhkXC+fZ2YlCE6NRb8eLPXIrbGCc8Eyt3sp4UzCpKMc1GsZsW1Jp3uKGclVFdsajcnFxqJwn
yLDupIBifd7lh5Ec0lrSnfhPyDpSu7YELJ5pDOrUW85D04aHCYavg//1ncVZvCUpW0GfsUWclFgf
Mu93kLv8XcrkkUK+jD1FPhkpJKbQc5P0c0IphRWMmMlZlckRcg/HICGPyv54Go1bav4rGPN09ySr
ia8IvYbUcbbDetq4Cs6qW4ww5vIAUaMZUhfmxWgR5eeamMJpeyUrxjgW30XqRHVuQaSmn9AVGyBR
lPHhYouO96EiJ1jYHFNZkju8L8gPzaR2FVrAEHBcqEJk8rDTZphtOuXkueE4mgXa7RQk89bnydZx
ZgQZB/PQYIRhwAsXgbDXMrr/MQyTMgJDPCM8MObnjCHStAN6q5Stl7zBmrpU//MhBd/2Xrw9tPMo
H9H01ctdy3kI+WdkIbXTXjrvRYFTeJvPFC1IYqYwI/RqMj29allgYjslFbpnjEvSdoOaCOZWXwOe
BO9uq4fD6+0qYTZ4a6UyEejSmftN+RP8xVviBla2EOgw9G4pGVMXNkVx+wZHNY+fbj0kcIvDXZVm
ZbU2GJD7SJM7arCqkx4qxCIb6IWt2RcFcWwIdOVSBM04+BRyj8wtmm3dI2QsFm/1gRN/nU0jehNg
rdCrK+y8jeV2oQ7FeY/5CLdLcdhfQqyFTa+p2E53lWFQ0BcDlerV3oTiJF7TmakBL47QopJU83Br
mPpUTVmVLy6SKEaKrf8a/FwrtBu13uSuqd/PE00vzL3MOpBjR6BXucW/UCJ6VNU8K7rpFUL+smTH
20h0Fv9fyMWuwm3157NEORtlm8/kdpBx1o3o3WLzt56tOtW7ZFa2sqBFGDMtxq/Vn9gE1wqD+ut5
8lUgp/TGtDHLeEV4ZGWE6RXIvLAauZP0cBWcqcMK4R1zScr5Bn57fbP0D2SOCQYbRdnHAP+IPXzZ
BQ4bnvh7aSMzICqlac6bAe+JiTy1zPSm/EHZqytjtmcbftupeqOFoTM5/HGnIbBfYEq4kQsSZfiJ
V5eEpjjwjKAX5Kzkzu+I7zidY/goftLXG+yGaH9ZSQEcfCIf5brDM94QKKESiyic9I6CsDOutrpF
RRuuhkbQYQYZgXoLChe3YEr1UVg9v71rdfxnGFlELWDOC3Xmu+Tj54S8HYIS+0WLKAfiUJ4Q5yoH
PKzXJBd7qth83N6LmqwmVtGruCMOO0MqlU/qXttWlt8UPi3zSxdi8PoFmvRVNNYp7YLXRM60owiq
cpV2WvJgPnO13LnzIXuwapdv4lfe+rmtiFyjBqqMHQejAINIfW5p2rk8rdJbvJBlPLPyduWRwfWi
G/gduDgIYDfAGrOobGYVNPsvTUZN/sYB6Fvi2l5e2q6L3BQ8iggV6OvjiP/kyJimQdDcFDzz3D8F
JuFB0tEA8hJ/9KvTDheqAwLZRqoo818mokCkkK/ENtq41DgFqkmqXjoONCiUkvHyqQ5pygMi1mL7
btaENbQK93lm/sIxWoi8bL2jnPhxoJSbSDrseirr9deoBZ1+r9flAgsYz996z+oZFnVEuJD4Saoz
qjcgNfZMPc06T2ixxL/AXHcFF5+yjCGoBQ/5fSYB0qJK+jKvT5oj4WWrvy+h4EgkKdnyCB1mMiUK
0ygWgrVrALjwhNT56msCaTn4ZVF04A9jHOzmGtAEU9wzHalrMm48xTdHQPlyRw3j5DTZbV3ZqzUH
W75XPJMO0sEYvYIi2KNWODtwwcHMN+FDlTFMdc9l3X7Bn3xrefCZvFschJVx/uUsWpV4DbrPLYNx
xB0PxFKJOR9eQzbewhi7vldLvaLbT5df0Iipw7yXUu/tedq35lJaa1nRLyyQmIoDcGNhbNL/1n4F
omtOwCNBFFccXIgV8/cNzG1+ACRVxDVtMwxJWFaAhDxBCTOwDA9eEt2BDfCREB3roNbsxJPIZzn8
zHnMeeCK1GtMGCfI66HhYSRDyA8zgB22jCup/uw0G95WsLeqlo1qEdpOMa29KoIeCDjOk03YWHo4
s3MQxuSC5qx/8G3ZqnWGlua0dktFC0ktoXN7eZ870txpMTFZ5jKZSaQhjjJLqKAYUP/d8UHP8S7m
oGGwbSY/iH5De89xCuHhCLYqQRBmJBNHwoh4Rt9XwcvHWj3XqDM0j3+yalFTf43bw8da7uTO+HJE
w9+XNPuyO1c8T6/muFU3BUuPX24adLCEeDli7+zhhyubPozA+AfKU+RFBn+mSSbivYAXN8fkp+79
LKsUCagEHe1GkYOJemPQ1x0tHkKZcLpdRQvpULWY0mauls0a/RMAHsxDC6XnBcMTO1Ir5GMxtBZd
SgifyIg0j/a/SxSeTaeogDHFaHEbqkwA6S7a6Ryuibo9slRy8u/87yL6UK6ZNl+ey/lw8wR4uCTg
VV5bD7i09aMIW2mvgsU0zU+cmwspKwtIEAtfa7jx9RKUpgW2RLWQzoTLtuEjN5KH34Lwvpgc3lhX
xyGGJDnawvWSDJSpPtQrNL28jOUdzcsc35XGR3WrlZtL6ExI6lqjytc8+O6fWpqGHeWiBvCt1HJh
TkF6/li/7IGqlwabEe9u1fIbgSrvIqQtDXUsgAOKJLjvyDvBHRdFHhfbO5b/HVOCNLD04oNySTwg
X3TMGFiOc4Vuf2Qhoht4HFs5j3d2eq0LtQccs169wYXMPWV2soFSINKHydbyi9UUkLvx+4AOrXCQ
YQ6rcPmLbIWCtKNCUCkhUJ1GKCmbtB3hbcGOwQ5NAnhg72JMXXJTyh6+7AMNfRVXaqZ4/RvGJ5Dt
kRnLeMce5VLWfYpTZ2EAQHlsb6W2JzNWzcnYR9hl9QNbX7hktaKYCrxP5ArpnOqr8ozcaBikEDqA
hutBpiFPvRIhbQSeHqbqTM3Jil85s33d+/mJkEYLD2cOiUYlg4jKqYIpQl+WEzLN1qwy4UgyeG54
bKgXQSngbzc4O4uZRY14S7sX6oWHBRRvAFxxCvuMjBE+URQaA2jBOWMxVJ6TH2bYB1BevceRY+jD
mjLsCyKAk+wFyYcldu4TPCz39fU36B7wWm45tI9wQr/RZDMV36LojMbRIk/m9meOuWC0o4q4XZXO
4rbE+mUotwGw+ILfX7ci2ui4854EvZzDg72FlsS3cnBiAsONo2uGMbQAjqowcf47q6dYrqQtDU25
iA5wFutFa24mBjV8sDMLnf+Rv58cg9mAORlMzeV8mG9j3To/6Xh53XgoBtKnVyiDJ0FFu9bguTwE
HgI0THNhrgwVh0pwPvswSHSinojgNkDNO+GRsTnnxoLnoYgQGTebu1PORPPnuSqmW3ladpNI270e
Kq1ZS8NjIk3d6lL9KqeeHqCzKrG9n+RdvS7b2PQ06R3FT81t6zI4uw2QqJU9JY9hnzu1PoQRV4hl
xAgBcQjlNkTNvbgMBon1BSBcK8u/B0kBKhE9tXDJkJI3gTke00kVzQxjHJj7C9ibGlfARiafznt7
s8TJM28Iqe3ce82AJoYRa8d8gm2qrtKuRLktdF/bvpV8B2vd8yMAbQctJ6WhE54/xhfIXxyg4Anx
iAodCkUOOO2APTiPWUWUAUQ17REzvESkwhz7PYqo1aAtVBibiClUQvDeCx0qRoRASXGl1ZzT/gVi
nSY2Ht6n4uV0anRYNj3TtMGi4Df01VglpzbRf5Pe4DMik+LhN3KVuyob3jfUQTzm4PWJbT0MgEDm
zVoJzMGdQ/I9+gnW+R+0PoOcXOeckqnOIdGZJlVm1Iu3CsF3lHzEyW3ORoZggsbLWngdcO62gIfI
FQeRIrC0KFOw67nPtscIpxumJ9TSvsxYhNZEwco/qMyF5oygO7Py3mLjXJ8EXcPZZmLo+ZzMd/AC
ZJXo3vgSR1oytMWB6MLhUprjF4dbRc0Hoj62cGPuNBAHdpmkXE5DQHYdQ1EOOX4J3ihM3h3AxlIm
8dZE2PErCqtAyY8VE7nki7+OkWToSPRFgUG/AQjAB3rbSHgEcr5rbaJBW+u6nEkDJqRuxDzfVP3S
SdTVFxdXo4ZKz2NDY0beUbxVjbmSVUxLJMVdNAe3x+ezOViAcGcVADl+SeKLf+5IrIuQvxozEfn5
Oa22HGCfdRlno9T+xAlsnuLR6c/V4m6o8LCSzRNCqJpjTTwzGdinBb0AntMURaGkKyMjsiBeh6wc
fvH+PdrR79stEW5ZRjZrrTU4rbEVwxEolKWfPrCoFBvrcOtRzA2iHiHYQUg++dUj/4OQrunI2uvx
5oHDFhM8ROYaiFD/NKzCD1y9vpnT75Yw0zlVQ4sqcREe3TC5ADN7HeR0VxUxgKhafv49iho1Uis5
cLhgoTVeo3RwgkJLMudArzuXzH98QqbhqQC/vb+B5V4aY/z3s5A9wCpZUpwfMOxQf5dCwwyMQTrp
M85hZWc3ygLG+i1elfXG4YVGBJaTXCncF7vmnhWK74WOuOx36FOOakNtbpsX3EldqBb1VQhVTffu
R029iRPKVvrNVQICkOWZXdhfAtsWC/qc2CZ4bywAzyspRW0rBtdaFftcrq2JE8BjrbROlJ0yrw4r
iLuVbQEApo3nruVN7cbTnemlmsb+aXa3acoanLgo+MYqy+VeUEvqN9QUnjg1oAhI2T0jUJAEucEF
sH0XmFc0CdUnm8UrOXEzYAUjDF7XlT9noyNmRmnSvZ21obTHourp/KCOJh+4K3VshLiJddTKZgGq
LSJPYJGX2pqRYKF65IofWA7WsNE3mqWau6bDvqQ3kvnKeUegeELz/zcRAibAhvnpRW7PxlCi7Y8E
KRp8/R51wkWGOmvprvyfBzttwh4rLIqFzGsT1vvSV2TSv6WLXKBrhn9WPQXzsSZBWBZ7gkIa2Oaz
QhqviqJbokWR4OHJh9/zZR8V9z7mQjJkXfx7kizRulXN/ooNccWV7VPfD6D3ncD5zzgaQ1S0onlK
nm7753ABfBNBjPUGmBn9CY5OkLdQ+LyQQJfhbi+NnbZeS7UM4TXMQ4BzlXqMu2o+HASAvwcpbMd9
Q/pc3CA2vpiKcIMAlAQXwqprwnwoNbNHGiyi2aFt+HcY876fv3y/QYSeNoEvj2SrBSt0Y/X5vbSd
ASeNZ0qX7MnExPf3Sj2UeO0UX0v192jx19tBDce1L0p6PwHjO/EBhy2WM6+MWZOYndx1hnNFnJO0
C5f5/1j2xGQxDFCGBgkpuQ6dw9RM9yBzOuxXUWM/Q30uDv4V9mKmnzkHPaFL8jbG5WPyMlTgxoAy
U3VPOEhu9xJAVVbXGOzqTUUdESo9xdcv6GL5WG9yOWOlljFtEUjlCvOi3BkE6faGzVXdolWvZMgi
ZYwUmkLosGtF1fSy6bY6QR8KcphDhohH2DpuHObrQUBjgWAon96TSvJBaNV7hbTlyg/Fjw5SfCp7
IjnIJvb+xSBYdi4IfQXaZ1JNHmS29PZaWU4ztqe5/b7aQP9N6Rj0qHJb5DqPIG7pRKVdpaQWzMlY
ad0ya/vJSeQJQmiAnGPt+Xo5EgkpE7lO3uIenWInSOj7duFGFQGW0TAWKRsFaPa46wPd54ya8JW5
+nlz3QtqmGcYmEoIhH+BxmtaRQjaV0dlL1P6ao8Ay7p30HWoKdxRvXo6Mq+b4PglsnjUUqWDji1r
B4HYstQMV5P2rdrGpBpPV85EAhIlgs20Ocg3An1Bsp0MtsGkAKcvjvZuo4YY+n3x2bO+L1dNUBRv
8zVy4U1wVUqdPEOBOiJpopVYCfVDv4Rv/3sBrcWUrpxXydTSaFSLvIeN3XVQmsYzerAN5J1XFnmj
IDE2H1mMwyrH+x9ZwrEpEctsw3055/+eUpfSpvJTzZYqBb8blN0tVrD20DSy/7pHbB4vCWiquxSi
HPg0k/unvq19kJCRHbkDD+DFg3aNrPPugB2qbw21oHTa+RaJxxrYUybfa9zUaQuyxaMSjsjVyIIt
3c6lSEf9cbnqfA0pNa70NZ3b3VtZjroMfIhBTARIMhknJdA4bllfUcrZUKolsFfkqYOXJEId2bNI
ouP0Cb+8Zpf/Hl+qfVZRS0P0Qq6Ksdl694O5YuIa2cH4xy+LjmVJIyHe5Sfj34V/7E1LLX7jrbVa
N/5371vS2DgkIhgvl310t2ebArO4pSk+KadFXSy3BIwU4ML7YFBcHeDEL1n6C0bsgZeBWn2FIPgx
dDaVs8TLajkK1SCAWjJ3TR+3yLctuIEJ7DtcMbXJVTRTmQ7EZ3dxDXrnzJ/S9mWrpoPo5GW9ICDS
y8nLM2ENdBkxqOnG4vt/At6DPrC4mXooDIT0gf3M9YlvpMrKxyCmqWcos3uQy4XAOlN2PtJRDns6
/8qA+JHcdskxbbXGutQx/Ly3QYOICK0diAozhtEjaGb485Apic9QXgD5SOpEtEg45zbhdjHM02SJ
L4HPZmk1UvsvcSJ/vRKPOhWrKsALDUQvp8gs7P2QL6u2eL2Olj1HTJN3+y5wFYLLqMxlD+w/NrpM
bVfAQ4ZRNirUgCdbMNZuTCuJ5TMsa3BBpW+FXHxuFOYrUPi39Nij02EQCr/eioA10W9tHvcz3OKb
3hrF5UjdX5GGcP3p6XLpXOCuLghi0355olT0QjNXOCLafKU4vF9ojeAcdlbJCDSp5qgE2jxgPkR1
cZat0hMeME3QGWC2+yej9E62S+eMwLFVEssSRnZgMPy/9zy8Ofou1qBH9l7g/652UviUIt6cj87D
KsXEkE3YPPTi33XOyGFkk5wCEbnhN4kmYzOLDF6cRCbvORJ+DO68nFKDjdxmt7jaTTST4IGaLJo9
/6WR26Ln7AQe1x+k1CmYEgLEHNLU9qdoMWHbccgWs+9RmaekZqnR3iI9Zdu1s9y6sesuPdKcUjfO
unO6oDz2L+wtNmJ8KZdBGbhTZyfNHfoVO19rdTqFish17nK/xAUxCOJNTFulXyz66QctVZBZb5UE
opYZcO9Dpy/l+c4fpwjMoAPQhM8xN6zrur4pErmDsCpPlvQo0OMtVFEbhjQNR/kp47IRX9aVbzhc
Tt/rArktFM8uYSC9Is8qm5gbua2RSOGySYtsnn+RRlLPUh+vv2deuMhmdmpJfWQ7ZOmr7HH0Lq2d
IbS8PgHwMrNe5pBxq231B/zj1DNc9RmOL6u52kbVQ6guL4YeuOBSi7+amOhSHfPYsPZyCeGMCX83
boOdb38+AEaS/qmH9MivCHzb32plq+sigtFueO6GPd1pT9cEO+tmRNbuMe+DE0WJQAkXx1Fd7RQz
rm5vw9Cp3oleFUsS9is/t3aQn8SIRum/OroQM7UvzwaEpTJ7wMzYC5BZwRyrTHZruGJbinSriAxe
1Z8hOIX9d7nJ5XmnI5SUJVSjpl5gjwOKBRfApLHwu6Qh9SOeKL7EhqHY1v0DlQhDn6FfpGBTAdP+
lp9PkqUYYnxvnGfF4AtnjYo4/zMIl2lublc0ANEZQmq0aw8nyPEynC7BAUaist2RXS/Cs7rlFkGD
tX4P4glQwnpfw44zXneobGs8R8Zoq9vNvOtDrC0QeL6nb2IZxW1fdw4e+oEQ09WoPc22Y4YpzIuP
zU25V0W2DDPH0vRCJoa1VD0gyGA/Rb+OfojE4mwEMjclA2k+JokGTygrgVLNxkOI4VSMDQIyjsg3
4Wx6m7T8w+r1phlgDVo/NzWBpLcqvo63R8tYtDq7ipcSwm9MUJwzOvEyaTrGFNmQ4nQWYY6fiVg0
pY1muzvhD4LaVgkrz3feUQngHCwNGmF0+9A1FpACMwo9Mu6/whwUlve9fBwLVMKcLSC+66zNCe5I
UGCu0sOb+XZMLeJasmMnTKYY4NHvkK+A37XbCRZjK9RM2hBZHjMjA5JThhwE9INqOXokaM4NW08f
TFxqf8Nf2r/fuw6grtzzMWAk6SwEUv4VFekH2PpC2J7u4CP0uQKXaBnegI9rncVHiWWRpUbPwd34
4A2MhkXPfRyfOSql7zen2YdLNn1eezNG5C3/mwR1pGLiY/4tmTHXgzceGyL0yR+b54l7XW1zeWIm
a0JklHswQSKFfFO2jArDTifiOr/euBe6fAFU7vBsmEFH1CCNE0xNjhBoES/eWS2+fS9pA5EnIRnQ
ESIJZ9DhY26pMLezyRYQv1oYEE9+AmhTv+jwEZE+kwTaft//RexLoVD5QhkaCoIoDmsJFScJKMFx
0v0ggC7AaqLor266QDHZDup1OuMVIXGdyCQoY28k4mE30oMjejScO1+aL79nZZw+8Z3VGLz+vidx
lVGCOlXKTv/zzv5weDeOLDxsqyryarfm59oCEWSm6ySXWUF1F99jrVdEZ5iBFv0ygVm/EMmBRm4J
bvngisYbq8OaAO0iR4SrgmYSlLXcYz1cSfFoH+4/8QpZ86CLU/7tr0bDngJHRpNEsy1h4oj/4WGe
5kHDt6mxjOAk5hzzEGOhRjvDmnavE8YgEerJrHyDCf4/P4o6WvDfQvAZ45GSV8ZUtJSRgUTGf3RO
YMIdz06CyGUo0qXAj0+I9/NvDKIKlm9kkmu7jqWjVi83U2HW8IqFl6cv0qGSKg7RxXbl9bre0GxI
8UrZyJ4HSP819T1qpYpXZJySFiiK86jpRsZp64Z1ytSAJxRPez8b6xv9IyM7DNy0Ya0WsxAhY6Fv
W3S8b5g0m384gjs+tO7zqUyX5E4fMmJYGfdG/1aEWEsmgs+aZDfUVOaY5pBktWWjIhRxZk+pcnBQ
r5P5czXOdUQa0wRCESTxXmCgUiMkjPkkllAGmAEUwYdB+limlkxwPWx0EiqkKNS9TYrA7qfmH89a
zwhYAzFU5kEPgFk6NxwTAKmE1ZmkX6XIFWBmneL4RbxtasgJdXSh+UFz6tDw9rFGQkkpnytPkUKJ
XJXOpA0rJU2OfrYv0e+3MtHhrk3gNcOVDqzdI8ywonnaBCuGgMCDRUN8/20clTQJoazG2uzMXsM6
x+4b/FoALXD8QSi5tjyeoucBV58lXH2Bj1UZsZSTtryYrSfR0hD0Je2UantwXTK8I76TjG6BR4+6
zX+yWDPxD2rkkSORPLwj7UMkU9lUe5VqC2QKRmuzIRYgekqm6kHR4lQrI6CGm/jA/84FQ/lm1KQd
oI+2SixUutV1h2N3cDjs8yXD2iL3bL9U5gk2EN3N82Uux7KaXdBxzeHSEnNpiD3SM+S3P9Skwy/l
uDtSMoPtvmN8n3GBIMzwlMXOe5Kmt/bRCsL+KV+3m5omudcU9khxpOaC7qm9KZ2HEKu1diRRMVN9
uvDn6+7ZfJBCQrZ3RfekL5BCZdhMXz+jEBSzrrFdFHuc/vVkIzgdrixia57NbIyWH/ZGmCyOQQdb
8fCqWyURMwZukavIUDo9bIyOlVXC5jTXiFLBOPi17U7jpsEJ3wJRGIbojHFl6AjHrrU626hu6uUo
prmD5RC6wnKjj2t4D8BqmIV3tzh53/PsvcatXYD6pfqyHNp7mTyxFLsBI5Fk2QgavCdruudvOoGD
rn+um1mttLr5Z3QX9NZYqYXFdrayv5heq9H7Btx63s0JOWUSVztyld8DYrcLcp8qvq6A+7B4KSh6
SRma+HrgGoi3t7KONzf3fnZy7IcyquffqjD5nVFCuNZ1MTUx0ezFcxKOMaFjuN5yfyBzTiQ7hCYX
D4yvufe+jUQ9qoBPgDRFmgKoXwxTwRUZ/EZ6ndlBmOr2TfkPMbKV5k8wO9/aEkSOpb/hvXxSWPCC
bFN8joR5KQ9oLwnqsL4gF9SpPFjTfXlZN4fv4+a8AbgwmWKiReYXEv4Ym8DBx90T8zFb9OUeq68H
3Jq9+DjdG+2e7bor3pIQzXfTfh8hf15uJ4+6e51+iR2Of06qLek7PTJlBZExBD4FOF/iSdNrGVvm
NyqFczmMb/jd7scyvCrdq34rrlsb4dKh9/tJ8hNdQNTeQw9jW5nRhwukurqtqGtKX1QbRNZFCKK1
CoM6JTnI0nZ4vKFrUk5t3d9xUu3sol3AOv7i5Uk/P0LIN5zTlPSN+e6UihW43MUDtjxd/CbLJctj
Gq1h9boU7HPlqFjf5xGNCfvK7PqN4mGJPzDj/70b9225vbHjgCC8+WH27YghQKfRmkZyauiYqEOf
rod9dt+x2iOiFu4INhdkfDdvmDgJTp/TVHmNf8hm4fADeoEc5TSI1KHe43L++fAXVMQhvKkNlz8E
AqQFstMhntCUJZKuQ8xfC7HEkeep+qvv2kYTMNmxHdttqpLkcBoKAYIrWvL+qGHKAFDm9z7GcPm/
FMIjrnsjqBGqXQDOQX1pfmypL3wTLWp2t/r6yWLvQcYwwXihs1Y4Z1m4tr1r00WbxHoq1wkUJb7N
qLCqqj2DgZEpoZG/RH/r2oI6pxjf5h1K4IMTa6KPKI5d/8Q+zwcf4HYut2U38nItCz2tIuafnCvs
4j8b7gXstATm9L8khXa2YVu07emcAnKCIrcObl8q4k2L5Br7ynirMgNHs6wUxmqdSHqt8RAN0nVV
tWeyroydJdz3RAErREwDMzTbR/iWpCxUmjXUuJGNn5FbT6TYmv0UEXyLGsSTVbxD2+zmiAtIPyq3
F3ZKwyS7w6zHyxRK9Ihw8luAo8QbhPMYb8IlnZ7UAkOUqbCMPge5xfIrBobn2z2ODv84NGvylU2x
aAblp1Nfl1vavb403Tcy4wuiYNx6BcTX3wlZXuZqKgQFFTlb9Z+po3OjC1qFhQxubIJPZ1nJj2yi
KZf1NNj22rlEW/nVrjBvx2JNYHBebE5R2vfm0zZzEuZ7CbaUyPDsH4Sy8N/cCXaDBNIinaDBZIZi
WOgH3Lvcgy+ILJHPKirI0KrgzhzXMCT0yCQDOL5lkEg3KnhY9j9BYZcBufKedun8USjW3dduY28s
dU+RJn6hy5uY7LJu/pK1OtztwjoJeC0b4q7ktfwnIQhzmUi73XpmcdQbneW6EPQT06wpSJ2XQFwU
Dtmm7+HK8N1lSiNes6futzVAz9i+Ekjv0wsXTtO46LbiMePuz+xdjbLZ90kBp+4qdgicva1Ovb0A
YxJDQLeNshQdtr/Xg1W3paER4bMYK1LY/DPkhzz7OeIhDWPFEWr1n31VUnhWdJUU2twXxVpnIhNx
Ozi4E2LLmr/8BBd72V4spONspzIQc57z9WbPUtrn5b6Z37lUkAM4mA2rlg0AKFbFTPB3PAXQW9Ff
G+q6sZCP/2UubKA+ypdYnMf9WoGFcK5JKjmFeWeYUQU7VjZm5c3iad9rQ55euxOHKbX5ceztiNz4
LKslxuAS0oPNPVK3reOj/tzdmnVLTbsjEA1pZJlvYXp3oq2AI6jsDhPYoyPR+rxqfhD0m+KoXlX0
P2MnHfU6FtOY5F8TyS1Ro/CG0SiQTnsmX3dwQg0W0bVbRb+WNClbpe8B8cXNCx2V8pu4JtNOD4E2
XE9wO188fykFgueEX2Ko75rtlY+VTvbNJzfzhALWcgTyDZnfe0yAQYuUhPtzwGkhmktvdNoVieZt
Ju+FC0t3m20ix1sYWbSNoohIdILTM+1vIa1H3DmqBnGTBWoG755+cOo8Ty6CwdLwoksVu7aubWZA
piXJJh6WPTxF5Ae7VZe+BxApQsvvtfenfq7VbB7LJowg37acNvMcjNc4d7lhqC2t3T11sXMbH7ez
Vq+/IQNs2y8tjIy1vp+UbFOaEhPdq7oQ9iH40eSIesUoweweilc1HmChiOWHkOIIuUqGTSCQcKbS
IsnBA04hpmTQpllYjF8CE5xLHrLPaSkdrzdCAkTWOm8pvjA5c2RkzaTtEKNwp7Hy1279Vcw1S12o
6x/f6k06nYBrpXO6ccW5/LBRUyoXdHerbt/39jN5QOfW5nnOHCUU0EbE/+ryDL5oOFKjDUCddXif
MkBLEdbnt50oXQNxvlYyjep4EeNJ84BG24YZmkvwzTNpO0hMAxloIcLRRbpa+EuFehoWHp8D12Rb
Y7ah34itnCWu7IAAMge8uXHz84fvL/Zi/sc4/XLSee7eldRZGr950/DoSE8wtjyaDMK5v+YA1Pwo
g+UHRAWq8hpUZ/Dofg4ApJXEzoGAwZ7KiK9uocpZZFkGRdf6LDpyDjUbOqHcv9zLw0e4H3PgOFQU
5mjgZC4shAxHLOHSrpT2ZTAQxopiEgB8LnS2MHCSijZmkypTRqJRIXpk2X5HBo3iros3U2JZIoCN
qZhgv/M6A3ERsOafkA/Q8+ZQxuBnX1PaRc4InrMurKLbw/glo+HJVl+77yONB7aQa9JPh40ANNJ3
T9K5rNiTWA6J9SYpE2SE/ioJmFRRUrYgM2Ucw4WWOH7WXdhGuTIx3BwZwW6QvsQ4qjaaw6RfZKUI
Up/Kj9GuysRu+XJRxXf/lr3YdOGPwNJhdExov+yJ8RpLtE7WnnQle4FWkh9tkh6/l1bLQe+mdRkN
lqYDQVl6sbUMX66CCsoIZ0G/GvuNEU/yhed4+rXT1t4q7NjKR5L+U/pi4mZqacA6n/AFx+rRRru1
XaE/iEUROJ2jy6t8dR8C/jd+5IV6AmMRNnMv6ene1RgdmFQDkZqaSgr04EHJn/45fgQ9QsUAm1fI
4HdHhYLmz3Pw2sOZShyhqUylrZauLoyULKZD11/vclfRCjCwRSl2cvsX5N4nK95pBnG/6tuh9yGj
2j3Rqgcz72gBw7DXGavQog0meDKXGEJhGsn1cCRYgO350MVuEJMYfrjc+rRYeYsVrS0/WMrtO4ZK
ptCshYps5fn0j5xfTn6AahY/+2BLn0afDFB+zMJaf5C1jomQVlGc+2vFfu5s9XvpHMk/WuxVBhjj
ptBm3Oyl08VMAwDrhBiuWpNXj05+CtxNN4GSpkzvbR7SgEYcI0XOnpB4/12IMv6/O2hrHAe0a2UN
qX2ErzJjsGH4QSxbrMPoO+1eVmnBye1euP43Xj3yVGU4GXlBjXnsMhQ3z0wE41CH2rPx46j/TG+I
+13M/L9ASCgRXOuJ5t6x5nWuIVfopX9OgyIu/4yVTgyxOFIydprS+40rDNAYlwJm4iA+YFFw9ZiN
AYysffC7N3ejWQpkg1gKdmggoXJxbM7Bp1Su8qcQ8UJS3DtG4OF73trCYEerkjZqy0PUGU+BLnE3
uu+Mqkks1c3HCnPCEQSouBGYRioZed2nc50yfQYpETo8x2vaObRPYQ0XHEbOIO5qo0pASn28x+k0
xq3OL5D1hhY+5ra4ppuPfj2pjGup3dAZyXDW7cxySoPjRRAvZ17N6LElBcb/Aq2yHPv24IAo+qov
KQH6SJs3G0PUS3cpgqFVdKKB+t3ufoXJEvqpbsWiIw5TicL72KhExmzLguQFZBOhYEQD0CR1tnLX
MZzitJ30QfiN5phkfn3krIwHdtRu7/jhcQBV9STGk+UPVkBeEmBsHH0dgDySI4eN5lSTZMMbcbgz
KnD6HMtbNlCLdsLuw7ZCmQUn2E48NqmCM6KqWoYU+xqM1qGjN//IEGT7F/ca7Zq0wI8UH2wCLFFx
D9LxHeNpBxhvwV8sSDa/XJvsTFX76KV3xPE7QA2OB62mxXXVQvN3Yn+5XKzTDTg6FDT0OyQu16Mh
m9CPIqIah7HNI0mNQGQ5/SiRItqvsbTx15NNRXxILTDwk2VB7na+wFAa1t9/T9P66XnMOyZzBQ9y
J3F5e8ICw6d+2Y3WsVKxcMSWUcuMCdmaeVGwOOAe6ptmKUEIWDh03tpoImZ8G4vAtIFTV0rVLzAR
MuOnPC9ZL4NfWGA5DvuYPlDf9jiDcIZN6EEV4OENuN3GIHN0B6JhLik4lDdIML/vRWJ/iFF24vSb
Z0eswhJ4pE18BF7hH2pJPrgLPC1aza5PEWq0qIrBmSLHFI0w+BTXlYOI5zRsUFWueMeGiuVE+xV8
zLi2ffxPWptIT2B3IBdIES8xq3xPb5S+yxsvpPcnQJhHqrvIWDBq+R7eipQhvgZiuYXrwUbjJw+n
HPKND4LYsCvCVaVo/nRKUHGk5+mxowYoO9bMH/flxIazSBl3bg1GThjJNVsA7ttZdK9P7JbYYiTD
L1oq1IVUsTzEHcpceeaxAyvKs3qT6VkZGYfo3B2JO24w4AFA8q4hHynnJYPYSjvzD6xu68PqlY5U
jgamNyiMad3I1/XWx/PYlbNf9KxtUob2gT6jITBDAhFq2AckfEAIHf31gaFO+gWD0i1C0DZG8HJl
Ikkym+Ajtat85pwAuXJ9a2AMDJgdVQNZNzr0Uk8wbOe1pEJgLV9PSTyF99ab7+wwuY4m8OZBgtp4
z0rF2orlVuvtY055uslaJ9gzNWaY5cuEtB8ta/wsdbpMGTl0jbvOuZy7RWtcx/sxWg/Zeww7RujV
m5p1UDQQbQszIMOtaVuBNj87V0v2pF+PJ1uZiCBCz9e6FSwEMJAdWB9rVgBFJR0mWpeoBYW5UB+Q
jB9cxhs9dE/WvGyMrRsJ/xMbmWLcJ9v1zkTjogNllAorxydL3npHicknZzMWASQqHnIfUUB9CBHI
2dea4hZ3s6qtFDUKJWKz9JKQNd+waA2sl1MLUyI8AOo1Td0k8bReVjxJCbcFW1y5xRA903a8srr9
aemR0ROInjA8a22W94a5UioTkM3xt/aY7CSsEeVd4Vmf5aWuefwenLC1URsjhp8LlxUY393I0bac
g5K336l6/CeS717Fpez9l4rHFxEelMvDp3gplNw1G7CreMatkd/hUPaXQ91ooqgbZRJ+8fR9ibYP
IgaEBzHIaLGvrW9uAIcgzzZECdDiPULlijnMWxJedEOggvEXCsth8Xq1FPaa3U7COPW/YHYDvDu/
My0lA1vAEqGqA2jENIP+kxvwNaVC3Bhx26CpOfxcqxN4B7JUmMgO0HbVAGOTQ2FBEdUxNnbULRl7
/PuIJAhqYXuUoyu6Fy0VYBK9yK7nDxOX1N1CHtTUSUPQKgwZCgDy1kScBCZJ2dFX8QT1GKO9Bejs
GmxgNsAoVn+fEGdQAdnyIc5LJfOoeZ0a78pXvj3ced7g1TdOPBCR4Gvv+/Ih88hx8uIBJjUMbiZt
plz6TDfYskuWdrcBT4fLjavRtFjqrOhFdR01rN4veXtL1NiymtypKTrQN07JpxBeMwfAjrf//lUK
q3h9bEwOUNc6Xxs4DUpmkYAkiD5WmXCFLFlBBmX2nXxIXk6BBq5c2WCoQD8nhpLuoK6WmiFMhoUI
8b9W5sRJoQSJh5QkHZ9mo6ymHCkjxqkZ3gMvfhTW2QCROw52E1wj8QONep6+cB8teiW7V7zuRqvZ
EeF9vDPirGX9CksKGueo24ukH5BeJGrrsYos1XBxuevj3LfQl3DPtULJqWuo7bQaw0vESXyXXbIR
Fmt3oInHWvaaalfgmpMoZG5CnMtugDr/XxBMRAXHCmoKwaed+AMbjZ4quPPRi74gPWJ0EWVLTi7m
Fgm/F6mn8OvfCq77t633HKn/YpnKbdIjx2rhKyC530wyJhkk2dEOKkZoiExjL2kUYClSvpGiswM8
kRRi76mxAsBK93GNINkkCvdfYikrl7DxOtm8sBPHPG4FpnxqftqNtTADXjSERlo9Tyxlv/2xKYqM
Co1v2rCfaZLgcMH7AAkFQzZ8wVCzXgzb1/hCbOYxB5jGI/Uudt3cmWBCeqw9q1dWRS1a0lfAPrYD
o/AA2bJg7TfkBpuvfwlD0iPkkWWXiac1RZnsaTSppr6ahiCIOYjuJXCOKNbTWE5DukwvK7/+PliN
sgl1+Y7QGJipWyB06YolRQG0Nk/KotnXByH/65m7avXF4ZDQFv4YyIfILlEgQhC/JKdbi6fAj+oS
anM2davyMLCOTMOMuOOeq15Wms7xP5YfPIrk0UwlPb7n71mIa1k44XXhc/Ja67R+JDWfpDIDi+bL
diqxwL9zyFmvCKx+Z1zlJ5W9JuQVjT8SC9r5byN1ktOWJ3c0gr0B8kV9XOP+0fYKt9attsZ407sq
nQHvqYySsQhwebCnLOFKWUFIn3G8juXZlps2X74Unnyz9bM9nTxCE1Kx1NJuIIo0dElnLaM7+3x/
mY9/UcTPTt4fyhhPCcP/ogE6xiD1t7s9kObh+GH7ViqLEtrsMihdl9/i3PVRlhQ3n3uRVu5H2FnA
U0yhiV2vAV88Bn9lvMt5pc1Wj9pn/qA8qSCJKC0PDn1Bw7XZ6ob8znSorcElWYbvry7qAKfotq2U
AM1hCXqPNxFvcw8z3bBkcGf7IGTWWwNdvwf+htUW7AiJDiaXAj5h6R+C1DzLs24oSJT/IOyfrmFT
MdxvXFbpOEpBBXPjQy60VdJnEdUOkbmNeGqzcNqh5rSgHP0lTykITypCmPVO01SkwsUvwzxn5tdl
py5e57aL2ORTv6dLWiTUIc8iGAPy17AwExbjva9aXqK/+LlwfGwgxYioFo1ZP/uRoG83BDfeO7nC
zPvDNCy5NN+dDCZi1hwSIhxYhY4FAPoWpSm/6ejXC70mtiND6/C8Z9bhKC46sRP8h5EUysDKLn2k
HI0uNi51007NC5SneGId6x+yk3SwxLEPxfYhv1blghJ+VFku+/gSP/TYSdqeQh1XxBOqAAYRtLtI
ULJoOlqsWwn3jJyaa+8/dZ8Jmzv7jJsYzlHdC/MBCMEu4RW9xfjQgLvbhf6O0V2nyf9bn9DTt++G
koVa3+8oS9B2bGLvB1BjcIVM86Mi5Ari0QLrOinRovuruvR48V9PYfUEFH5H7M4cnri4UAhFb1d3
Tvl0Um9HVnMKnasoXY2/TTcVftBs1vm148eY+F97CdExFuhUeNBHhvUFQ64bPVYTdv7WAlPcHYTp
0/PCvcbLE6FtGSkuIbAGcLs1lQLqae+oXteO804v7Asb5fVXabOOrmVuJfuG4Cf+g/A93qBgtnTq
wmePV12SOA+RVKIepcYGxQwJxSLpdpV5/HDzfBsdaDclKKzjPoCpgCgh7at9ozIWuEE49jNEjWhJ
xY198PaplGS8X3ge7xXCSXZ8kQXYqNnos7t5mtpJupel+9laqLXbLj4zd+tGgvZFqovWXXA3Udhw
n9CKiUQxKGAOabK2v9divTIGsEB+0VvvdUEeFjv/LqCZmbBTOek3wbIIAY2v4nFMSp8qX7Dn4+vc
qeb4g14NenjvdjBZmm98vgx18Ld3VclpAvlF0PQec0YcWhKDgyK0l/OEsT8crYyPCvtPLj9Aja1j
zVMGMzXfEPn1jT5KnxkasT+PPbJPW0USPIJ6qkS9HTvuvQwsUeFHlsnIfJcK8kxF/QqtcF0ajy6Y
KfrNSjgCCLIxLlbrwt8GUAWQ0wa+0ShgMxt4J1z1spimuU0mOHvmhsEwUTnUaE2sbwQWgBeLZ5iz
u2BcFVNP/7GAqtDz/DNI9AtL/uj3xlKsoaC5GKW3In310P0YQQs3O1gf3gXd7mWj/JpN8UA9EO1F
9QOiZghkCNlhbeRIa9FrDBr9SlWzJcYRxaaPg+tNkCXaDfqa26fAVQ8uipAQ3L2E/2n1qlEVffIT
YXdJomi8VQ/0MpSGZA+Frd8heUDdCkuG2B5RwMKa71HJ8t8qXP7uqC7m4axTpnI/NUhEjhTCvfXc
hJeEPTjkCHdRkyiBnW+1eQDuqsYSSO5zY9Bd2REiik8NDmFgqfgDDu2qLsweGJZJ5Os7qoeYRJBj
fBmIiEmc6QltXYdPKzA/nrb7YvvtPVl75fJdq93VZDREtxjJomHPSDnal19BdVkXXgD5L6btbVDR
oh2YVbh5WXSNYNJhmrCMhP0Kx2s65I6MXNGu0iVFLb4/3HmqEDc6xlhcKHK3iGlJGTMH6Qim0p5z
l3yx6S2gN/2o6EXfqihdCc2+UlwV2jb5WWvhpq2PLC/YKBIjf7mwIw3hY56St8bCvSK1YUrfZK5B
7bbMGla2NBiZVRrES8GZzwmjbhOYwd/3Rj/eK5D6ywR9L4ojW1/Y070o5sl2ZuOJhDf9qi0DcFZt
V1ZMsQpZt33PB2OX/ln7SZ2yPkhYxIaYYT93LxMPjXvzImARxmCeijU5FBXrX+y2WSq/WmJRiETK
tEjdIaV7fovrLn3WA5S6RDLhslvSgTLSZIzVvyOctBVuc6eDWAf/Sws7kPZ0/GsSmW+rSIiWw+lL
gX1lk/D8UoEp/l7OY836OtRkRXynSVBVlSC411TMcJDGQK7oU7E5NFYsS5+B1GtrwtGEgpM8N7Av
ck6qjc1XXT+XBsz2jYw9F3vuX3aMqOwXs0F2LqOVISZ56BeGLOk1SQjnENnESrWdlQb0N/gZEiAh
0o09EbdvV5KPhHZ8Pey4EPMxbSuHrjlNKgeV7KEMUV3LC3Uc2SctLKccAzLoFSY3U0qZYmLMUWJY
pQKtS4JvfcfFJdOl3ts+AkeL3r4vAuN41xrBgAjTKPxGKDPC5P2WAzxBlFVGFhZMJIuKvD35G+yt
3npF5Bs0kEKoX7T/pU/BteIcTPSFEdvHkWGTJBsRQLtjRYGbvZUzpSuEO4p/jl9XNY1gAml2raBf
FOvkufonZsPHZEa1jX1cMJ/PSil7PhksDu9fi6+EXjxBxj1w58BOhIXAeguwAWVfHA732b0fREvf
xEBgzLS3UIudH93eqf6lmPfkZLOqG7E0JIS8pJb6kxon8IlugQrRVaulysmJaGYtiInlSjSn8v9a
Nxio+GFHNIbOSGn5LZL8xgtsQDkiOJKl+E8fsp5EpSBlZnYLP2nypRAwBQEkfv8mrtc4lW8lVv0i
nPWf1YE7kiUGhKgJ1qcZPDbPwH6N6v7UrjR527Us6Okrp5Liud4GZ+5HsbENBJPN+GO714nAfDrc
dN76rhW8DEfRhpHEbRutPfMbraCy7TUQuS8RuIOdE1EQ8SjRVoUGZg+xNIFSdD5agGGZ36OEJCCx
4vWeHWH2qRekXFxBHxcHJjgDBAMUI4+oAmnJbcuV89SrMRofqlrBN3O1P4qzZ1dt5lX8I3ZAMUTU
FTL1LjSJKLMd/ddY0q4asmEWH8QJzIVSDWRCeu9Y3blyavpfP9zh7xg1s5txWgzcLTF5KEG0U5I/
LwcmtAplpH0BCgv2APrJ45s1pOyexa0spS205/Bo01v0HnlxUIrZhdIWuOwFwGbaNXwbQU6Lzov5
3/bN+yjWUdMah3o1Oztra2BOJeqEMWVn4j0Pl/Y6l9Ha/vlmNOK3DEFp08sYwX8Os3dNWGsAaPYF
LT6WR62cy3erxgReLGZhnrwLF/PtbqSrRMe66tvZ3bMbjIP9gKh1d46HqIoHo6UqTjxJFZDI6On1
IZZt4Bh9JSy71+A/XdHyKOs2rqpoZsVIIiKXla+eKkDI6whbYMe8ZYjHa5XTEiXXdVEpe4YiAA4g
ECrQl5WT3h4c26wEcFDRs8lw6dsLrzq8CQ+Cp6S2fZ58014AA4IQxj5zTprwl4XLafD8ebuNV2eR
ofArGPlmI7QbMlcx5SSTH/XMCPpmStpkWZzk7xPEPDLOibO9Wgc3uvB6CklZdc5Z6F8PXaFk2ZAI
SYIN4qUE1EdYFLLGCn7A4ftwJ4Z6vEwoAyMHp1f6ZzZKL2jJ9RG4B5f/Te4iLi0RfrUGz3Er4Ctq
G3YbqNCnjO0/TRVSb2FjWH5N3JXrPr91yuC5O726f0w5IK5Xz96i3hVT4nPVDkDJqvkjfGMd72+A
vlc6gnLN3h4H8J9DeuIaNhA5VxAl0HXBSe/iBtv4MVIydj8uk/oUF2U8UztJGWU8brX+ycrJoACx
6IWQWN6wklrHl0eG6RrpmUhoEOJa6mTOZW2KjnKh+o5EIYdlPeF6vKBb1yHSXGl4rjWa0jnTwl44
5+t+CHoNEM1LCpeF0PzIe6gPiBq34gHeMYmeMn/qPLcZA1Ybbv/SpSks1Q5c4A5nscKXndKMqIQ/
urgL75KsS7et1pOaOGuK9sJmh3n8D1A5arEhPSdSCq97YcHGyoRtzSfFUx+cwXRlHU8R/UhY4mhF
aEbHHw0ixTC9/DzY2TAeOZ+HL/G/F94WLZI3CYDXLkLYh3kNhmpywxrUA2A28WSJlPDuKnLepR9N
cpzKw65eQlWzo7Z3/L0L4jlA2FLXoa0fIWQYIVf0ooguztRDUYbryYaF9gBEMPDdt5IeM7gdNTxb
eMUE3fFIijnOKCDzY//O433IC82GY3APQnq03dCsffEAXObWHzH0lk0aDsjevEojvahmE3VoI9BG
Qa7gldAyaQcDMVdeG7/l0g/zV2pxSzkeY3E6G993WUtrq7JYi7C4f33DKC3FliJRCYHQg7q8Nwos
dq2eWt5vZfrc/JyEFQJW3f5Kx8oh8cOkuUoVXon+MeQza2qXF1LvlhFn7v8L5bD6LAcvtUFXj+o5
mCPUHYHprLxqPL9vn+86Tg00VohEf5XUAzzS5CVxOIx08nth+f6lFpXQqUPWcOWVs42tkAcEZFAU
M6s9xNeeJnciym7t64rpR0i36xoT+506om8lqLGYF87d6la8W7C7iUp25UlhzEa9tLV2nEEFwmsk
TlOoE+BbWVnn7KbR+E/1PbYYO+kOn558KwW9tRgIy6QiuZ10ffiem85E9Zt7Wwa2KpG9sAWpV+bz
H/Kf6zCUKMPQaI4B+oSV0sHWdOd8T56S75qeHFbRlih97Q+eOQIhUhqWBGG+aakvTHSSjBqayKrl
P1ZQbfFI91o7JxSXynFKQgEU/6+yEg7iC6HCv28Vh2Je0SW0CsgFLslI904tS8+l5phjSNqWkDJu
cIlF6aqFKPTavuI8zcPIDkgGKR5DFQ/9EgTKiuKGMcV41UFahLTVd37wAMZ5iCC+FQqc/OY1kru2
jIzZeN3piuEj260r213fvpU9uPA0NW32jd07uqriQVgylBs4T3eWUFlkVxdz1ME6bT2I47JNIMYp
YAOES/fpcQjDZG41OeArvSdOM1ZFgn1qMfCi1I8hD1lBU3Ss0PIvxZHBd//zQAARXDbf183Liy32
a5V3YHxvDjR0k1kx/MqVMZPhu5LIA/zGQrenr3Z2/FWXSDi9xJaMc//Z7VEMFLqDKSGXgl7qIhbL
1cCkhSO7Lz6k2Mn3a2yYI7JHl9AJN/1ZJ5GfLe8NVtM/n8JPPrY4tU4EIrk0DOx56Du0dIBR5DeU
zG6prXV3sTSQLpfNMS9kuv1UJ9Huqt6W0wn616jo6tYJxIvDJwk1oo6Sa0qCB2nDoQnh0vrRu85p
5VVTZ7rF+y6mL1D70KCey11u9BFvAdzf/IDZqCDQHbTUKdbe4dd0Z2TnYMXmIDb3rqdT90xdjOa/
HYxuh0umQEbePMjqOfkz2zyIfkbxO9nkBrFKmjwz0LQvIucuaWvtdvjLXfyH3As3RRv0lmSwySpl
W6gPGNGFVdozGgFyayZbll6c7dCpte8/P/FySBqXZgbA1JpO+IN1wWRBOumeWnhTlYp1cm5IUwKI
aVPIBvm7bwKW1KQwviXY89Cda9wvzmFTI6FfYCTlklX58GJjFSpog53TkZEjM8rcSWcJERlY6FLi
Bm58bmp4UByEle4Wjj8h6zNox1fkOur0XPZpd7mZYRJ8qUexDMq8S4VTE3LeFz0iCcl2RPRwWB+8
IA2BEUk+RqgEq8jJwlkjHAcHu9HPP/GvHW7SexVlAtVuF1kv12Xp4XUg8sDLGWbD+NmjGatJfkwJ
FnNkDIOftnkKACF5E+yt4DlhUsRH2bzexj3tQOapmK27EkOgWrVS75VwXYWWJkUfP0eMTrlw99vx
v+sYTlh44a9XqC/uVQpAww4MsnbzfgDLmuo9izaZscEDTAgUJgheIhxPM5SsFmOqMGJzN3NK+iTY
3olVKQ1E+MjIyBF28g7ythMiRWExA/eE2PvKvbrouQrV40pR4KWr3RY7KVG57x+NyyVw5eOAAlzN
4HugPAI2dl0ecS99iVWYIiEYNbnmLR1w7weDedcPlbqGb88wMdNa59qzwtMNw7gblr35a/GEFBT9
eZf+nVPW9zNYo0TcY2B+yhSt94RXtPbq+c8mXsVRjCjDunzbAgY7RkH1uF6jnX9mlM2lbV5PLvM3
TO7RC6BAm4OwXY+jVi8y5DutI3xcYmcT8EqEooH6uf2PoXk35O1QVCbbtJyzxZKWJe+s+WNYR/H5
rbBl+N7Z95qv2nckMcQOs/UY3OySu4REzvX4vDB1WolxKSBhhkC8wcUYfvwyYdldaK9CW59xaDQh
uX2bMSWdUe+XNgEF0VQ8u91AAUpUtyhSqiIb1rmby2P8SU6lssghHO5axx1bZaoiZpVeJCQBBoVk
Qriy43d7ES0sTwrm7hvAMjAFfUEVEPrCQ6MMQ1erUNu9T1C26fUbsZOsJK9AAU5p0tbmEwWf6HOS
oDDPKrEQO7wd2Min8wOwJtqBjZy3tj747/+N+MHqO33carkSgBhENoRJk7AbIeYlnUipDrR8bDOW
PN1+D/PPqOh57CpwQD5BC2aiPIQNl7XwulXigKtUgUkBKvW0pzIaLZW41+DF0/M96qBk2/dhKAmV
iTO0ATsycKdTQrKU/ZeXU2PA35mr8zb2X/OzG7ciSYQKL22SXJ/Ox42/TKZLfLYXSDVxXU/Z2TG/
eAHJqVDetC1JkCeRolh/7jmBxJJ5r4zMuRWi2zbGHvbc+lYQLpyy7DhKAZjowPH/krWPpLIgr86Q
K7hVlRyHsP9W6Bd9cGfAt2Wa40q5owKfDoNi4ASwalpEbpN9KBqOiJJdWBGLR9mg+q7a9rTJF5Gk
hRzD8tTkWhPiEvK96xujzCUuGO3clRL6o8goy5cBhYOmj+lTCdQmpASh58PkNdOuGfJvXY+/P9Q0
RQUbcPI1i5lvViAIZG+A7gwIbStM7xx3tzmOPBzYVMtAIBruNQtl4i9SOqY3Wnue+Qob4zaYBGbm
4jdlurbai7EOuZck7qfw5CsoKEnaxIbgYu0J+CTKDP7bWQJKQTHDrKacNQD6pgTNz8LRvmDAhtKK
Zt7LYtblcTX2bbkYpEy+KEevQxtiP+KSy/Ya2fulfnvC5QMP3wAp6TRh1Qxvai+AjraeP+7NN/Ev
ZqPy2d68WqmQUC28XXRbR48QLWt71ugNmK1vVLKZPghcEJ3P6GSNcKNm3VTDs3mJdWxh1LnVN5vE
TUe2MFth9BElxqxcblFshbT9MukOaSVUblU43aDk81XMtJlCmirj14piJwbYpGJZ56hyoz5opesP
atI1C7ziZAfBbVtPpDHvM4dBYV3JmfaNbONbyg5hXXk5O7Vf4r4vupW+RN+a61iLEM9UXQ7UPJUm
yPCyIRw434O2P95B+wKf2BiuRM0qyIMlzaRWdo94ZlW5333TEWQLLFG7ZnMf+d5y9ZHEbGcU41nT
ZNfkeQGIf6tMlNU1HKdsoUrw29TZYjtuC+EvmDd72oNbtvrh7IAtwEcV/cQEXfzJrA68hRQxzhlo
Ijpg8VmD0miEL2k+yoeiwjX9FG8tsCy8Viz7BQI/kmamcr09kKQphwd0rzLxhp8b5TBFdnVnAX03
Xw2ACLtvXclYDaEaSjyq4AIyeIpgUKvbKTC2VcwKQ8BwAalnSK2XhEmqiT1O0pzLnN/ctizXMC8v
XYwDgooWDMkJ9H+qbVRpM2WERzCKwS6Ig625qQorcrfmCRYhq+eGFdzVdE7KMo/0pN2Vm4As+oEf
fd2UL9Lrqu7+pr7XKW0IoUHsCnB9JjD+X3ai/vWLtHL7JkgNn9W4R3F0l3rcUT0DMzkfvdvFgsI0
1GH+40uveW9HKnYr6TBqG+EMURTc/BzT4Azvjfp7djYb/GgVt1onQCwwGgdx5Thv1eOg0rd32yRJ
UcftRSsudigDm9jypZD2k0+TyZe0cSmvFvbxLerjCU6uM2HosakYCXzBe3LmLqEoQonuHo0Bol3U
qn1w48PbC2oFAV5ChAOhAzr4JmZShMhWtuw3AHRev2o/jILxPGzRKfHVG5OCg6kzZWJ5u+wvh+mY
W4AFYH2Vvtw1g1mnC/IqTMnqCBi+Pfn690wGH8/qeeGgB5AE4KC5+DmGwggj7soznfHjTZF0y7oS
We8LqMTCsDSpEBzzR8o+7okkJmpAp2NCU/DVfGGiKXH5brw/SgXhMztOgFzFF+7voAqBWMcb2Arj
W4R3W4hv9Ro2MWEfJhfEO4VYSMJLCvinvt6ki7UWUJBeStOerdXvZNjUPh/m6P0lAYCFxDl1AT4/
lmk+30zBQlXDRE190N3ZXb7mo7SJnBkAOrTirxYlRlZxV7VLlktAUBR5mYc5pGQOA7fY+M0TNIfU
iRJO/G8ayiQNRrR/h7PT5uKvp1B91dJKafWqCTKlfzUz9+0NxIhvHsTs42nW8Q8j3ANLYs8JxA3u
YvjgsA5TT8sy8QIuHVhTpTgwVbhYaSM0T0H1QETCuL6xiu5yOJksQ7x0tClp3U9O4hQ8UDsINIne
37loGtqbCOMDQSxeK+KVf3hzqkKJQCdSdTg7Y2b+OfncaL8HPF+zfe4Jnn64yxdKer0tTDHF/dBk
5qJWGPcVejvQNk1vi+3U+moxWXZh6y+9odyM3QwCqEZH5ICATqYpOXFjaBspsyhbXQDF7ZUL0TY/
pdg4R+ErhVaCgtaThvDO+F3+g1iA+UU/F6m++QfDJFmgxVZdU3hRrAecfnTzn5Ey2EFenIZwtUqk
CO6RoxU/4+i5OCXXducB/io9wiZoiCNstjX89OGZ2Dl/zThDRQJwIuE0bPQEkrYKUYumaGwChpcz
X1YyWiO07WEgEVpLxOWadAMR3Q0fy0kmWlSx6m40THHw0qj4wLS1wL+jAPCEg4OOA2gL4H4SHKyd
iQ/iY3Uob5oG7+OKVVV6u1Lt/tTd6tgDXE9quR+dBKV0ft0mnEw1PKQq5rtat80h/lc2J/E7kTiS
yeFEaQ2vhV7vYOgxIFkLDAlyZ3LdbSc8HVXIl2E8GEoSGkhV2PT77crTKPzMJpZfZ8HjPZlzGAHz
nF0qq7UtAk3svahCy5JY5/4UvPdg4pcxys6aJzgxv3Fbv/O1n1McXSHp1Oyodr+eIHyKO5eJJw9e
s6L4p0+52X3dUS6vx8HSh8TLR7W0Sqwx1kpv4J6UWt/ho8nmewew6CyX0+SJTqRw1kNLHvagc+4G
27dI3Mf2CVXGdsHVxtJipIlDTMyZdfjoAXm9BAYh6fiKmb7IhfYF4gBkJjhb4KQXDsgMgKGZnANW
8kvKjMgCS5CwVu4TV658ndn6uFryKhSakAvdYCsEZM6FBTBrhF+tlTyQaYLAmy4Tx4hvwoeybJ9W
/vBHg5Ckdm15DrsHxdMFZ7+Jm5xBFONr+C6djMYrJVmmwMDoT4PsZE1CltpwRl6fLL+Q7ysmI33T
OWD67Kq7aqWRv9he8wOID/CMSkQ3Gl8OKac9Ya5p45OJVflD2j9bBKFs2u0jrm1OLFF/Tppb4ak1
2WwFUFZGgGDPrECwmLpTOvGY0XXmNVcnNLwMlpZcu3/6fYBODRsMgSW0wmt7AOjFQaD4ZTzd42WB
jAZg4nfI8bGnca/AaLMG5J5BcXqcu+/RHtjc1M0mmh4ikDTGC145gnvM8+Lgx4JW6ZCbadXser0J
/nOmk8KDUJhKSUcfMlHQt+K0fy1cbeZORiqVcLCHfzQP9MwwdaIS7jqZXAI4vSQdDyiza5FWOgwc
30gWybUbAIrAAhZ3uNsbfFLRcwlZHII1xQP6Rtn+ZFDrvoeqoYLXiUr7NlLp+KbJT/D8eL3nmKFe
LkQzrVr460M56BXq46zVw71+GKWQtdGGQ0IjyxHAXH0GnkMNvf2F4rWeSAdQt/nhjBU/UZHPbTIH
0Ip/sI5tI1Yv6uQL8MdEYJh71Bpf2SdJHZR5e8ni6+a18XbKEY2ZlfZojQ7SBqxZfEXXDa63DTpn
P5Kz5Ux8LHdT1tRn0NQucpYx1wi+VxGLmmi7dx9KJDeTTUtrdf3RCBdrB/QcOcjGaRTnNWzfQzi6
xUWmBvwsoqaLM1gK+gyWGOSjwZWn0tHJPnWHkv4meeEB1tYkG67teHzcm2jsJVbqqvTy4d+AmvuV
S3+5eYDOwsdOAezZ9pPENte2h54RGhiRZzud+2Zx5dpEOFkMZAsc5MCVy1sjtplZi154it+uR03G
bd8oBMPfcM39yOu8dyTcJ8I//vqpiaBf3JSa+tmE06MrPDi6aRGjrw4DeLNPdRj1zNM9UC3RUWcf
PsX7xHmZoSvzs1RHwi6C1oXR6z153jW+MI11dxbHCCtaVccdAk20jhiyNV5t6TX0vi+XEZL+lufh
H1g+mTMl3c6MGAc8jeex9NQpC7TnpjEK2nH/pPpLP1x9clcwd7Z1fwEnMR1r2jcoLRqFl58LC5WZ
fm+BALUoLKG66QJFbtiQLw406LS5EFP4DBOT60GO9rhXSrrSE007njsMBdYcXFDkYtjDUIKhokI2
haGrauH4D9vAwW93CMZv+OxbDubsgrjwdqyOK60+kzokxbxPuf6qQN9SkqDDp4ywytQhiQtoMHyv
MRLdVG9lQ24fGvYuVADqWCrsk6uGvYCroAc7mxl9IqO6QdtilJnchRTuWRRmdxu9whO08gyfGAk2
qnePvAWiLYumzk6dRoR/zjVh1Z+GKH01TMjrHIw4R0PoCSoqUNgQKaxwi1EaRxjU4EDF0ujjt6eq
wrUh8vfTstwngenq8EIUeJYlU+cPwJRMdioN6cWKXKNGM+iAT2xpU9tkW7vja1x6MeTcfLfLcUea
ihfXjA+omOukhgS1T/5ju9EMqU5Q+jJsXc9Rx7DSvkqMICYSGh9HmEq1yrz85YZmMdWlgckeJ3Ky
hLWs4hJayZVu9zZ0HQtxGuv8huYTRn4USYKD8GL0qC3DUdWPXYDsSkJGXj2fok8hT8iJCbR6GT0f
YAS/ENfdIif9TnYrpVQLQbgTr5d9n0L346l2zZMZJTe0f0w0LoPNNtjt2/tLM0sO8OeR1gLlGw0F
FlxTFagVvlN2svSWSAexhIHE3zCeTFfWl4Z7kHcZ43Eem0+qUxB3CImGn3VXl2ls8p1v9ssyljqv
wzURqVHnmbDV4G6kqNCd5GSHgpz14W6VYI9EM8V5IIG87TO5VCFwAFp8mHB85YjjBG6GZcqzsIZm
SjZQL43R9MXJpgQAy345mQ3FZR0oQJZUPHpKESdyxiqurJIIzBtqMcD7ZWzWjmV7yNPgh41J9KVh
LiPyNx9FJGseOYFQ0I9JqF3S8W6ZEWr3HOiDt8GcRg7Y1tGMp54XGsRJfi5i41XNj1TTHCaSSIkK
LmyvB2hxaC1KcrNchU0P8f8XkXhSIKzB7tJGRgCKyoNhY1jL8nYTI6jqStGmTVsQf3QuzlKWey4g
82BWCWBu4eemlWo5GRtKKuRayDm6GaeJEBXEyh2vcMtABk8BR8ibnL0JWo++GmYRLAkFSOYgYa/c
ovQQ887KiNYU/dAoWIE4RS9apI6X7+TEg52hI7jAbjzr6SONnKGe9WOCvGzIZArIi3cchmkUrvWV
w8cwQ8WS6x4egQ8J1Z/VvxufN19yZstxWE+Bb1YPqN2U7l3daF1FlNoMYpZkOufhe4NXBT88y8n+
/uGviuacefv9bzhccMmdH9lqmVC1N8IetMlXQa2ydB6buptof3OrFq406sfhMdyOSvuCzq0Lvtca
QdBCtvxjFbM9YRoCECKvxXbb+AB+lbOq0BUoJCYFetsvKghgeRqJzsyESBOeonSFD+6/sIBdH0/V
fut/ZzbIDTPYHZgEKw4WLbWtk4uaWzPG1ow3S2xnPv3ZfMIE7I4lIVwUIBLStfUAA1Y4lQLjylev
4Ez+JGO2NGFBWnJ7jbwhJOD4/eZR+Hkh9vzW1CvvwDnosU9E53TzYWLt8mfJ/1TjwS2C/199Z1vK
G9c4WizkZkcevYMsNDdC1kYS0rikpRsVHCJ6iJPK4/zpipYQfe8cCV86jj44ycPeMJ7J255tgvpu
5BqFNisdJMIeEi9LXpVMqesIarRBMxvapTkKyyeseXBdvJORL1v0w1lzzkf7R7d7hLGrf6eFAFRq
94QfHCQikalKy2K33Ws5e3pZF0l9Sa7asml9ENt0CX3gnLnt8oDRsNYChiA1s2wur9JeKA+w882w
PYyGOx2stuwVqcwWzSbd1bBN8tv/4vFpAiW1uI/I9/tT1fBWQi0TZNnfBYp6GE++wMEW+YXgcv+9
DTB78fjyKaVx3qnPTife8Bwd1dSnR8NvQmMihJLh7e9sWBkPJCJ1o0C5IqY181CUxyxY/ooRoFJ3
gqH+GbFr9fuxBwp5/vAem1cTRPEBIc2mBp1q4TGECxNK2kNwEAFheKSQI0VSvKcrIAfpJ4jp7QxM
l3F/c9a1dki+KDTOyx8NTPDcqJxHhONYkWcUFkdx6gaf4fzc30iGRZ7Lhoxc3QuX86jLwEmW0AZ2
Y/e7rqPNTlRtoktw1Mb85ETW3o1tqsRsi0oZyG7LYeUxFO3SU05GbUG3pZpmqSMxYfvfpWGjKE4s
DlAr1GA/TCwLLTO3HKnfMs4NVkCsPF/ZqvHq1DOvoV8V/k5ouHi8x1dceJlc456kup2osmSs7hxB
IacaOzaQUm6lzCnd9zuX0g+JVwfSyhaT2TaNpj9WwASUcZLKQ8GeyyWlGIBxE1Bhd9sm0GGeiXH2
IH4oHDpIYkB3xqXfpQAUX9WDL/xVNVXNea2VEACnWiekvgoJsfa5fEEJeLGKOA6GRQrM1gYQXJjp
tl83mAkWEC4TncaFIlGCVXdK+VZzKOc/NgXQ0S3ZSLgXkNgismCYYO9IF4lTywi77vRYkj8ykvwB
bXc5ozN2Gj7y0MxLCW5tRjhpUdKTKp4mspzFY5FYKs6nv/V74h0pRlka8KlbSXNAPA8IvGC0WA33
ycxqXKEvEzYyI0HftwaErtvPoPeesZdOXUNqzd6hse6TI/qD+Aw899nN1r8f+glQtA7HkI+G35ML
3fmriUEd8B9Rufi9OCaRXOEjsbwr0sdrRrvV2YS5T/3KTTN3ji0M3r08sjtRLquWFIzqkeJWV1oY
2ERUS0FJ6ZM/oK939kQmQ8w1srUwsQUfbJo+eMKIyZ2cAob0LvZQN+rJci+AD1iPcyy99/G8SIx+
5/MPKpUByuBNz5PNHKctH/9VUMkl96sLrNUjb0XaU/eGL+RwYYjLALkyT+cm1N7HCL9qvOUWxf1x
QQuV5Fc+xzo+cfagUbCtCVXTposriQSrULtgoxXNSuICg4ed4Uirfst6W/vPdoeh/c35jKzqIJLZ
Yod8UZe77Dmk5bTEQJwXghvXJCDcyXrw+AaBeVA7aRGKFja7NS5PAP0fL6a+c1aQ2nVNkGabSr9/
CwdXoe5FAEZoYqs1LTA67wTH4TY6ao7QBgVYOQkUb2K9vbQwv1re22n7MIk8q/eCUbc0lzZ4FXbH
Hx9sxlJrRMElUrVx2JtuU8na9sV9H2Nqcm50PoK+4HOq2A2oxPA1V6/eqX4NfEtuFtE4b9d91WtR
kJ9UkKNd/VQUzAVfWsiZEk3Lgno7t+IfPAFwA9019/8195wOZBAMclggRXiyQRY/K1JCKC9pVDB8
I+kctKEnTkwMggYxks3OuvW8bflJi6p0Wqe+TtiNmA9Z6lJV2oiE4NF2ceNvQE+Yqu5VP+B1MOTy
xuSDUN/kQueQcZQnBpOXQ5N2QGP/l41XuSe560KzMi3q6bXL1WfU+xjSnTL3bagqnF585UORhJG5
cuhVBxTT100H0jbyXGUfGD6ry0qHzv9J4XXYsGPfrxxv89JCcz0Zz0FLDpMVNDK5v5k76WoS0xT7
q3kJ8lzWUVpxFvfhVNDf4bryghB4oiS/6ZXiDljDjc8PLDWboNCWu5HpeRp4gK8t4gRrq5yE3tZd
0EB/Mr9E/rPP+dOGCmQeaCIaqv8xvIKb52bOtCQIxwZ0pMcb2e6F4tvaHekFwMi7kSmxttS3pSd5
rVo86PHwOESXIEHO1jpcoI6sFGq29a0VA+abuldqsKis6cbsqyo8LFZQ9cm8VzZLJ1nETzbN1JXk
9SlfRl0MenZapqwtBVIxBw/BTfStpt2KHzcW3Fp4863yqGMN4eW2ldo7+DsZdCnuHENVnYH1uXIP
NbkDroHcV7mZq0BL6oMK1YLM36kjOZaYYJjQZ/twvnSDPppXxIUbAUIYiW7yUdKJhObOZGKlZv54
0qloQjfhXIl4vqY07uWjxaW8Rx660wniaehHbREUtLRxGeMsEzxo+rofWe2ow3XQnidZfuedCe5h
W3rqMU42M5Y4sGLlDk1hK7NbOVLNcGhIffj4kKVRb1cyrKsEZMWT1ST0kaPpH5mFNSOuv7iWc7TA
3vZlNbSlNTE9G46Jb+HdcWDLWJ84HisE0h26uBX/nW8RwHVfWPUKcASzHdoSMF30ucRFkrso9uex
MZ9zqbP3VHQY9JhOdLFJRNf6wjy2+rEYWp+uEeAKdr3A/3KK0N7lgRk8HdlZ3jSwvt6piv9EG80y
xMRCOtEkzOBvSewOh9jt39dUcMcirK7XagFbPuLP5UVaEA5/NGhnFFe8Ucz7cFWhdOFYQsrfX6H+
mEiBR8AFi1RBjMj7Vvha/z/zuuYtS194Yu09JaqzY2DAVUeIB5SnVrP/6FIyfWRiCKV6qxUXX92G
lmuZLRCRMKOSu7L7kz/KeNkNpqvIhl/6r6MZe1GAaQGjbHFcAF8j6L46I9QRIZo/Vwqj8f4OR1Nv
SaVk/5i+0Jvz5KEkTHjqlb95by+fIOE0X++2DaioeYpDchnqal7whxxs/DUG4k87WEw2hDvvu4Tq
5niz3MIj7na43s1td4t5VNBhF/kB+NKatsb5gmYVNKn4M1TmwWPdv6mxOcurozI9I3BwKdcdTDeD
woro93T/7tZgJk90wMrkpprP8gLryFzT1J/cUvg/Fqq/2xpo+ovjvcB2Z4NUD9vf6oLun8SWI8Qx
jbcBcSLCJ26YaNUjAM0NtcslsUZ1t/bwwfT5O/4odpC5eSa9TAjBn9wy99MOGoEH7TDTnhagVcHd
ojr4a6FsVTujD+VUUEIxvYiEkOD2y72Pr+LuhietBDnJKnT6U4Y7jS0Qdzvs2wyGls/abuOSgGyC
E8/uVhY2u3lGk8SjugYeGzmDMNUrVZFWpq0BjAIXrigCJIygJHCZvafYeol0ZfuU8xPpChl5Ekzq
5j+R1NMa7cGVapCG9UFk3+3BECmbMQietb7avr8cUYlH1OOyO1TB1Bq1sLzx0HyyuC0oi38n+NqS
PQL7r9QtEwldTmPPJ5xuqGw03rBav7LLvZjjm8NhoQRO46vTWTCPd4mIzPuz4t+1ykkJBRapyGsZ
akeph31EwoSs3NUwvncb5vGxW3uhf7Gia0oAlooh7Jift1bXDrW2EQJECw/SBmEs3tFu8sjvSrl9
LcoersspyBOerg3FVA1tV5Gaw4/i8cZ+yEGlDQ8qlYAKLgm5i3pD7yKaluWTBPozPFJ4ayA4trh/
K0glnBo48l+90sPmcl8oE96WMX1qBytt0vKMZ4nMu7cNunaPubDmEz5MGf2ZeZQFemqghwWi7Il4
9uyJaRTuhuNL0qDcpNXGez/QhhVQQUTfC5I1MD0NTpmVYGd17ya76kR33a1M//C6+xEMltyhweGJ
3yISt8OfNAv70vBq5rHW+2vcOP1l2Jc8QCTeNLlJunbKnepT/d+Pvxm1Wm2wTWAIQIIL0bUx7bfr
DQdIBmRsBQNKi9nuCOkFyrTm3snulA/VI+hFnxU9NHPWZ/OkDd44VZ8h3wUmryGJ7m1JGQSbEo+k
4mTEDZT++aktCYjjJc5s2cYAhO5gq8+zYclsvA2gBOa2e/95LiBg0o9L9wh0FQ7mhWYFCkA8M5MB
O+lNoU4+2wX0BmcvRbf7WtGCed5ozh3QXMrPxELrd1aOGkGmu63or+tr+nOJ2P10LPFkgha/2PCm
+e3QVEoLFfLiwFNp4oTdFDuXtaKWSm2TInU+zFrxt6Ekq6ev6eDxpo0djmHqKF9JS1fQHUZ0HqZu
3L7mFgYaOxsEEzeblWqZz21S4qvxwptWet7unB7jmU2CARG4LIxjb9TS4bt0BoSvRw+auN0BAZQt
H+hKgVQbdLEX+c5JPWJJhmjRhfA9admoCVpfl43yzqz1i3FStOhLaT54mEqum+ux0wiZiitepdo6
Tj5A5dzEpVN+sE9NPuw8V+4AK/qnPTUBC5UjMAjRHbcHrzIPoIHN0wTBKSeQZI1d2goLhVb6HLFB
VnIl8yqFBpzBuWDyxGdTUFD807lgPrUFTfnx4O8d0XHosRHMoMYaLYwZUHk1hlaH0KqlGLz1zl0Y
s2DpS78AyIjBEBVqknwtqAf/FGG6iZW/Sx/vDjNmEhmtLEJspB1BwOo14+JC9tUxAV3YiKLvOVKS
l+98XLSJH+ulkwUytmqxLiF29CkuO+ScE+tJZqr01iZ7M4vOMDrXOO6AXC9S9JajzOV4IDFX4hZi
K54laLJK95zh8yaIpM1bxOnHZh3O3/p+141TEKI7VNbEoC+GB5wCZQZCUagX/5+K6u/XQsmNtmXL
7p47rVLAXXvT7BVTAtof4alOocZ7FuKLw8bA+VqQ1T3XoLiFiqTmbQB9pQxG5XI6YpB6arqXFvF8
qszezqhpRLduaqBrxwLV1eEgZore3PVT1d2OrHJ39u0m0vyUO3iPllmioj+W77jrAvK/gGk2Mk2N
lvZjLetyIgwFDWU/jyTPKf6wYru2+GwiHRJHYUMkF3ADCGDaKbUYRVtCELvaBdwmmrZQU2PD3DRx
hprvH9A1fkxOSPOzzkZ2mPBLndwMwkFdCdhKeUXylwDaCulRbQW9htmM0Bsj/FE/AWHA/AFFZWW9
pHv3I3S2qW9x3IbNj+On19ZNDmQt9HEfaM5lRD+jkNLktQe+qdukUCCI+k1twYU84FByDgKUZGkF
aCFQexltu9N2ksjjw0Ss3OPHIHawEWkeHWtqGd6r90RlpPVPNOIh4jyFIPslPglfx1V4x29EE0Hz
awEp/nFx5EKJatoyF5J+kYzeT+7CIcG8Nj9wsCeL8Ay95RGJ5+fap8FETPrjJ9X6SQdnJAplIUht
zKjnQTblzR4X0EpHTogQxS8JcbJ2i4lVqnFcaBhyVdO/OojCj/Zqz5yNTTqX/uHTHHTqVim9jpdC
cSeU0vA+yOpmTbNXZ2KmIZgaU/GegyaCPjIgs7sRkvWksQ80Du5tocIzFsxWd4aaWdjLBHb+kNFx
CEq/bq43Y7wuA95+JUO/HP+dt5OQ00VHMivggzHSclx8KAJp/6FRd4hXvi0DiK2jEsbHh0YuXtvv
+M4XxLezJKuthD6antPzq6W4/GS+Fh0WqlYG2WcySBxUJbT3H1WfVjPe0orFRViO7gdXnTDLzlwn
6OuYjvuIckxwdxRrQWyoDSFj1j/WSWVXlEak7AZOngzYWakSak4zQDv5LmLjOrKtJHC7AIOpFrk3
u4w+9iFGVCOGwgwY1ilP73dWfYfQzIghV5tnp+YI5ZP+g0zsmQAKHSPidELv88KpXUf3+G3kkD5i
Stg0NawCbey7kKLUJydRzN69ll386GcSqFMP6Sw/ASwJVYCnm9uWHQ6Q27HZqBtX7dZoCzJkYVt/
ungwiIAc/roswirCqGxg4N5JFv/6ocvVZzKtNeo/Id04uOIydFQAGvKbj3PmXUlr3736R5zOSHOp
b0hQpOaosvuvvtjdol+69s/tbmxsqs7p61winGKXztl0o+aToIY4FnkkWFENDsxrEPWO8LycpCd8
+MZNvP46EMlO5LBcWKtdcT1YRD4pdASYP2mWalsgbTcwBieLgqP4b7531Z3DI+SLYo1Wig5NSYKJ
damxLok0KVCljss05Kw0NoY0Nt25lXYa72AFJqspX3NAUgnTlB/lG+fBKburaXW+LoNCFKoP4PbH
Lzkh5x6NRqD2gdi8806t4CZdM7vjd3XN3u0UAhxngeyS0YilJPWsVtJ2NuSGqECFDZq7ILjz7M6z
Tw/X511ZTHO2PD7+2+IOUW1SzfhP1Z2tb9dMndVJT1nDNymm9mETjJ+q3XbKL+YSr4lgMmonsFjU
QSkoW/Co95v4JWnUwOTpXfeDjQdLa2MD+F187tl5fue5xW4VdS+mDqqeRTc1NOrUNHphL07NAhbS
JAr+7ny0F6vD9Mgcqd8sI+lFC0gb3WvNXywVf8GQnLQkoSHF+Svi2c0H6jWWroT/vsVEH2xG9V1d
yBbpQcZ6W2dnK9hQhbrwbKbEyyCumzLVQnnkbDyyudds6R8ac19Omm3yPrElpj1cckJirwbYDj8y
Ht6hlOlt2L8cSTgpJDRFKDrn+KaKuFHUtf037QMUZPpC9TwunSoT2HKw/IpBHCjszUTudufIeybC
srMR1hmRVlbHGnJPWOcdRnpzAqfhJa6rdbjdnoOhsHrzMT1pvU33WX1224RBdsg+E4H5+BW5q5XY
5senE2FQT2WgYM4ApSoo2/bKVFQV8Mb1Z/vIt0gos1oeVbDok6+vWBxyy5ZmcePbWvUyD4Zh9rOO
WiZo0gkIa3/OB7Xp1M2p2/XuWojwxLMxbtu2C4DAD7fJ6wI9aRnYFVteJ1HyTJ4H5vsU/8QnQ4ne
nc7oWvHYGS6La3ge86210WlzhD70M5nWXxnTS3EhP8ONiAtVyp3Bk3SZd5/eSW2dEWFRM8a/9Ho1
XCqDO8FCUBvPHNBNghVrk0D8BcOJ0X3QD+vveflk13AlD0+HJTVcYToUfbfQh4G2Mjt2Lanz/Mn9
deTCY6RAzSNS4DolALACC7g0vCHSjvaF7/qdPlBdamBLGl4g1dxBVfLZF95oEEtsJBi8W1ceUecM
PxS8pOOCSoOAjYnwZ0C/CDxOFEF2SaAZ78uL/kIgLzFKXY8YhTeQq1fAUEt2I2AOJ8DWWIpINoxX
6vQtiw9Dd5V/uuwfTVMPmRPrDTPVXyklbHE13quw32uLgiC3BOh4gXO8gKKB1uIxBi0asJ5D6qSU
dtJ+7+29HMpZy0B1YmRA8LleZEEWy+25rjpd9HnSmXw7HtN1Trp0SpjmKVn3kRR8VqEft5E/THFS
A096C0JQemjHvCRY9ShJNw3du4gmgIT9/U3NUVz5j2QJAB15/szIRQz0AkuXKeS7ezLaZQ1msGO4
oZFcANKFkWobh1I3RWniVM3d2uxVNiZTDzBXka8nn15MVjRlq8DACE1Zpdr1uwNUEOw+wGNjwHZY
/knRXTS7P2IdbLELRkRZ+kEn61r/qw3ZKe2d7lza3pdulBnMzwx287LfC8kJ4JzH7+dCl0zT6Oau
NdiVDTg/1GPImgHMfgfkgcI+TyUZlbamCc+zcdajECZ+9Ts9Y9cC5TZLUMX/IUgLSZpWdE+XvFrZ
yoKMgRZVjnIG+lWSXROLMJT1zuiPlAcpRahw8jwrqvMETO84YMTxCbb+mtjUiuBDPcu82XbWmIeV
X1KXzzh2IJPhE/SUe8jI0pDGtcBYN9EAMVnxAFEeUDD3eBrndzuHEb28MyatN2Va5I6h8/hroSJl
8ogi8Xxu5ysvkhxeDVfW66EjNtAnPwLYxNf1LcmhcvWUYxCQMq3x3sxL2wy20XQ/uwDkuxtbLs7t
ynaPNkKhNfIIL/A67syIakGgDSEaEaLcSLlKu91q7WYoehax18/2frc5Tguehvf6ZSijGg06ZTgM
F9If8QJ2Y0UtjUgV27li4LeVCnWA609pSuMH+jbN0+wdv0fLYXt8nB7GeUulL37MTWwOAMJtLvMH
o3nCbMSryURoWxu7k4J1BJuFrL/fOdmQayHT7zgz+Rn9Q9g9y6dMqDtSBBVi92X+KSFaWMX8ZKFt
1vtajh7eCCoiQWwblJtx9jQ6MVV7hLgM8WxSEVbQ83YWTqjknMSd5Jd87wlyqleupYy+mjMGXeIj
51HCaWwu7jrICN6L1MTRpk/eh1EkEk3Ub2K8Nc/zTATd8WjCpciBVizwYMkiDKESCKCRzYY1vHNE
y0b1wzbMS3NC9MdLgPRQQJZBUZIAvJUsVWykqVIolM1q56aX0Uvr/Vc4Ai7PeFcPIL3Gbe7AzKho
X/FS9ZM1V+ThqDZKiI8UrZqgCCM7cTzpckU8rk6UDpjS6jNpNeYbvE50FNcTgLU0kePW584ED1xR
vK4r0VGxc1K7flBjcjGnIUfn66QFFRDj4abHpK0cUQoaj98oFdhb5Md7mT6ATzb0ITNr3KgmkfXy
iplRRI/lGAgIfRQSjaKQqgSacunEq6rI19RaTKKgPGqvPBhAgLqeff9q0+3R7Ud6V/CM2a3+35K5
JxPvIIZuO8AxdmSE0vIRkrNUFHWXZK6e/1Jd/+by+1OfDMjrjoDxHAwU0TVjg0GWjgGjuPgvdyVd
cK0i2LDsgfBm/V1cj2/xDi8vSFYWeMKh/1dFWpPOlGr0D7fVuSaZMGrppwOpGOt1umzSBqKOXDe/
VPcVUAtkACfl7wohvySnbTcDiIKn0b4vVHGiE9laAhLzZkUdgLnybFvZ2KLU/SQ4+pCCZCRvErZU
R4/TosP7jLB0f2oumVadd0mhNm2L/0bgc7T4N5N7Nz9zf44lnNfI+gevVKlkDqc21rxDb8STugWE
y7dSXddq7+/tAMMiE33Uquq11pggGjMAUjEsDcnix9SLOrroi/gZsplcNflnRdtrqfdmZdDuBLZr
QieLfRKxS00osLRG6tMfc+dMXow310TIMg6slWDJitSxLBUQHRmbtLYE8l/7jrliSDtTntdpjFbs
RKXAhARtSmLr39fJ4GK0FaeTBrelgC3eRn2qc62zxzc7xXZ3l5HFi1lzMCydLWetsfew1lOTX/4c
KEZFcHyfsxGpCNTcUMsiBRP09SgA2fMgHsatqJToJwl97WxpW0kEmS+tuKfwwz6bmYgZJvXEIlYP
Td/R6+P1MuJxelG9+bXOMiDaEdp/KxDU2rtKRlUg1Z2gy3SwE+0P8+a94FveHVcgbjY0tzNRxqNm
APLAJHy3vW8eHszQVyNHXqJtx13EREQLMVD/U4SiCmKysgA8yFYm0iD9TYxG6AzP4hodifMh1YNS
87g3NJSQhM3iQdCq0451VW0IKhQn52SA7p+iOnUPNZ6PGmixxpLjF3a3KcwNsHielUITtGu9hy6B
u4Ql4cmUZJbZp+UIiw2nUIWQa57Ft+VWsSifiz5ZRMbUMzOjxohzL8B9PHgrlEUU5uek4E2yhUh6
5tX6wGyMo5J6pXc6qFQE+ZwQcOMM/05C+8/39fE8bVIjspHlJPoQx2UQ7JzIRlvBZQrozLHNue0d
D4K6vPVsGH2s4j3vc/eNyTP06lvf8CXPjxAjrFouUYRt8CErfQwvbnnkPGJMGK7DjQ4gxOlfgBSo
yUrDfHEfcQ2uSX/zCjzPJ69fv80slxOnWCRB0a+7in7KCqCzlS1jz+SOfP5tNvRDyfdSThXmRcFa
vEuiK8Rg3difJkETnxbZvblA3mYa5ayYcu6niu3jU3xHquBMyZwbwZj2UIK97rnVYpk4KIFHcdsd
WTvDuOrjN6DbWtzB9DykuLRN3J8TtYTUn7ELctgaR3B7AwCxH9Ll0/k+zdlj1iJ9aIXpafJfDDFY
SMXmSe0TNi2Ty1no9YxBIX3lBAsVTn+90XIFQHMeYYpyhDpVEeKSSGBQPiQk1SMnxOadrXvHebGJ
NSo5F5GYXrW/y4GkDAFLN25zIT8rcZsIKvAM54bbDEffKdnPBZVmnjF3nk/e1wIWHGh/9kOf3Gwe
TFnl1jOi6FV0KagM0xHuyWrELhpco7JckYXwQQC+6Q0IO8Z3ViMGv5IVYDbkLUHMYpDtRRld5scx
OTP1gSVtxXyuX0zB+dTal3PUaQT2UiKi8DmZ6iPlg6PmL9zCeDkhtQnw57mCEYSCVkUSKQnVnMQc
hSJq3YJqx5q4zP/YcMVtS3LtG70RgZS/PyX/lOMNwR2UmtJm1zXCwIQGoB5tXjwvSuH8sYwgOwOx
fCjigUwvpfO9wZJAnyJTXMjyF8/+oJs2XCfeeyJVX1Izzqe64Rd07N6AeIkA4pgOXwhHcVwpZy2h
XHoIywRMwE/pkxkl+6sHxqsDBJ8/rhWEqzBlrASVYwiitpFEL73yJ4H3OWAPMgngcIZGwEp0OHRh
m9I+Ov8FCL2nAjh3HcY7eupukODpqB8jkhJa3Jdv75gJWLFoowK6Wv5y7zTZ3PhXR/QzBk5Uiz4Z
HBOpwbvAlvBHsrLSR8Q3iZvt0+UM1+0WhoxOvgqPfInrlwCm4O+9mRXzq7Ht3J6971Bga4S60DKf
xjho58HoIxOjhKDvzrv3MRLSpz93S44GsTHf9M0T/3SgU9KUS3tt8QwhKpzgFr9r63OqipftDEEz
YKSUbrBkrOVKuc+MRTmMpvhhL6sS5JunURDHmVnR/DIwdo/5Acr5HwmRbmcQHxMIwFqjhP35CZwp
bdcwrEj2c6mQX4E3gQQtnKC3hwXKNUJcb6hRvOSUSbx5LITxXsIVboclQDJouk1S4y2/44WVXjJi
8d13G41mMd7oYXv/eRvyu0hkzZih11JFAGsJn64xWHILXiDQkDSidowNaoCZ2SFlh+ZxtZHbyYsE
yAUi/lyU92i9m+3cNK6gTo3dDhfysDw3ypz0UPvk9stxEdKTXFLaA8iOIwWkXwR+R4kUVg8DsesN
Xrh6W8n1kRr7Y50BwCiek4Xn8SiiZ0gLRUxsI3btxTWlldtp0y1IkWRiw8h4d/t6a6iu+2uXZnXx
58Voyi4Rv1ULwq1oO8Eoqvnn/DFWMm3eB3nsK1Mftz5GdKIP9YzqbwXJ7DsBjTHFRLB7bOeOrbKz
EFrc4/+rh5W/STXkWpTgjSNuROk4ncem3TPixokc//oitCmURmUB5eWKEgTMtbQ5VXzgHCMzcCcr
nZ/uTatWlECzftk5WfdO7H2TjwJUO1M8beGEDrvdLjhQyGhzs+ofm61RKbCP42DzXpCbdWg9DAmG
f8UzeSERCwoGaqXAO8pJ4Ytjeh1MXcxO3RQouIrK2rRk45UySduaRHxI11sQhQ2dwmAv0/lt/td9
W07AOPmH/82ruQUlhKLBx1mu4c53/Kgdleih/mnQ5zQ/COgluHSEUgKOYJQu9UjQ7K6Ral6oCkJ6
norWeogvLk8vnNnXmZtI1f1L7zAKzXObatXCUHtHwOweOke8WA9OGYEv8llJQ5NdsZvU4dhHX/f1
njYLdZ7SIsCb2o06QCiDC5W9AaZ5vvwoOa8SZ+bb5a1eGua6wG2Npki9+TCpF601VjKb53NmsA0F
4/Q3qsOixNxV83SRpQgFgNi+FP7bKo0GM79Ru8OAIjIjLqv2gIC4PlNWpAxTHovyqTmcMsiXVyK6
5qRrOB2hDdbzaAWEncPxgQa0puw8+/ZaMgoswp71P2CgpFckEaDA78ijiJVO1YpyrgqfsHKct9mI
Eiu762z9+K0X40YNC2AYvunkAkHLxje5Yey0jjyvUxfYQ5UqAnujqymoN119yrL/LdmZmV7OHkjK
+bGp8dJAr2GGnsRj+7H+RdUnQjwoHGv/G2lK6Wn5dFB4ewwkfmsIus+1DbkbHQqFaNFtlXE0HSx/
k7nORrad5VVjXYGkyaZD85LDl6pfXcuBHy/Ht9GphcCmlg/bht+azzfKRCvDkZPHbxovLaV2ny8W
s2sC8Yu/g4KG7o24g8r0eEljiZ+Bg5KZPN7P3gzylZDRLandeIO2MoH/kxp7kSlcIAKomVUY6IH8
34ZkJ9coKpc7E1w37XZ3ET7wR0se4GhrBcdq+GzgNBUMWsq05+lC2Bgdoqjr0QQYY374dQ2QZib+
AcGRMZDxsUKPwtJNgynyLk1w0HWOtqFhzyJjVtPylvE4ttKC/qnSIhmFsssIvcuWSwuUOVDPtbHo
prBVrlAfH08jTy98dVMpiU+JuPVXMj5nc0Rv4GODj/AwiqRtEIOPvCicGctV2rGG1R1F/nnPBmhv
k6Wc4E7ZJUbjA6Q65+156NTtYL3w3l1nGcdJi/wG3B8hK0865J6jLDDB31gOJWpyjnXQWON3Xzec
xmq2auEfLOxRh9fqFYTxtqH/4LP1s7oHdJJ/i90ky0aMaeIAhG12Ex7slXnDdy+yVIxbDbLIfFMR
AMZa4oU0FKm2CRNxa+dGOJESMtquNPwSA365m2YwLDMBiReFJEdazGutR2+QTHM8540FRQXHo21x
dBragZf1FJQJnTn+sH+O1rdEH/OJFlRt0Y4VSLGfcBnlGlDR+HTUTNzLwf6VSLqtR+yc4CGHd+VJ
Ql8zlCutVfFxq1fpwzaICawWENmtGK9rnSxscSshNo8MKuHV+Wm81nahhmuMJ0VX3acRtvWqVreC
WD0Y3VCXxwiXxMLbPg+jGhKxMLp673M3OIVjkhOeOQ9CA4E2p+pvmvcJK2Sa3rLPHml9r3a0UXlJ
CtViN4NsWH5cc9SWejU7kCBa8J6gX48ZlPdxDUCtgQPMIUQ3HRghm7A7g/gYxYWg5TX5l5Uog6ci
By9AJ9TFXEBsnvdqpQTErFIfdv2B2WmathKeJps8mVPhgkulMzAf0squ7Bx5O6SGIN4+UH+ZOt1H
zPjEhJBeM0mEINb3RbYF3/yRtPaHFAYSvHUid5GERYRtO78CKGko62DC4lGEysCacZHtoDEI8aZ4
Fi4PswRYZJntIv+mHSw+buRmb73i/fhtnWT85WKCJ+aKoqvbwaEHmGc0fDNb+uv5awumfiTFoVnu
kdImiCPevKIySt2DpyQQKcEHWj5TXtX3OtshQivD5nPkWMgzPHOWLJ8Yzgi014qVV6kNmXNNY//l
tK+Mc8N8FsY+S9a6vvRRJN9M2UKUlHLt8GcZPftY4sEvu47aF95n8HpY2sdTwayv0+0TKAnsbeoc
YPjby5TzCxD2R59WbxzBJcTOcjg2oRr0ZowScUx2FWclY7mO+wXeQZzSkunwSIyb8qf3mXWjwx+K
GlfEnjRFKcnSoz8RR8iZ6fr4F7jUr+zw+w3iooIdcQGGHBEwGHkXLA9vtV81RHU+P/YZrWIOI6yh
IH7Az45nV2dsxPgIXmUM7HLa8T4sCgqILkLDtTD9WYykkXdA5md4TCprZWNtcgQCUIRePxMjOP71
S55Mj0aUldNVV0FqEILclfFW3S3RP8Za+Bf1CAJqrhHhTL9/GrZEWL1cp+YX+oNfOHgjrSq216l7
3xKmSajYSAKS5U/7bEfiFb8hAIHMsiLoWpgSMa0KcrkCWgdSh8RHrV9n2Flh95AJk62f1Lp1ZfiD
0Ag/H1CBvhuHFWUdehjZU3iZa1AQzXbnD6AKF3Gbvm04PUeURQy7sVgun6Sar5g4ZCD+azZl+h/n
ZjjLFrI9CYCpA7Aw0FLnR78Bi5uRu2d5EAXAwuAMJ5jhwD3aQvaCr/vxCwIVlaS/w+l8vIqyxAI3
RXbpJRS1f9reC3tYCd76/Kc6YLO54wtpDdBDYtzdx+QvZiKDeBmTFp5WpnbRlE1V3MXYNdVLJo1B
xKUlu/81c5pZBWncW1E/qCCv8yR5Ka/W/uxnPKF0V4+6C0e68Y90F4grZbCjmShRkMxIw8qrfIIz
gHdsQYzuYpNcwkLICHTI27jjY3MaAA13CxJmFqr9PD8/qsZ4cH+CZVGRzL4QBSqoRicAr2g5rA+e
trPRRJ4wY0fuYNLD+6QOjBF7q4I/k72hcA71zSo9GBxvZrPbHytmGM1Erl2YjGQbmIrMQCHY5L+N
qyjIM1h8Olh0EF96lyoR3FFdj+0IYvffa52BIzJToUN8uqO3gpjpE8cOca/b0+uacMVeooL4+8h7
zZHmodcqSfJvA0MDYMd9HNh3LVWagLHwaWkYdNDaD8sJAaV4SWTzsczpoHMi2zEvL6Zz5hqu9SZO
gyxKdGpXbSrUYOOzX1UDmTYPxg0X4gi+hAJRkBN+aRm4XVb2RLRt/PrJ7GVoorHC20XCpIC+POHm
smTj8smArJLxo/OfOhb3708XYr8KiI0j3ISOJYTKtKLmoHXBt8HszfFtf/9/F5T0oFjIEzxvBAWI
PuKuEXWogeajl3Of6AvCVENhdLR64O/N0MunYrv+egrhvPqMvqpMQxS1k6VEyyKmCb+Zy1MLmuqx
DtpelzU3ZwxXatmMXLh+iC6d1kkDr1Zo326X1zNtubO985yQQi3MckLQHPj77E7KXGQ/kYZp5DXy
eTop8k1zSNqRyL0W+mY/xZ07SuepfMO7moe9+OHfdm8YYLP+nwvZEFYF4RRGdwGmbRV3MjdneSZX
elYwT/RuvUdM5ojRGW9im3PTl5RRirjwURBn2oC+l1TNsvMNdaxF1nUS98QxvhYeAepx5wKJ3M/d
lMCEUFZxscZEWGI8s9zMQ3DViXcldLbPJ6fyqo9NBDprD+kyr/dnQDx/+cwBrwC3BBgC7INmQHyR
xZ5Isu1El7rozWxJ9iF0yYo067Wjv/c4T2XqHOhS1y0SzfNUdS4cQARg+A6LVK8mJhH7wNMpBFLX
GzIR5pgBAODxuzYq6tWr/uVYp3ubSohwGr5k7DG+oD2XIMBOM4q5IyXfCqSgKeO7bkxLReYPqQNV
I+hpnHZrl2Vc88NvEZAMgsSTnQs2gcwf5XbMVJGCnywx+mwC6TYDfzIyWXAq+r0Mkbi4G0f8lr/m
K9krvuAGPdghmFAfHqsHEiilP7kTuUMQHp3xj0o/Lv7ZhHd7U/xunWFlVZrcJaSdeF7iM80Rcnil
cdcquyM+17tcZDQ7/yK2vn/OK6xZy/Ftzk14Eyag9OD/VlV/8wzBOovY3l4w93WTF3vooZ8n1679
l6hHjxafzvIglMknamb+a22tU4JT2rqw1dfBXMhSvdt+KZzQItX79a70jxyn6vaVTwCqdceXnfVx
eq6aryd086oukOZUE5Px/OrOJUQ4myL/AAEd+EbjHiOVJPa+s6ebL7nH8WRv5XQ5q3gSUTrcOeO9
OHaDj0yjExR9QQlNONVrk9DHKxF41c9Z8OSwNuxqZnuxkpGcgQLlhfJrXwKIkL1XAnJ3HcdYKYhO
KYgOZegOiMJXxusJd7vAsdt68LpdF9cTYl9pop+rs72RLVYiqVJ5tMfzcWYxYP5juyrw9pFtcIZX
uI29xxRvofuhhMc/FL1so3GSWz8bK6B/ZlH3/J4pqR992LT7gUczMPAmQjaTuvILpcK2PduPINDk
GUvOCS7rEAUOsTyGCFkTzRzWw2wKVRY38X9yUyxvm9MvH49bQAZckFn95fXnyWGzpFL+8jL7ewg3
x2cLKr2cDatzbWHYJfOmpFK07EKt43AvsuSFboj0bs9+GfU80aRbvk7EdUmU+OC4KkZeazHnGkuW
LYyPOiMzzX6BC0MXaF0lQR6lG4Kv4Ewd13rs2KXHdWFZBin1ksYwxGiJrDLqygEw6U/SagT68OS1
DABTB6IlHOYRx5K4QgZxZbRFQHkxpMCaQwdg6bnfufP2x+5XE9p6s/J3ckSt6dG+aJEX8P9jBJ5U
tJFX425KyWz2w37uTnFOiB8DeZjGrCAB9fjUIlmyxxD+DRbokaYRYKwEcO4z6EkdxbIuBUzsWhjf
MY8dEcK34hzI0Ok6sesaBCvTCfEZTox3bkqM+xOQgE8Cb8UuAxudcqTb0m7a2zeFE4wQbubB4J1j
8e51+kSfxv2TrS4ExVgj5fewahUQr6lIEvB7DFi5gXqPQrybdyoEPDa/rQ7MV4gj36AVroaOiAL7
+QwHfNy9j8q7Oz53q9aEKdY//YnOArPpP0Bw8wSNLTx2UtTmeK8k6V7T+EW+7W6EoXTkp5HIEW1t
q6Yz+8W/HEZIAfEXZ1atz+V1ex7Y6dG+6MqwDpssDhqHd/97s997TZOTY7nGmQTX+/GIGAKmivXG
g4fjMrhDCQR0y6CNTq/Vohx8vzAuVtGr+cOpwF2ypwNnqJUEzx0bvsXP2h+C2wxfWtmhcuQ9FSQR
McfcvolRhefZ/ziu4shZ1kKlLN1QrEDl6nN4lfeNG4BXk8f1leVxFptFFDRULP7oQADmjFFB1MHJ
jxweIXErsf4jwK/P5k3IarbkFqyU+T4BMxMCTGMjUZpp23i/1+qAxxKYJ622dQZXbrliYQMRcpJx
zfYXSSkHjAQ6swg+/++rv6y7RdGALG2+WvAidrKl3/FjAKWvQ9VuTpMDGG+zXMORgBIYh9DAhpjs
Ct1ZzGOCaRMPbSYHh/6mBiICgVW30MIpMJycwglk51CEP/PMg/rb3MVEe2i2PNwGnffC5/DZBpVE
Aud4XvCIQmykSzYb1CVxbLvt9fFSh01B2DxFJuJ9k4aRv2uh5EDwIKTLUEj5+8yBcTxMXTo6uEF1
Q4J0tTXH4To337bcHxlOWqCyZv6KfLI5O9Nfn5AasMslmc38PtrQ9ESkSDtTeFlxjYHg4ym8DSIm
+16v19NxUxnBM5JoFyh0HOpo4wDftW/b8O0C5Y2gUvQiFa+hjob/08qpPhRFeaaEBeg6Gd+z5bhk
nA9rde5sLQUdLqODncdZkkFqgg6FNUJeZ8EUqKOicj6CRqM3oZVJagYrpM3gX5ezVthXYEBVFvHZ
D8nc7SCuwvfLNNn1YSmAOH9ya5yLGuhTlvVAr+p/6DcTi6TJcLhnFEZEnr6Ha0keHO1H0VQbvlO3
Tl5h6m+BGjKrPUIz/xcx95WNdtjTzgpGIDPuR4ciDFwjxgTDj1fF5hzyMghpOyMIs7WNK5/VB3ni
l5L2bEIeMFZxEroYp/MgYfKPYsWq8z/f6ebdtX3T2M5rHatf/pHY4z8XG5aPIAmfWIyJI+/FztRg
dGSe8tzNGPsUT3uQUDxLMS3eS7wWbLwZ4dVqDqgp5bkUcdMPaPyrwV5QAyKhcgqalTDO3V3hSxhp
kEMKXPFSi3JJl0S+IoFNgm9js9S9Hc9pY7Z4BqyzqGen83FpxczwBG7vibgYiZEah4cuoaVwkUSL
Cdd+YIjnJgDANe0HMBzh1YpnmjR1KyM08voOB1hmgWZH/gxF+U9xQxPQKYFYKwnSW7IZ8i0xk1+u
eQSL+DudlypI79cpxOI5KLm3RFDP8xJeVuUPfB0PDBli2SWINvPah4AlXi665Sq5Wb103bwWsMkZ
XCS//ns5RLrRKQ/VMcnVm3vcuAltpwwQFr/w9+tKsm5nwF75g6quMtBS65eCvGFdWuzh3d3+R9UA
NyoLvZ9W8OpeZVo/GNp0YjL2zTE3GlIROqgiwfpqdaMyvSjsJUXT+iBe6WVEN29yAcvFFKMYID1J
MQr+oLGJDRmN6QgtwBjDZDsXhdsoTJgXYXe97vZA6NslrIg4XprRs7vZfUlxauR6AL9DnEg8cDoB
ShiUIH+dqjk3nX7HfHiD3HHBJquhT8HreQurAIMVUxWjhNygU8WmJxYnpNqbSTwLu0grTSTF8WMa
9jU/6UNh7amrBWggwqyJBYi4M9hwBsbFy5wx9o+WO+ChGsM/UVNNrKD7G57YSmLTu7x05jCDFQ7b
qKuX6mJ1yJ5r7FFtdLc61hcdWk4c+scM+knGGRRs/5CAwlnFggbJ7KDX11ApGL9+ddnENbc+ERLu
lspeByGssFQdgwO3ECozofyMx1Ai8xYlxDIobWN9F3iYdxlFP96hQq9lzQT7vgA1qD6blUfhXpgB
W5lolLwP6X6LJqA9IqRatgDKvBQXX+ld2pvoblGDQcAeRMZfuByvZoaz1N9PgkM0qPkB2gkjKWF2
/fPP/MR8MYm8qSqRmAMk4XhhsxR9Na+7ACGVqRhtSHuctejkBkVjD49TT6025SyXtN/YtXPC6G3y
Baj96AWx5HSFraR6PyZVsYqQy1LFP9mnFvmllSmuRKgCVqulv6JDWzL1Zzy8HKuIiLdbGyQd9L33
tGytpQsuI/MN2+wwGajaDM/TL0Riebyl35Hxas5Cg83jQc2BnkArrOIjAeSwkMDL2cxAbGRT6DVI
gMXUdiLO7m27XWMBH0rc425h4sGdX+uDdx70k6k9WRckohiGWmwrOZIY0YG15lWXixf6087o169x
h14H5LnFOrNpKCzdBHRHNRvel49GGsrZdeqzvfcRqBMSFKfQG64QB1PLDem9+8GJs7apLy/Qs1n+
xCYf+gwKxLe3p7ZOFDAX+CSdj5sJUS7dAfGCKs2SpkJdAXrnkoDn+4Fhb4HfnXSwcGJNWTVimjsP
0JjDGl2L937RQ0D5J3vDkmgU+D+N9lAlPA5J3hBpALuSPZi8mqQ/bpc8a3Q+H2FkrXO2SQQR4ZTs
vN//tY7Zh2XyiCREUneYhpcDH9r0GyS+6G/VSQKChrZCZoOuPLC2WmIk167Hi4ODj4Am+IwuWV8m
U3o2iqVuQa3eb7pRTyryU8PCERiO0CFgy7cjJGXiIi67mkCzn1LQH0P2NIZKCO01Zv/ZV9NwRhC3
W34FEpWB9nnhm1zki7l/8GY8o2Rc+HSDYl9B7j0dfbuT4GWgR2NhQueoxCBjNSDNB3CJ/xo+34gQ
DMpL4tLFnqUPhfWyixvMG/Dk4wAzesBKu6zrMFe3lx/9b1UZJpNhBFYu+xwOVfBoh+TEu9S2BFzm
KtTiph3nMX0HC9lKK3rex4BfEvlcfzRl8tIX0zcUTTsu2qJg3xiDuXPUALbLScjmvz3DiXFraOmd
bAUKrPgSLdxzkxlUks8vOWPXMq8ha+9+AjdEG9qzSfh28ObkIt4XYt07uWki1Ri/6tyLuZkOxntS
uyFsSiYgbsw511+4Je93iXGtSsTOaSbrjHIDVcj258b4COnXSSU7/XqbhVCJW2IgJcs8ftorJAK8
pW5cQcMJFu5pxqkkciMl1yQhQecHmFz5yHwbF61quC6sb2CzD+OWSWS8c69cY818vKum4qttUNTi
axko46J6hRRu7Z4GRkRGgaltxXXmsXqUC4VlhBCD6YdMF8hC98nwqQez84Wmfkcps0ljnFW1kYMf
Wkh2fh9RZqeu04eoZi0nfTn1H85iSXEwR0NHNSKhewQsb4LYiY76LlgvXAFWpklRHX19oJ6vrdWE
5EZnUBug29K/THSVeJdzmCbESLHrluyFi2aeOK24cGDd1ayIuwDeoPK8cJ2xb2qADG+qPHgLKDPS
54M+y5wBiZ74ywat87dVWg/FwDib1dLMbUH3Q48WTeqya5Etot+iHFQR08l7u6fiEFnWsu/tFoB1
7T5CTdesO7gXMxzH6I5tE84t93ge+4N8Iw7VOXxpWk1VQSHB1E8ce/5p679ipHObmofMJ9LK88PE
3h512c9+8KPA3k6viXPa2l57jTplyuHLnm/xZc/Vv/W7NaX9CzJf+AgKEEZ+5vzshwMcvrCzUEWS
jvibVZpFWpgHbcd/BFq3L4nNB2IVkEb4cecePyoVTWjQ64PZDeT7xa35hCF0a0BsfsajwPWhY4wU
dlRKY6AIp4nmdz92OoKh2yx5nOJTKXxuBULAMBv46MDJhWtmBiPufRt8SfPwwZamefQ+cqweJgpz
x4Vj8zV1lcH1R4Qgea2fyhTHQHfDnHw15m37udH+Q0Pt3KDYr187faUNLhXS6/ekFOs9AoC8bMRe
8vthhsjUkop+P2FbewKgdkI/nfvELm4nhXeUcqUo+wWyJt60Vbwjclb6mpgJIpUHR9OHs44EN1eG
ONnd67PbAHpbIl5OO8s/DvUK+CjB6xcbUhEL0Dr8aSXXDMIhQ7xA2nRW59zECrg4DRQtEuV+g3t9
g/Yuhmo1jrq0uzILtvrnPfaaFUisxRrBT5eDhcvg7cmtBCJEFrlDYyPLvRrcm/C/K2U10J23zGHi
i30QCd1SLh0jbDRvLVC2qkEDuHDoHRzEFyHrCHnPN2u3RxxshC+gZuJ9dTxcJ78ncIMmYU/vvOSe
pHajsbnxbnQRH9g5ZwAsW0Wq86pvS7qliHnbomgzIpJrsXHYClgfMPk6KPg4aFb4uFoC9klpEJPR
kL0pthiCycbNtn49K9Gg9hYJyrm4iilBXUPr/WKwbA+hMOP/kQMojrbx5Pt5Dmf90jhj8cqJsHCG
bFU5fBTSaLe9882xhE6bFVVQE5CakmYx4StACPTIZ0VCoefOJ+b1g9uqkLKmZscC87CxBlkGDDG7
Puo1nhZCpgcxPOlp+gWIPUpxa+dhKFws1UdDQNhPDHrKCva3QFetC/bu3RAiN+Xe1bqT8/czHNC9
+GRb3BcptzeuAj/fBcj4fKJFVGkn6AHerYBEAG4JPDlHzJizvQk/zuLIvrMxVQNFvUNBhSNR1rBI
a/ePh2FIk0ni0nI3151VlS38Lald1rnWhj+6Gp595H9DAHvak4Pbymr0JefdKzMg8ZN048uCBddj
fp//Zj8JuSiRW3euVS2CirMJ98O7RRcPkZT7OcLKbnxhE2aMRWJz2VbYLj8NzxQmSwuT9/rMgahj
5ggqBARVRoLpmJTlUvTSKyKOcb8KII3fjdQueNVaNvizXGL9qY1qujn6VHWjk2oGhcUdL1ZOGLGI
ALDYj78vT5McJut1AdSsXDHUDFJo0Rd3m8WQsLa+xqgKLP5gkPtFYdtUOElLSUF2YJQSQ+TVulZl
CgtODnOAx99LmLBM4wJwb1hpbV4QdnaKi6ZZaKqAIytwYy1SrDeRCJAwYjiP5kPxSmhv8H6txw8x
iC3ngCI2yMh0jixXb80dlz1ivFtq//mJ2PE/Q83/AHSvN8dc8dbXFQCMt4PwCUzE7fjCdhj9QZeY
/MNf7hlGfmMVOi48lkxbEEMfjXJWEXK4kM1P1w0Sp2+cQdEtEgtZPsPSC2X12YdYXAsVx4jBg7aX
8MqHdXke7rtamRKvvukqQKYVkY4J8RwaCsmrxQ97M+br6BSg3glmMLKKDvIEcgDLD+VSf3J1+3JX
2rblNPXbZe85wg2YsfVhlpz6pxHUMRkHIW/HFzm/d0tssuJyVzwdZJucjx0zP/Jxyo8eIVWCBaUg
J5psASzNuL+xJIqV4U3nNTJjzIdXorcX+aFPXK3bMkXoRdBQLEtyTfXkpZNRjbiz+/KCCdw+fR+5
UDdHS/rB87o+u9dOBEJ96r9KUh1ns6+eLP19FHjz2+Xp9n6q1kfIiwoHN7/OJ62iKyT1xK6q/F7r
eWzfJ6FOV/E88ZUTxxKYNZK/Lsb65ZxhimOGnHeXSO+XowrUorNxtCbQ/Iv2FperIeCCuC/p5EKT
AqiQITW0R6FcyQnYmeLy+SAiAs5o0G7uWVFxhFiWjhA2aPlOLC5PBzJ1aKdHegZnoDw8CY22m6dk
fUZOmbn2k6TtqVd0zRKjkX5u7bCsPZs3xTCZaUqlzhvDpmks+9jRZVjTauPrEE1Ay8hTsz5VBIyD
uyq4ggDc4wDg/AkvXi2SHBbgu1NdXyU8K4o/6HRI6RCfevk3W+0455PSb4UcSViTUhbGcUUgLXvI
rapGDs2iqlDDg/68GYb0FwRrOXZq2e9ENCkiTAWjFvpXrUxLgGc5BEPEbA/s4JYK2YP1TDp92qqk
aWW8xarNzQqIoFO67D+i/0RM6A2IlFC083ne+gkRrb+mQLwE/59vSSi1sGlYoKmDo6DVau8gZGRN
zMPna0wUcW7Q38mQnzkLEFhy8OtbHLBfIUjOuxpy09oNGOS4vDRVQbkY7E+0rpU7YVlFHdhlg7hi
h1GwZU9nB1vyrLgR8SgPRhqtrCqJlX0nHwHv0EhKpF20BxsK15HnZJ+qDjqp/y0YMys/V1c6+Ovy
c8bMaRbG9N2aSVgE8Puz2jmwzRuWgsQrrwqD6ApQRGlPd1CG/m/fxxqVhxNiqlw6QKzY/h6i2asm
+brpOnhoRVhtQSQEO3y0r9CC4QrUf2O1Qh6J7/t1t3CgUZ7cOU7FmMMxnPZRBZ5L7Clm25mYajFh
jgEchpcEBT34rlxBbca8F6KLrDFRWzodUU4BfMtqDXVAqAzHUx6OtvYTE4H+lsRvQ2s5Ps3OWUnE
9gOisG/YxnQv6UsXynmE8iVBS/rb3BnrAnd/0HJtRGkGmGeZQNh6bMf7/T3fsuZf0ge1/YkuBQnx
ZJHF3jx02W3e/m977fSUG2tL+31xikwfZJudtUw5QnLa0Evu+K+hcPr5j17nL8KrEjs7PAMOJktU
TNCFH6LlV8BblkTuMG6Ezmv3/bKrCSFN5m4LFBAOAppF+yYRNZOkHBPWqTosbc5OLaC+Es79+uVL
1A8l+Ay9jCvuORJvCakDQmgpmoEUaIGIk48N22sWdov6kx3OP1MnbCSjbln+/BZbuSI5d9VSIDLK
6xtVkfcQejuiXvulDu4w9F1hWYLi6DD4HKxj+3062afFTdKmHCnl7Ic/GzvkeGAnf+9eNZ1tkb8o
1t1G48yrBSOpeLF6718GSfbKMdo1KYIQR+n3xMcqelrz8ifd/kbiNd0zQEibHDIe1ffIaHviDpEb
wXb2eoNkU+LSmJuwU5zCrr+s12hAbcV6veLhwH9Lp1VPY5i1s1lts9cOpYcIyNYuMqOQEPyR/wG2
8L2k/0+9nTBTsO5e+MUXYcJAAocCKjN3afci4D2eVfwus1uXAACzfz9a3qQMDm7mKPtw5Qku2+5i
Pa0b8sBZdOEfYecthFPfxtPehRHyJoEeRvxFNiAJkqIWGw4hE/j0uAKcEpqOZ93elzaFFVZKBKZb
wNM/Ee4uxgCBkICE4E/mHiiOefqHoM3IhAn5w7qNwahndAmECaw8HScp5UctGFg8H2u+K0iJEaO1
V6fzHdpVdVwNJ4sM8HvNTLqKolL95W1bJS1xdQkTERTCgJJYpBsQjaSbbmaEY5nSxR7T60xaetQV
7cVUySS15d89PzqcdgE6xKVBQd8F1hCWkCh2AvIFvsWDqTyhUBSEx0j+IGY3Mu1Kmk8mn+QOBk6l
pa4GzMBjUb0Mfc2VAJ8vlkt0xC/QfC3/oSq7ULvtowXtJzpisN+ok9SgfvPSF69v69JThkr1KAxy
BoWzJPr2D2Ct015NWay9UzU6OuKEB2u/vs+nPSem2bXmqSVWNQ1wfjkG090+p1OnJ6DKm9NhYl2a
Zz9G6DvfO5qY2d5ts91/7hQG45YS0iKwdaZHTx+auij8MYoP69JwiMhbVvGBku1hbdUZRadAmbag
bU+7EFBKoqFzQ3SCVXCIV03t5P7oEdoPe9iBiWMkJ89+o41CgPMNqcwphKroYKLGtUag8cDNzau1
mLDZ49JKtwAZvw6TuNhN6T0fl8lja2kGAbXLyu7Nz93NIqbQfcb8Yh+wfZV8MqlqOE4VcJPTIlDe
WwILLWzlQmG5OucljoICIaziQHkD9FcdIaJ1TxpLrUakkBCgJnVDKgjlCF2ayPH7qjNJiFO3R8B5
/h4JqsQzxa8/U3WWfvyeDuHQkbMrqeXXSMwCw5tbKlDo6O1xjMzYXGJzzcS5J1mt+wwv5mjRc0Xo
b7+cn5jPCHrYH+V5UJPUf/CHJ1XfgxVlGmSHbDPNmNfK4ERMYh+xJCvwCSsTeY5iWxPYULT/QFtZ
F/r+3nMLbomfDm0pYPSwy3zTjxRF1vCsEMBarXq7F9SftpKhiru4dXdqHQwUkCZpf+EMPYTfeNww
8b565Ahvg5SwSnFtWRmVzrDu2gK97ldBUkoXVRyO7qpCktCL6OaSoSBvYUXLQJM+AsP/JUDTtDRM
UAmaYdjz8yX6hxt6ENTVZfDaRpjkzpcZAxsRQ6qH6vv6euPgbsSSB1guvxO5mhwflpwk4XYcKWur
6t8wPA6RhZ+qh9efuiQa4w3bx1j++KyQNYbBEgAkgNLCE3GJz92jhwIitPf+cScOy052QwLhp8kv
lB8OCox6G9sXQfBs2MRO/+NcIFgP9TmzXrYaz9m/AaYuf5dU0QynXGmLsX6KflfF0Rm2yLYLoL9T
y9FQeW1ScUkvVprvuM9L/bpPcWOkbVCvPDwJph6anv/UNfbEH+h+HRqayC+vBvTa69InwlK4Z2d2
4xAqI8X1txmGhblS0c7kax8P/Gt4HIgWuCCir+ttScBGQkVYEQVuuHDmCdF1LXhCNmyS9pt4x9P/
MZUc3ghrmJSDmHc5athGEMTvZr2POcUtRwDnFsXrBDUUgPA3lwUz/xw43BFXpiOq3yu0XHerTIJw
WMspS6lmkMLGcGdp4Yzw+SUaf6uaHwMD9U8gO5LCY5NFKvgJgUIxbA5zI0AmuZJEiYXLwzQu4RRu
NQUCouIrzAOParyN7eJrnfRu3wzSCEJYxeTE0J8oFpcLx6NrqWI/Bam7CBmssOvuZVCwmvylolrK
WXlZOtO6SLYjWAxSJJPD96SeT2ddVPKHzeqg9KpNcFgME3TmUoHpHRTiF2ynI8JOVNIRtA0s+J/J
mJM/0oomD0/EbH0OYn9hFr68xqqlWKuxlpnPka/cVHlZdC3jhVeYRjHrxpUtPABYY01OHBgsw9Ou
rHMrn9JveTl3Tb2VGXQXj1JRNvfGppP8MAm3RwZ2wy06rpGdrxggJCh5KivHuBKoTTrrI9k1TSzi
4IgEuBUgL6Deumgv7JmD8g/LbXytcvqH0oGWVuRHYO7GcQhgWgzigkxacBGceNnz2ee/ev4mEZDZ
H3DfSwZQQVCGzokJ4zXjK807iykjAymd5JndAxRsYEoJmUa1m7orLfUQACaoSV8YnCiswnBxe84O
uXi73Xk/N2nPk5xDw0MW88xLnN3Z0Jg1TpwuaTuAPYqgsr26ACUU0EWISYQtBmty+WjiNrX4ABMl
Nsq64qpF9VmHWmQc6ojiWyM5hYlEO2cYhWO3Xoa6k4A2Ksa9/TZG+UXA4BQbWUL0wjV8u1XWd3zy
iOBzyR/CVViSujQfguxY8/FKEslagVf0UMnUwWn0VzVCLw1xwLIOIN6WHaBYrwR/zvKH/6J7tpqn
T+dI1sM9aZH5W2sKaUp4+AkZMC86sTCGo0JuHgWuH469JWyALbcpXIEE7eNxsvhwnkL5xRG6WTfu
SY9Jk0fSkPSOhVJYMvMdFt+BwXZkLOc3XMT1R1QM++2l16Z/jS4iK6CXoDRgLPfEblWrhqCB9wIr
4KgM4I1fx1b5mMK74VjIaei7kE+MmhzrfF4N6Ili9IrQ+q9Rbw9f2a5VMROkOzB9sBv+ENjBuJ+R
jS5OXbScBDDE0RW3/xsCAX4MObd5kgrQAyBpo/Mw3Ne/WBo8A6FFUhMLdsCYYY2CESJj9V+zkuTs
kHw9l3b54La0Q7EI8E/F+4F85PLUp5ozzAAhk8xK3LjhULnY/f425HcVtNICRSIy+Ljc16UnoSQi
tW7clLE2JzxgiNA9mOyUGWUa7aXNaSaWDkeRzlb64IzC1UrvZlwv7ut6Tze+KaXvBDSWDNjZrPW9
9y+RLC7BWrDNtvgl1WZuPmSRF8OcidxpJOXNmmx24MGruZwgULJFWbCC/aQE9k1KkWl8EwuyiyxY
FBubH71VBIIr+fYfta+1rcysRu20AS0AGMIdMxzYGosljOFYnFwxSJyd1Nw3esO25vMJ+8NmTGvN
66pGM5827xKGZ7te3C2L+t7tuNqQE/1coJnEPMF+DuWc96DsEZFywoSYRXIN46I9aw/LeiopN8Bm
2KHXWGYk9RsmSFeIqXjqcv+e34U099+xs/074VlJzRvAHUiKE50+0Q5tpP7u2cqvLXqhW2orxrio
0l6+6KJj80UqRkTYPAnSou8XkPqoB75yD3sPYMiJY81oTzyUIxGU4nGEs6Ya//EhnrL/sN+oZNCB
gH83JMKlHH4083OCSAZVaKeR3qMKYbK94GlklIYXcQ05RAdTka7qArLao57llY76TqemkV/zwqu2
evNP3AxVKCjIrfQOzZqBceMrdnx3XNW+m/1DGleklZp4mPRc6HMlCvy9clJViRV/3VZ4xauOkeZg
ZDAThimsAeIXVUu5krkuewt4ws8ljbfXSnTb8ZYtFckEQSFY+ZQnK3X+w7XA4p3kChOAgGItfrJO
Z11ei9w45ginEWa9s84c4+GsTiktqcHju+l75rjGN+DXtK2Qu8NOqdGWPDPUtRRRmkcYn9m2Go5D
UjNlm9n2Bn7eb9yKa7f4U8noJizhKHQ+4xv2/kFc0dkn5wY7yctHLl35uyUT+T10uQZYHX+Oe+3/
8IWpO0+oHEzMP8Ij6STd797marrE25VbMaP/N3LyP6Khjp5WnAmexYQDDVulebns/Ue6kkuu7Bz8
2qLkq8dxL7ehMh2OzWOtn4TJc2POpyx73qoLTzsEHy/EHHw0LCfFGH876681QzcY2vE113EmqzuC
6mbbJz+U/GotI2k9yewx7kvsG3K3M+kbcHjNSWayeHIjopn0h1VmP/+CtXVfOYNgtqvLUEgOg0Vm
UPLGXNpiWVOuXNktQTXQDtDcZNvL1D3bJbkfV5WrUW5MFaOwX+uhvdAp87gjW4TAmgBM3jzVOG4n
JLgPiBlFyInlJGLLl+4m7+sxDhZOllHlf9PmK47OqGstR5g/DPK2oPXkPTLm2s2vuI53q/7wcTFq
uQFRg+donMhhKY/d1Hf9GO+i8zwuXlxh7yX0nnlqIt7M7KK33NlUwEC9J4aByoXDoxKjby/wAdK9
6qYQ5E+/aOXwUFsGnEfNoDHaIa/JI1XNGwDkjB+c+tW+W+RsqkRjrD9UpVfdhfVQpnbG++PZvH37
Mm018WZoC2rAuxIQrJ2TxCYesjCru3YyE3q+2rqb3jRfgAw3WGVRxBZWG4LKCDEdnQ+z6mjzfoBy
CV0T+Cmnv3axlhdw/Xp/EiYPreGcTLo1oW9HHI7xsQk9a9x8N3qTEHoEYieNeo/4hHSzAeaf0VDc
/yOhEpTVvrzfa8w38zhJlLOGoOknWHaGalQfKoufh4zPcAKk90msAodfLNwfwzNtAiRXtixaaHuh
DM3kh7Mzn1v8WejrTgTRKJkffVxR63DESqFM6rsaDg1QYTyLg+w29S8V8hCsjko1YG3tfbeRUGTp
db6NeV2HRofaRSVRSTNYTyW4aWWiYIVYPf76bdEi8BkdBRxBVibU/iCRPiRggwdsY9H48EHfgyjl
fnQIBBTzxwezGJmlyLhULauyh1ovJ73Q6tfvq7ilR2/r5CsoN20FLyLDQsuH2uJPm8zxYx1SCu9Q
PimFLdozh6VGZzjlKLMtOYsT4eTSXbR4z5Mr3LHCsR22M0UKsjtpkUHeG68yN5Cgxr5VBAxGyK/A
qrwn20A+xrw7Hn+rxSnb+GAN3HSwQUME8VZFL4gvFykfKBIcZgz2Dngxg29QX5RHyKHxA0VdzmfP
CrKl5MnFIy1MLeLmSxgGRcoB8qJtyH2S7bqN5fSmu9iDFN4KArU8zNcvRa0AinYJa4sDjxfzMNBo
D1TJ/FdOPE5ZB4mzSi8QXST56Xd6q+iYBNAB51eoTRsLxfYgnc4mI0/gzh67GRslqC9iliHkamaV
X2Q0fbSufGMtCfzcS/v72nKnPlqvgxsNO+HGm5xVCQ2Ro4nUfLEX1qQQgbApFtusn8rS6+ut2kj0
EeM7v3r70W3xyELYkhjVB4rS92oGwFzxwfpCY2t4RmMCID88hz/EL/K0jxQWwa1yzkzwU00AaQtq
OPFo8iFVmR5JDTwVnd40Yi46pxT52ktV9KsG/c90y95ElyTMESXsG3susgvv0RDjo9SCPYKO0GGM
LGvZboG15nlbnNr0Y1usfK3JL5kGDsWYV1s+NO7MnBdx8YnPngTPlDQUaVKAbBAlrOSKFR5sFugl
QvJVRDA8e3DCh9rQjp9cFbE4FOkk9BUylNeNZg8j8jIiDwrQENyNtCaSzdZot2x/tJxZKpXy2XBM
3ULQ/QF0sXZcS81jIlpnC3gwOy6rT5DpA/9VL4Sgk1HN/CZ2q/tEUTjzkoOdjjEOluCqGKYO/3Pg
4XzI9wQbw844G8JUG6+lamn1+cY4dysiphJ+HMudRmbp6ie9B/hduDougl6PfPVWRyyKptbL866G
WMiCzQP/nuOIDOFbNBlC6xhpR9OzSbmj3o52AJwbkNGfERwYTmX757DWPgcsIspO6skG7grXIChQ
Jk1bpdLj8Q4jWbIinGjYAcUcr2rOheefOhXYf9fYFay/j75e9FSUXqgX4y0G28icc3KBhoLvmAAQ
t2m/igvoPGhrKjdkzNbq+A2qjgnEHPpen1e5Ihs9/1txBh0Suv/G/AR3bnpWv1LbLUSmI6Wk0mIn
BUf6Hxb0t4nQpVvJDNt0rxkwlxFfLJitoFW4sZZdwg7Jk7cFaKZ25LAXDvjTX5zUMs/cv5IIpSmD
dNhEX984ARm5ZO8LKwAQL2VFCSR/3DVO+QVyIclOaFPVgZLuzfdIx4wCByxHD/27mmCD74A9S+81
vW/fKwwxlSKhf8fXMQHwwBlxKL9y7YGGzBGOQJYDhIErs/H/BYXkk4ONYlumB9O0VEptiLQYj8kE
orj9Lt6RnfZmric8oi6jaYtM9wgBIcW9R747s2HZo5/og2UNJp03VbxbdGfupD6xPAbFHnZeCUi7
ngYTpmTslyvuFRIMavjXJI1WjOP5eE4vjss+AW5Bk5L/F9rz/H/A5W2Zihc3F1We0xpfo4FhTuNa
HEX8mp8wAtVRYLYsDixI2g+DWwE1XlTR9R5EwNMKt39RTir2xNePfJcay4rSAH5ELQt86XXJtayv
vKZk2GaQgTSEUnX44HMA5U0KE2bEMrc3zFKW61f3WLTSX4xDvw99l/vxmgMu6VPT7vDN+gd7AsEI
FZAsWNdS2qylkzg/sOowIRUyQyFNjpdLK7ItnFzoTUkbeQEOkOpA6qJm33cWmUQJp2/SnTvLR9sX
sw0y2uAcfErlw1SDhkQ34P+vNnvv0TzbO6KPgX8tU/791kJa4SESVV3hhYr/qw7MRXPcxBYE5VIT
PPyXOsmB8GZJChbVfchr1z/sxNtWN1Z2UFgNRFNMkx3XyLWjzwlNbsjd7LPDLCLcEGIIRCPD2mG5
UAZRA5+zvEOBPAARFxF25k1lLEjdIMryvO6Dn+f490WrT6WRh0MGSBllcYjrOr1becz0+Lg9JR3k
uCxL6sDApcFFPtwZRyQeNP/swIP7nuex+8QbJH/pwgobxCd7bL3oJUrHGqKCUgLOGh3LF65rOX5Z
S8/3x8AahUj+ZAkrS9d+SC8Rza2u9honNJQv4sPzSRxEt3it9a2RjYtvcCK7cf40mECRH2vTv+NV
OXLWBGyjaZtr2hnAFWE1qsyKB1MMxxB9MIcgXhg63MArWUrJSKsuj7SiSV74kRKMVmabqoK16dn1
YLBNifV/MvWqai/oNnsDmCQTn1gmIpQk+6gKOmooutEOfhNY2YEQWoVfqoOyiYs990Jh6x+bSPZb
s/mQMuQXsl4KEXWJOEHl8b4TltbiJLlJxKrwwgD4bOvB4hld7y4829K2ldvWI2mHy9A0lNwrpn/s
Acko+qvmY5sewYRwpONg+nks5pgwDcU3reF+dTUcXC4N107JroW/4QIAvD/AJoYxDI6CA4MPsfDr
S54q5tEWufbgGkK4sHmY2ObtaOLxan5wWfhwX/HP8byBhJ6/rO9mGkrqIih4FKrXbk2dm6oIl9bQ
Hu8VV1Ln60txYGzGZyHzU+ymqq25fiEph7PqSx9GVMeHUcoXJX6Czunf5rHdpqpmThfYMGw0qOBR
7uuPJHGHnJ08TrUJMiNIgg6//EXHPYE0IYODStjoF3cfrXkg2AMSaqtBpP0vJLC1PPaQiTOZO46M
Jjv/TsFSBTF1MntIrXxfcph0g0ESc0MMeNI4Q6J1Aow19nLmU2705oXecBOADa9iYLCqgcbKb5ZS
v6H+A1mdItcYw6YnO+j3/Rfyr50bE9Nw6sS2OFYIqWfV0X9srCG9YYYFnkfOQMc7PnjLYv7H7iA7
qu1pfuZti7mXOYgLZQQDcK4/5upDocBxeiclpLW4B7uNDIqdWIpOkn6LEwHjfiMjDA9MCqSXWKgv
hXaKCFgMnI5nNWLyQvdOPnL3H8NLeyZEr/KZj65yZ4S+jjmBXtv9kQUdtnOccTf5NgHmpk9dXjFK
F6bXN6OFrECHG+L1Vpkpw7LE23Wba4pOcxDb3+dZybXd2qGT/bfv37MrzbJKQjC+f3AQPcbaCg6I
G3+oqMiFzyHsZ4OK9WlVk+HgEVzkzpTddXZmIHRUnZUcJT/h51f3Pw4Wyia3rk8CQ2p3ZBseQz8p
dC18jNyl3Rsg7i8COOHyjd3kVWOcQql7yuq5NK1JoR875RLzfkFZiLwNuvO+JVoX+WER2BOPG4bU
jhOI1pWxxLTyTlFAIbGWrNUxfKIR7KECsXqEaVzhLOpdI+cim9vUHx6pIl+4ynd/6aInb//bykWJ
y7jl7SSJd0vMM6ZNUqC6ZiZGHq53yDFBxV9M00SeG8IPs7Sl9l2wxp35fLWyfUzdeojO7b7vvGuf
RucWn0b6MsODugQqqesSZkBaGslmkZSr6IyxHR6+4OTD2/CgoVQQIJXwCT2tS5vwv42zcfXhrRrN
a0daTfxlKpV7Rosu+7a/Dz/6yvRl3eqmD3xLKx09Ry0U2e/1MMPY8YBIsgYWVBVYfFZImka0QNCX
lS8vpwj/iOTzuV3GnV63tvNnHGAoOni8+lg9Vx20tJXWb575O4IyReLzi7rCoLB8QDyBL2cLYpf2
EHXKPTm8eJ5C0Lzdc2577e9n84T84d/6uqXLKRqrOQzNyala9fvkFjoUKEIWY2umFUdcyDNFNgD2
YUsjDZvQ3AtKomoncjkKhy12n045HVMDVOMd4u4kuAehq3vyUevuvqfFD3oDs5NBtKyzajgPzyZm
cL27ZgqQqiVWudXe71JkhFtzFy8YQPp2lO7lqv9MOcwO46Yemoyh/xP/OSDCjG+LOc05cLgTMVN2
LboBjqvbtH47Bve+MEEuNO7eXkc6XpfnncM6VHeSlUI57/doQ9oJklhWsLxa372aiV2e9ECay4xM
/dHoaTN+tP2ZnJcuQmri6Y+EmBZt5oYzYBcC8Dxt97KWEt4E/QZQ4bEXq1WmcjL/bqmGcfbBBqFV
Z9VM7xysinNx/+Wb20x+1KrdZHxsr0a3RKxMlwUtod26hcReu80fpUF8LO9bYoPcJ5ovkGuKRjyr
TNcjI6+CISwog3t2T2l/BpDkhAcMHi3rxpLrRnv9o/KCbAasaQcTLdIvG2ZAxgUgT7s69twMAe6m
I6zVtrkfiFgayKCp5OJgzdYGSulR6oBKymfjEpExc5oFkpnFK80f+fpgK73dr+6p4XE+azPdjlU1
BpEIziPPG2B/TBws8BH+Sw+7/i+76aOtTjT2XYO+AvuaZR9md7La+gn9707syjGm2pJUjQ2f/ZT5
W6l7anqvveKMFdAFifTBtRuOZ10F773aDyy9qUvzq8JbDjMNh3afRTrpz8Ce0X+zxg9lDjHGXGAb
/+pyJ5Rvpo8//6MICUhQNnqzl7V51YKuq4p4gzo3oIyFvenh0mBHahqeh7L+pdJvAHAt+dahnTpb
5UXDIfPZKQdGpf/1ffKKRkRi2Z8Ue+HVqX/BMSAmmEsc68dbzZ/scdV6aOxS64KMfKX6mm7lBYC6
8MCkH0YrosbtXcxRPgQ4vHX6ZsWqicFKnMatmDiPtbJei82q7iaALPswBuEOgL+Krf2/JJyGxHYb
g8VqNoC9qmvHrifbUoYnxs172Hc4aqxh8J/AbMwhnMttsqB2o2nOfotz9wOi5huWBoJXL7LEPnsT
3DjYC+HVQol8nsFfXhAXVCokXlcFVNSBVEvzN80DAX39WZuVEYueM+gpvj1Wgn4EQDXSnwCuZy7x
YozxeDWSfPUXFZE5ntBxwYC867q1PyQWM9X7CK7lfJMHolHCwMq0NKy5/yNypfQkMAe1vcv6WGoz
CVo93bK/iqz1k8JR3WUck03Vz8OWkgabpMaB2v1MI2M8fF12OPeV/truvh3czSqcXrpkIlYLUF0b
6wupmGpwloFZofQ8oxYwKmWmTKktyrVhVaI7PukwNl8wSLNYlwcDwYhQCd7vUhMVDhZoj94QFi2Z
L9dGn2r6J29kMSF4DurjfGpg13mCFUYHC7hWkEpOzg7amcOQ043BSlYducNM5jkAk1oDU3hq8pDM
z2aDprYppDKBaq0fgTgYB1MeZDyREVx9QIeg8pJIGhqA9ZG53TXsKVOIvD5i/gZbgZfvpbr5RMN7
hch6kuZt3LAmJbIjI+2YK+ARAeO132GiCzlW0DyRZJXSJSAckSNSbE5Tqr65CIhs0CoNp8S/i4Gf
GRE5S/PJztnqs/g8G25ifbJ+OS4aPFejH7rWqQtvhOyqnav3/7OoCPWX7dvmxVsmF5OFtHPXxCqq
XUl+GpUwnH7pbF/N0OLbmwrxm+nlwVSgB2EV2DfnLN77GEv2AkVHaoHgSe6SmOXcRvFPlk9qb4Qk
qAFmKLlTQ2kHtc0JdcMeqvK9tS9uijSGG/CTF7O8QMU9VAPR7fQmzExqSu8M+NklzNSbU5gV+1nV
zXMFI76fN7ZpmcfkKnOrSO5TR+71BPAwxtbeGnNxo0Szq4nurNZ3LgkoUxv+aCaRdJjHzUwRiTCv
FgytL2s7TKghxeUedTAPxJgPaA/JDHxjz5Z4MLmQPUyTti4H769kAojC+GMuTxy14eXNIwunNW7/
AWyIM98sY0WTBvLRB86PRK9izUI6FyFUWW1We2roqTV2Fu9FwP3yH7W7d1M0PNXSU7q5ARwREoSm
ljKeayFg8hXrXFJr5ZXaFqMgfB1WqFtBQVfQrJBs7PpPn9Ps5eUidiEgZZqIsnFz0aBeeuSLoJ8h
R9tvwwoObGgI+rtH5dSXgByprpUoifDX9TPV73N1g2ilzFjnkjoMdLaawDyy4PV5chDmKDaXFhur
SplRcBrJhsDQR0Mg7dGkUOUyopE2d5xqqSjEMkD+ojNJGHysmnhAlR3k5XaFVxxbID5EvKTX98QG
iSmCdCCkB588XWjJ8A75mKPnj4VVa4pj1F2ObR1qsItYpcwsGYajv8EqiEcpti4RwUX/K8vPx3LP
xu5ON5U6mIkHSJpK7cDaYgYnDN854njmZNr37r+BRG3duz+W0xFBaNh1mLjwWH8mXT/O7qLEnaY0
qUsYLwjQYMFVoSApp1/pujIzlPL1k0BG6VQvC4WbZuy9MHrikUHYw01FbWTARKviyPF6uQNqaLa9
JFCA2GJQw+fRGE1IQDf1sC0rdJ44/53XuzIwklQ0g6sOK6r2A4WZ7laqwysHxkL7YoxXhadpf6JT
L6S9HiYLwHJx8sDJLipp6H8qXpuHXfUGf9xwrS7CsHq8idqBHzPXSBirMt72pxXj2GixWFRlaPTB
dCUZ2F8ds3+DPl8U/kZD/Jv6b3nTxMio8QhXn7fLmlFwN5L0ifZwgjsDgnriLpx2ZmYCaI3jOV/w
U/Yi/5isf6tewCEOItlQHd2dlvCDGb1TxkOvZbNi/zRa2yCRbChfLlHdDWhpXC45XfxIXitEfxUB
/9/GhxNx7XyK2BV+nTkP0PyC0o1Q3RBoY2YpaCPxZ3hWQ74CK2n+X7wWAWjGslzPllghHlIl3KtN
i0z4WvmYLBoymaNNn8c53p3W/AaUrLT/ntG1jY93EnVFkggX/ZUZpV3wEVDp/ZsYEzjJZo11Szey
dRNYp14h93GkSBQx8KF2ficvqpixllRZ2yG7jOcp5Br/wEfm3kmab/fQcASC/iLAossSAmrBwRqu
r1/4Xud/oelxcGEvK7nLP0H60L5DvZd128BTFbTWSv/jxTn0bGZCwNfuGgHKrf6cK19twF0KCLkf
Y3XYqsdwJqRPPWq0PKioQ6oLDCE7lDn/8RkQwujDyJdusUWps8RDhAL7rOlmWIqd81nSG41bA/CD
JFLYyPhy3mtsYXvG2TO8f+xmylcfFzv1ZNA0lyl3FiDDLKzMXVNuHQWpoCMMkCm+AUaKELcxYssX
iqhJ9cEqludlvtbPREjSfoLXuPPqQZzhvGN7iNPHeYEfWrmLyMtAQwTBUa6ole/ieO1nFfoTMVqh
dlT4//+L6znB5eqfb5xHXP+KofeMd/IeAElbbVx23gNeVCbX6M9zVslB8WtdvP4cua6Srad/1Guf
irEoaWj/DDd1jFB6qFZ/YtKAqESn5F9l0czJQeuPVPE8QJvGfEJSkXi7YBFFZ6iElLL35EkR+z0i
/jQgmiXByMPckPOjnFk298atOqVXqx2YeHC2abQfcM0HXnodUvFG7ptw26wJ6tNOOfzPqfMRvUgR
ZYTuYuRulLklBOETpVOLWbBhyIxI26hibuaxPRfFh9aJMmigDFFeLUa4VD9emnGZjHkHwfyTweEH
JeZWODPUiezl9g77jcJ1ax7lgS1wliOBI6CRQ9YxQljbxXosdf5WswIifdqcoFhFvNV5SsDkN51K
mU4UBkIJoI+W6Ci3ESpKMeAZdNzsycFdVc/7ixyJUjT9hb52y/gcQtzeqfUxWdUUy0tu1Wb0taJa
g+BeJq4zWZ48EY0LgpP/fT3SOg6MZhyNHBaDD7GakkQqg6aJ20UigNkhN2ER5Tc1ackExrIvRJ/5
j52Lrse1vrJ1+12wzUrTRvxfZgp7V6gwQkVeGJBdPjMhvRxo6xINYwuF+grBLA47fK5LqyANa8In
l0iVRbw27w5ayOf70xwz1BHs4ZZBgPkPiqwVfWiSOrAOGf3h1XpZfmdtfevZLSBGF3RU1Icn+vvP
7189to8fXRS7x7vuyr3mCc0CqxYgw7Ic0t866CeH6QGTJbevwHPIwBCyUdV7WUOikIBsLjNClWig
otw6Tkwg53mv+JQFd7CuIRC92fZW+ExH6eRXSHY2pH55pcQ1AVvEXz3rkKoK84Sz0A29uZACIUH4
24Qo5bESl3zxapeIIK4TEisZtu/CEy8Lk/QSrNjPcvuIqMo+L6ggDA7a7wQQKZbX9+kUfKw+qHi/
OW6+qT63q5NXwYbtgGel3hq8ExyfDHP/y/db6WwpJ9CkNxv/AtQH61uweaM3Z9tqLecjg/qRHRd/
tiQybKLkVzOJjoIvAM9/d5K2R+yT1VYDj5zdz1HSM28q2lmUP2cCwigt4Y7AEls50+y3Cw+LNWt8
mvdmhjEGqG4zx4fq7yS8tkbM4kfTecgElljkzt3LvEnX4/9WnX6omHQZHiLFjQhkyK0a4nNFS5k1
TFf94G5gEiIkzFnSrVKZZIHI5wgLJCBqx3aTxXiNMc5W0ycAOpJ7MwpR/I5O8u1wB3xtIeqEexkQ
3hxQgGAOyfxel0TDZMs/seS6J4PjIv8J1Axg+foNkFguRVyiR8+ATzzcH4N739IfH/ySHs2Zbs2G
fqwq/d4y5YVkon+pBJajm3syH+Aw4SBwe8i6zKdYuofkOBl+HmUREsubQQDw0YezVpQaB0YBLQ30
acf1xGXA+NriwDfGgDpYBzfX37V2B1pDey0Xem0Sr8Poia1v+m5bn5SdHqYPX+Iwp7rkG8hBFRwR
P8+un11uvOPeO9kjFNUTeLbiXku6+r1lCN280/xKYlXUZuwMztVwJM8sEVK0UF35xk5cNmTgUT/E
s9hMg19TeITccw8feYFLbKyPTZYaw3udYG5n4XOGz3eOBkVi9ssmRp/eEUTrxUy8o7hksRojLupP
+HFWgl/mfQ58FCsS9vAWKPKzYXRkH9hr5oohsZ73wR4yJ2yaVOXtdSM25L9fjaOqEHRItVEbjhDM
nlVap74j1XsVR2mnOmbtpwWc4xNLFbru3Un7QSYyPZnCu3ktQEld3JedhTT3bODdGhgkw11aahh3
6jX3eqGbvx8odK56f/1CZNtTGEIWhc0t0FEWwSUBpfUFiLkwM5NZXKndPkN1z/G8L/HHN1V46p+T
vARbLWaY1qDHZ3DaW0+KJ3w0ZlOpAGdTht3xwz3iLYgMjx0RZjL5XYwGrCqmur+JwmLVNRTBVdEh
a1fejHfQG63WTH4tDoOlBMypFITqsOIMAy5aNFt3DNtyVCKDb3GIZPuOtC1He+//q+HnpNdGlvo+
4YM2si/EGvyfOX52qEG4U0bIDl5ytlWKdtWTSUb8gMe/wGPoRzZnbFZSjrMS4Ospw17kHRJVM2hu
t1km5+THoHqDPUp0ULzrMMBF6Ewej9fOy176ryPg0XhxnMdXrCq4kIPYJvIoq/TAjI/Hji6STMkP
848tDwO4O/zl2HRQEKCvWhSwKLu3wOwvHI7UawlXKcAbCyopvZjs9kHGRK1tsEct1k7qheXv+LXd
Ibb6DeGIDi/tBi5BFAsJO+VQxRMGrbr60rA55x/5wK5hzu3HlCxhp78srZmvuWSdR1GScKEEn6nl
zEHhM4u9iITB3BZTTp2CpRB22sLP5HIJDMc/4mvZzcfPNpAuYMPywtGo5xDddrn3TezBKDbBd8IQ
FymClTDBS3WLOidZfTddp/qi63WOOPkmgUH4qGYfRdpAS4Zz6PwF0g3s5zgmJ1G4VuNDagZXcAJ/
/mb9iOGo1VR0/7qcLTFhZOUluOKt8A6SGRkY/uUbLooJMYSM5j1BTmTMQIvL6FB8ii7P9I95u+OF
y2aOQX6NXgDr8SS3QYi+8x6sVf/jXZYNiEgPbETpfaNAg/HxD45Rak/2QlOCSeP0bQdbEEAWhcJ+
rjLEBWVZ7o2ioBQvM93nydjC10DX2P5YGz9LPGUbay0n63+68fgerhhwVUV+DVBVtzF62rqzyHHl
+TwQwGdD56Ap3mYQq1RkWvQNgggBmY+Br3d71M65s5Y0KLwrKZ6iFPpeXL78cKHNFl74LtKLnW73
mrqtVaXqH8JbHdEgsxGMfRZPshrMP9FDiief2LPs4z9ltZRIvSolGbwpekFdIY64F6zR/TWNhBvN
V9i5JuIAU6q9wVnfEd0pleRY7CnGphTP6jC225Aen7kSwVeSOMgJPg4Kge5uGa4oTGfQQY7Ru6pf
AWFI+R+OrhQYusjKfrkz01hoMpUqlkonVP36q6LuUJITH5PKvXuUN99pZwyVIekZWOs+5is8aZ2p
Rrc+myJ5PFyH9AePGy/bYSP0VlWaj14syooKyjgjZsPtRg9vrtL5b9O6ZTvv2VXLOW2WK3OszPNE
BZr0gwPNWmJ5Epn8GWPplR4/BY/ggAxcNC/Dh23L9n6FKQvltSuRjem8feT75lNPJwd8VyyM+ULh
dQBQptVTRtEvWgrkgra72S2aCNM3RkRIjLtLY7x54BeNp2qOCLRyLvXZnx9dILdI9FCddIrIzB+Z
lWj2VtqJj+vdVzLgNbRbsTGdjlBv0826GVE1PF5Rf/FAGNgd+rA3cp+qMo2Nhrpdn+uBzzkPpf9p
HBnNR81XKzgp3QZ24A8eymr08e5Ni2NFmKIR1odWD00xW4ZMgrYqLtDkSRozWXzniEO1xSxG1b9H
zB4AtTF9SPUcdMLxgLFQAHq6MAandoGVSwGjpvzu+i17La8ZXeuZSu1t8ZtQ4RTTBlFpm2a0aRy7
ryCJXdLXG4cdTgy9DkFE9oZvbHoYFR/93h2KqFYaJV27ZHGb0ZwZs0kKMRHRhIcXQgwQfGV7GaFa
XuRAyDFonEA2iSAuvLIMykg627KcjlXibJZ05KEu+MZBxbrOxMpsq74w+oF51uSeic2b7Sfwr8BU
Wc3Z5jJciEOHc/krVjQem/OJuA2erANMgDI9eW55oCfu0RoQCiPnl0t+N3Xv1hWL835x+NvIOvoI
nhMc3GwBp56A+Q2jDrgLavw7vNwCj0lesAFMOLxMRh9+oLvJ2k/90iSdzdWGBrFIZjs4iZrY8l2o
t6seS1jbsIkCipk9TiPBM+xFKxeEEv2GweCIR/r3rqvEFU60eKAnLtBWd0NZMrKhVRmti/veklIv
EFLqH3T9ERno0R2SDnLZTRoVEB38jQ6s09kBBcgWBgyDIRCKgglzeTz89IY74LlEXfc3mytw4pRT
funm33FVvz7NFm9GRN0RMXV+vuBNg0R3Kh+d65X6GrOTwf1jEoBgMJZcfIt0VLplFk4yVBzQVNMX
p5zZz/rNWAQgD5FaXlJaWL/p5hBRwdtx/BKyrMPiWD40hF9tdeKzyLLr+ZkMUuU+mud9BLxjqSno
qpvBnvDzyG229qA2n3Oz2NBuHTQOcewVRRFRrkcXfY17I+s/soC8fX/MSUo7bkd/ySzEBPioh94X
lKa4fy1Pwl11gzpvezm0FAiSiT2fME7O+RK0GJ7r2SykL474o3tCIdmy5myW3+jPk6E/BDp6DGx/
B3mkv0z9YOWlGRrUQn4RXPdSy1m1UtQtPeb89j1LdU2+Xmt4hxVJX6HtBqIq0eGq92N/jb1RPn+T
cjrF2za+scun2wSVAzQu7Zfpkh6WwKSSjv7CAFQCoidWPURTH1j9lA8CBKUlNYUUymKz9PA+NIYZ
ME47arIMqX31w6fB8Yon3WS49kxwvbab3tZM9QZAR/60Pb+2i1iy81GRpXwSWIhGGKwhX8oJJc88
dRwjC7HRsn7Yg/AuWYCKrF2IH6+NGJmweeJHu/pa9j19FEVxZMFp1gdwpDq28DxIYI/8wz+KeUWQ
oc/EmifteIMBX4b2h6JensJyOCJ9LLQOjKJf6sIw6v8RScciGmv7nWXI4qnY22hHiHXQyiYkbaLw
sCma4PSJ+8IQJadp0clXx2hIo6X43JSVItRD5kZbRJjwY249G4tCPsWlsknQAy28CWCXY0fEmHvA
xWV4kHe809BLw4Is7CSYZqtLeQqmSdjHMLPmaopeEyxCKzGDeOEW1+wkpWjGqpQuoX5c8Fc7rzqe
ropdTpoKEcsJwSBYLpKNCnMjDvbji8MbaXcNWhdaKyjx1TjKCsQmDRMP1vVcUpUTRUi3ajgR2ujb
pd0knlrLabzWs9rKcJsJk2K/oYwjPSQNUuJzOA1x83aOdsujN494fCrdYA36gyjEi8S4L4CfTCOS
HCIrBHb+7KhU5JmjN9XVMfyia3Xc0eZeQH7VoQPyFHySNU9jnxfYdqWs1SMuaPtm3pC27CwTJOZD
F/0uxcI6xvTsiZADWYVoL3JUEt/Q5ddW46ksKFJhkViQmcUlc0hERjYns76EO77O2UBPojDH2+72
6T5mTpVOi2dMB8TbgofelWL+2lbjBL97xfv5+Bjtttb0FOU4Q1xCxyga0gn5kB7bxiZrjlpU8vIG
5FN5eZ+EOzQt4W+2dpQRF5cNg/cY1w2eOsKSGDd8LrMffdUkiKkcvacjdixg0Lh23R5kRW0kIGco
Fk7W2ptpBM2YbJYu1vFrRSPLKs27izMoVp3hW7UnAzchVBBlot0ML/Sg4NzAB1U48w0CftOfE0bi
03V89iX2wqQsS67EpC8McIwMxh/mThIk0CSzC9bOpZES+wQdWo6lgNpLb9oXHmOnfo+fbtajkNXp
bwoZmdQGUR+4gtycGt9ez+rPH615KOdfGBE6pfYLQTy3mBAPUeUx/NaCZw3rSx2yrMVFPMqRfxft
T9H353DkqsZoTBlwB6BbXcLcUBHUmIWka5pTesZQnZZVOUnN4Z0wbyvzCzI0rEZHKvdIE4qAoNaZ
wpRJI5U7irCwKAwn/aPVdF5Av+OdRbN+uIIcGkmQbyLU0l6B9aS89KDwybsxA/fF2bm3DK6flOWr
XxLr6eKzhLfzAU9yBNVlGrLpuEAn05kXSWGsAQQX3LAhWcNn0ttcFumC2/7LsG8rqGGvVfrrGTUN
hIsCWqYze6kLin53oCpvQmAhXjzcvN3HbJsxCzy7JUXPxqtftfK/KBuIbxxEmRQLkwt6HtnxKEcX
qRxOsUU/JiAhmumLWG2Z1/BkA32WDcVyqL+EPJHM1L1ao13r7uxtP0wdihsdmiURSF7hlsGYjJ6M
TunbeFUHUmvaM1owViMNg8Um0/fCi2fB2U1fC7LooO2Xfy/np8idl1gVo5+4bI4i09OUG82BMu7D
/NZVbLlfWcrnHpf4U0VCcj06Nccq3WA+nJr1i0GopBpE7cC2OWRSUIwWeApkRamDgufI/uEXVZVY
xjObGf4/t5lnjsg1xU7Gx6LGuI3Kth97SG44jMbrsHziSFva4dbbnQbhL9MNUUWkFG18fm1HRIVj
xQHII15bttgTeoFEmrZ1GCLIeyLg9aRCPbNGEL2bzZ74mJV/sVSQfv1uCdAJlkiBM9Ul0kjqkoWu
CxLPQ8Lwg8DteDP95iN/Xa+BaUG6ENa/rfIfrvQadaypoU/OFMENyorlYhYb2tyx4qd1boa31JOS
Xu2ARcy71ofXbYmKeW+mMkrph3bxCa8Z7lZxrDBQ227SBi/ey7PkYV49nQot6rSMFE3HwgrZo8Hk
O4RebBvS9R4YncbCENG8bO3TfVJOLRSMFZL39rLimJ1wPp8nH728+MZenfvSvUcvc68RWNjjaXx2
+SslIC9ejDzcP3ZG9gdYblUZjljhbEq1neDHxfCqiTMiuSJZRjV0OW/6De+oMNBE3MYJAv0FgOF5
qyzSZD3lAZCizj7iIt/WbtsLN74KlAk8gDpV6iGugw+9WDxVaLvgNNrFTKIOu+tB9A4s1aa77j+i
sLb1b02OWVS2LCYLuPdJHbM77odj6H9XjK5X/U7xJaDQacEkX9PIL0ynTVjRsxQNpINSCSvGKfQ0
WPTyfgDg9gOUBcSTS9jJnVzBOmjE+1wjuO/JxP5vnM2NdFXuZq8UgABdWnCcxdnBwBIClOId1qrn
yCdvywLCuU2A4HM+a3ealR7k3yzUe9SqS1P1rgfXcHdngfcBsUoRq3W2n1K8RgzoXcqbmuWR1Spt
rzZtzKQ7QS89Cn/GMBy3MxaOYOpAftLNmn1UYji0PJC+5ElQofYjH3YtCzipsCeMS9to3esxWxSw
CaQfy9FFjt/rianfCyCeh1ZVGixPOUrafZmXgnyRJFZJIfGduzDA4428RGQIFP2VQNMmBR7segpD
FTsqvHDMmawlALYuAQIWmDtt36oTEVsX1JU2JEwVOHpcQVHa//Oedqy29R4srgtQoi49BakcR/LL
rMc5dIAQCqvMpKFhpOpPUlNY4XahlYcf+rGSNWgY4KF4iq5BFX6ySZfeBRDM+LB4izGAZ4yGXOW9
+40LPCBVQGWhlaEEk4Tdi9WRzxX+62qj+IJAQJyYiB9hmqw1zf6jOgdSaZbxQb/H+s/FGdmUW9Vk
O3kRFiny4ylm2H9A39ujuZxEBwCRkH6HqPP8JcvFBoGD/z3XvqH9RkHKZtCNqdFOWcXGd1KBoSBt
nGufaCV5l5dDyocWs6ltj2btBPifK6txIoOdbA5zBNcSDuEh/1N5WPQb/uOZQHLbSZoeupjZPYdD
9Ked83SY0uHQnc1oKPK/1QAse344mPUVEOIIiUkAsT8oeVIljiFIsNaDmE6DkxW5biecBE4ZwanH
vLZTCunjkDbanLaEEtRYZ8oWBEFOxmTutDLzA5ZJSC0rQLU+0qNaSwhBsbG1JUDNgFT780YuxUiR
i6NBQEesX58Idw1ZIuneGmRJtmmG+HfhH02YTmA7zfTf8QBBTFTLuwSroD6P0qI/10AYQtKr7MjA
PvZhqlUXAeNrT0zYJAUbUV2U59oPVaui6/2mi49hX0jY76Z5bx5VQKmsIW9eZ/8WMXQEo78bs44q
pgc4amGB1ouXcdet+wdWCUUnfLNCAIik610bWWV3qLv3Ib1kigbjJNQp4U1Ok3+zC1NJIAiI7gMg
NkPr4kTE7eIDDQskxzaUWkPGgGhptsP/fernW+3wlbA5yywTs9qxDJbTqv24dS1yBUCSqxK+bNOZ
JW4CprXLZ4EbeH03MjoB2owhjsq43EGzxhiUL1sDXBuOOh03vpLbiIFHPb5vnZnAON1ownKE9+el
n1S1RsIeNZFnYcNFuhynptO/Wm/thi5hVKcwb0wJypvS2BL0YVizQGjQopqbhCZ8QUbPnTWmhLdn
CVmlFgtE2+UKuevUBYMhyOAmDlZsRUaH1Yta4++OLy4PeY1ukvr1JeICZDPpYJLUlUr6wMsUm99M
D9L7XvdB8FygusTdEO4bOG8Hpq1uf1zzxnsJh5Ce9q9eoVj0b7QiMrawY9t9hGlkYAmPy/Prdzqz
cBY/fEhraWulmAtNfIzgn5l5iVXfxj89bVhc+G8/mDd6UGi5Is0jLMLt+7zfNYdmWxol6O4mSSaR
9XHD/PGf7QQz0h3uvKdcnT9BVB+ECQQ3/AI2u61xz0FmHzw7lFRmFJtX3t5A4SfLTnOqAO0p5pFz
a9l+dLQbL5ZVoj+zFGJdNH7cXNPMet87RMxa4iF0vyJx9H+BQAGOzI1RHt99hTf7Zo6XgsurVTRn
298F4BRM84xemsIKOZhZsbiXJV3oCilwCSRjAWh9/kmLAX06MBVIrrJA9tgawxSPu+/jF/2iSMHD
iVNHyp8j9ufEIvwT3DdxcPHxwJpWh3pQQJPSImPOMhtMjM5XZHCKG8PczUCjJAEDjwlLb7XpnIhI
FAVPhjWXRbPKXVwg1lgJ0OupUQwSGeo25NbyST9jocySz4fAfyjfgE7Nv/0e333rpxM/JhKpCeaT
kvzCy+dzDUd1pavXjodEKbfIiM7Z1768jk3Md2IwSHuVokKEREnBIN12QGGYLmucvuAOT3HBcBBv
oLNYDV1/wmQMJab6RMUOBJRBXrJ/WYInQrfSOYbCPwq7c+1oddwuQbPfaLOOdXNO7IRYuSJud+Xh
msySjNfKspzxk7vQVDBIyrct4p6XmcjvyN4S0F3Usb5H4XVB5PckAX71OBUHbXEtmaVJKt/DoKoV
wfETEQgPM9SsY1HPB3h15PbPaPKe3Hxb4Ehia/ZOikg4K335gRB1+gae8Pi78v/dUTe6BYYTD2ba
25XsQWoQ7zNkm8OadR61ZajFzJrTI6y8qFexcJ70MI37MglPGCebKJSvK0L8k7Y9osxktx/82AZ7
B1teeFsjvo+UMIbM/tNIJUX/ZDXMIK2+y9t1EZ34e8MMTeFDR7C8khdcMAC1y2j6lgQ6KYwGyqw7
XwVswGl7AnPSZEnN+hdr6SJQZ3oXUO8Tc8DsOf9lRj9JiOJd/QMapN7zBmS3CToLAq3kKpWtYfqL
AYsUgBKOhuzegVAA7FQjr/7gG1qwyMDo5i0VRRkl3rx9PsY9dh2Y+o2QntQ+iLvgqlCwonLkVbDj
mdvLtM7TRwZRt79dKCXO8zDMSLnQWlJhhYc5N7NdgTLmaiGsbknKXkk61wOiEhuYS9NXVkNAZ7eC
OdSaYNqSFxDr6oYWDQpT9wDRlwVPTQ8TBU38umI+/zEeyx2m17+/cphvvYa9qFk9hY303a1pQ4ii
55IoEawjGyyJhu21yWdmvV2tfdF4AnPC06PgWdpBMJOegVXiq0yG75BCTEFgGTUCrh99l5pUhD1l
NO7oSSPMKsPxoaEAu7HedOVkTK5kvmLqo2ZKLABkoEScN5li+iCSM7Zdv5rgU3ZUWwI6NchepiJL
snlAvOnSa1E3hq1nslS0pxbysaJE0nuX/Rm22SlkGWga9XJF37eEGJkB7a2IiSa295GsGcdPbnCZ
4dp7Za28gQCvzZ5DYLkmIu2RrrwCbpNdx0xKw9HAfxaZffCfh4BykjBGS0DjCtKStHt4UUbubtje
qAUZVg03phxa4qBB/G8xH4d0STQ4KXGuxyeVOdAKdZEo7jqsWzCshhUxdiAVuLnJcPtxJwpp+HJg
EcxW45nUUwY7fRW5uOfcyMWmp65DFHJbvnC3adyeCYE+4uRYqARgXNx0y07glF3Dx/I0SAocY826
Ol/P0NQ/foxNKpeqH4OoO1nl72q3BLcPdJszUCRi/wRmBNtq7Fchv3euNCCCRwzi9HodNmx4hyxk
u8yfxXfw8FaYdqwuOiIn1vvGLpb7jngC+8EwjMNXxUzmV2HuWjg/po8GieuFh9hN7CbOdJe+mrEp
Sk/iuAO8qlgtLMZbHuZ0d8XR5qtNL91RzVsYwW/NXxMCX94ppGIHxfaZ9+84FGCaa9cV1OvDJfWr
NCkQa0Io6tI8Y3FEGy+smxu/oB7AAYj/N/K9zcaDTd/CvNvwPPBo4dtwxsIRuniAa/wcCw0x+lut
QlgmHOs5466WiLIT+zR6SnK3NQ5a0l2hZaTPfAfJATkfYuBNuNX1UrIWjkPQh9FnLsRqMyNMwqMQ
DIZTG5EWVwLZ+2GyRvp9nPalOlgui6ilwQANnDp6RCD5N+Q5O5Yh+cvmJXxWyy8x+XSGpfD/Yr9/
zV8rnu4aONgB3VOkEfPhquMDv62C19VF0Jfjn1GYReK1eDvtHL1MpAp534EUlOOwLPsM0zZNQqsv
a6fYwWs7uG3OVwzpNpMf3XlAX6zHg3EIPnHs9TXBhqEn5uqrqbjHQcB7zgRyAIHkQltPSkzCVksJ
G6ddK//HAIH82BXcHxVsr6RnLpJv1kr2O/NaHE2e0HcNBbOB4TJgfbDiljx6stCfCHaQryfpi+NC
rJMBifK6oQTa7p0vQQFP/dG6RZm1/uDybZbuTi8K+0P29NjfPCi3bE9x5i/85uATHmRkOef+B1Gz
BkK+CaBJzdK6taZdv4sItwp++cyjEPmCeotS6PzsLFLUc1xEgs7WDwtUdjG+ZNNT/3JTiiIx8Mzr
0odixmgGQnmR08tC5479+MIG9FqWmYFwPKRzLiLlvU27iNikYVAg6JhKI0XVFjhNJVzoCRrsGq2v
p7zZhtTzfUIgJEx07G5pwh5BqKUyjK4Nz+PlfAiKJapEKWK4kSIYy7Mex+6pBI+JTFVbSYvqgAfR
9+JB4ekoRX1lK1ZCgQHmZJGZw33IDh6Qd3lGk+AD6wv/R35Ei1XCe+GetPTBBoNK00VoK90YzihI
XGVHn1bwoNtY8sz8FqvY03TQlaJt0boUOPxUs/qOuSn/dEuBaWhUlJPwuwZAKuoIzruRZRjNm31Z
90cjs9oNycoYjR4a9k1+wfO9QbanZiEqB3fITdn5zxlRe/AoU0pddR0mxj2UeWku6Q4+olkukR95
mpTMkhXDvDS1SYmC53G62jq9hsR2VsTr5M0evgH0ppGc8phfkpUOBCXMPjV+6PvILZA38RNMI10e
MF7rEmlzpdMg8iPcGm7MPj3cdwdeYkax2hq680dDKXyhdbYOaJ2F3Zdek4jq6yBhky6U3648E0lu
1KEWkI1cKpAX068F+p3nspSklErDZclTGfdwjH4qp6qVs12dM6QQ+xzvotc2dcv3fuGm9Id9HWzl
gI+HXp2a+/Z06xpexXux52TOtyCVLYm3t6DRuCyh4cmd8juc7RxZdPU3q3Usb70jtAlyykwEBKD8
fhZtrLNTDt90kxpI0TjfnwiZyOxkvUDSpECcK86IpfJMEHXJmDT7yw7BRcziFfB+fakBBG0RLHTc
3gJ/RVa8aIQiSuH+ApDNQQ69YN3/8xQRt4US5RhZFkY16NHm0tvh/RQXiL0047kJa2d7LlI+tRDP
ODgzPjOq5WHM3U+qM3mTjggy/nLtBHsJuJ8xk9V71BJlMmYcUukq0izmhQrmo8WpZftUsYjGrNpF
PwNyR5R8j/HjdbQ63Ul03CbLL0Z3+igwzMbm1LXUxkPeaBcatHCAut9XPIm2dz54r5cmH+CnqHXe
8jTUjGK90fgXwtye3zgr0wM91XlYGQz7DgfpMyDoo3dZimsX/DdAlLLQhWqq/L0JYjMztcxea7r/
Aq0H4rNlwfQJ2jOMhkRstXjAzSLNXx5eTCEpqlnV9I04J47+5jzt2ekX//XRYS2QC0TIVMC4IWDc
LaJd27p5dzUB4lKxE+pK8ZP+6dsFaY5om/Kk4s138FiOk/sbmPo7V3Z+QzWXMbiA1nA6FqqT6AJy
vvGNt0xJq+dLu4pO+AbjefRfuL1FQ0LlDTdGet5cw0x/fcX/aZVZ6ebQJyePxWZvYa0nf54FSStP
t949oEg0VeH9BcdF2cGk6mVke9xVRR19DFucSogiu2MU/+cpcdJ145gFZ9+j2Rej6na5raiiMmKD
zQmRh01SHuczbsrE2Ozh2QKgrYZmqg3bHYETzOKRygBGj1oNIJyr1tgnmc+cNqhv/ygaXi0rpmx+
Sq7kHvj7QRW4hQf/M170RI9A+YReSWu+1QVkc2oUoQ+yocmLPepboAYoq2BdRWhntFt1vhsDuap4
9V8AtAiTkJaKJxNO9Gj4X3+4BwUXtsJ17ew3G1nknjJs/jKxXkVnnm095z6tZA/Q+6lwdvs+acqu
1vRoYsAOf0HsKCutRSEcX5hhAvZTV2fsvEKuuzavLPtnLiI+GdExLABIAAXPwTQaLYrFTVxJTnfo
QwATIzYLawXxfNYwea0MzdsSjVc+a2goVOGckFUln20W6560aVoLuCyJoCDwad32XrVigOLZAal8
TOoMQaEU/g7QDaiQ2fZrT4CRlycB+/su+VrJapLtpTImG5X98M4H5kjdrWpLejAnJ7d7ZUyfTt2I
HDryWSIoAW9tZ+fgrHzjEtGHLTrj987aLgQIF0io2VCxGWYimi/H0nvJCLXYIB/iI6Fv5Z94uR7S
MGM46nG4saRS+SvlOmDXV+87sjM4FTmOkNOpMAIsThv+I2ZEOGs3fQDc/Rb1JEX+kT5mxI9OJLh9
lTJRyW4HUyeU3SHDOcVFp7cYvSe77El7oiKcsovmrdVNGv79ivZqyRbyDL9TxZ8hZyC3JpJTS1dk
w7+f2NBJ4K0GK2B4Mt+pWLho8E0fOYFkPHirijb2TXVXKq9cHqk1U1bth4dgbK8R2e11PFTYjWuG
k/ygESr650tl0NKgtTUZx64kfQcbHEzN3mI7Cfa+g2RHhyzEtAfz237RVIU6ZALZoDDAbt6zsqFM
ZBFXAgZUDPfKLllHF5OwOkSTdcF31Qm41DRBetXGMNc0eLdls8VI5/Ldrz2C+3SUDDvCPX0AHmKc
8iDb3f6nxRC/n6us1xiHpstCcK6+hy9TzWPb9vQjnoNXP/p6soKZDRiCn6XoxcPv43sf46f+B7uI
Fv/k/o0+lfI7QE24qOsmmqrQWR43eqV+cwDGPOatAtaEdW7tLmRaS4VyWZjbyUfEj+Y6ZRnymcji
h1tTmJO/9gxM3xVVcrfjDJ8HqWBcW27KQUwXx/ILoZg22SuiQ2fW5140kWO1bAsbKV1+MYtN1yc+
qMipHIkPza9CRUVAfuavZj6ydmF+cKDD1VNwt3jP6wDluqr2uCy/IuSxdiMmOMEdvcem3gBcJFFK
gpE4jAbbYbgdNUXhwYyjJTTiGUJ2OFzxOXpc5AT/cltbs2jAX7hjCxNhyA4DvQc22nMglLNSeH2U
iacDXtdfvw5ixRHoY3DD1dRBF8Htt/o//+A3Tb13usHOPX4tAf5O6AMEbNjeRWgImaphZU4xNJLj
PmMd6prmIsTF9/JXn4SJupS3cgB3vWmX4eOLWGbtPprIqjpRI4BHhasIaqGq43AW5uy0JkNn9pS8
Hy0aoqJ1Wvd4fhjW960wj7gbCYD9JKVvqa/o6YW9k4XuVmW0qhusJuG7qJIb9sRIVX9uJQ65wSDl
yCdPqgHF8fUwDazd73QAKLiUIX6GlcQgbsiRU2pGY1sLuf9jUBFiTNovZUlv2Da1t/gT7QcVjgzn
o3acsrXXuihd5E3mUB/yz9k2aGHcHfH1/zhJ8T1kjzvhS460HwbcLBuJTiPiQ3uPzdflgO1XPTn8
3V1NKY1/ZkFIWvVb3ijeywmmULfL4MbTEWHz6zNsTK2PQkUnEyiyETs0KTm1/zIJ5vkLrmQfCEVL
pxCP31gGD8MVS/ItXHOM70FmjTP8WlTasIpSfIvdwlWUk8sRgtkOvHHx1bQpun8DA/Lv/ygg9392
+hWEQj1aR0NN/zQZTw9MJLdxt3oPUj8twhT7fjSWr6zO2t09IkOLfPK2Ubm5fbqiUUm/dhGQad5a
wvD3qoFb6PXH3J+RoosiptNIDHLSK+/6y8gLXD82vwV0GXWocXi/Mh3Pgc1wkfjv7w/nx+wfnESn
CibfEektBI+tVbR9Nw7e23y+jAWEFRtFz90kNfnSTN7K9Rj6pj55h3mjeNfyZiGDZK5Zwn2XJtv2
WmmemKexKMyMrM2lpS2jXYY/vXUFVuVp7CSZuHg8p/KAhVb0HoU0grb08N19b+Yhiz0usFLLyD7/
d9g3bJV/gBglV/Coe2ZRsXt/vZ0rzV0BmSKSfFiuUuNUmY+X4BgwGkbiVQMQyQ1wyv3Ocrp+io6s
9n0ARuH/sso3bRZu0xmEB4rsaaBHEgrH+RDPT3uASb3WQAngyjQD3MTfn1bDYN6TzsGC3GMJOtKv
veKkp3xSNFw5d1/aPGnno/3GDG1yK3prwKW4Q6Rt2SpG0yYARvOABR7IOP5GqGrrC7pv8qSa1apR
leXXUVmRGE42Y2BqQNhywdVHQXtQAVS+49wjGL6LtJWp2u7JyGLL0w2NJ08m+Z/7JLmtrZr82zFX
su1ZmfcQ8QMweWvhQnleSqHgix1pvlOKxie1X5F3sPQjd1R6fnLojV7eV7uPGsm/ICpsPkFEl7RM
MHC3X3O/kTcZBxgtL69oJJE3FCMhlyBTOVxndeKowzJ2R8jOS0A4hz+eUrEuDPMLqB/rvxVLdyCP
dsHPWFymQOw1lN/0RIIs9LgtcGah6bbbTr+TuLdmt8E41JmNrZRBpUendxYFH7rHmzW2cDYj/BbD
8fLGg8MgJ6+2jVxSV/3xmowQVgfqdeTIOUCtDfc+2dcDdP+MMqxA6Tbvmef5a30eLlzFcssPyoud
02bFF2RBgXFGXv0kvxJy6QYYdSjV3GOrqsehUQSieqaYVapeWlw5kfc5pTTIBTNRhLTQml3F/OKn
Fw10+F+KK4NBglrgebMOzjCc3b8pgGIJkWJb+5crOOrY9CTA0JAYd42c4DGTKcr1Bk94FnagH+0N
shEdkItD4TtogWdEsZIO6uyB4aZTmxH6oTIo4WaOyQcfnNY0xT1OCZPrc0GTfkdEVO/SsSnVynfP
iSxHKBNQTydJqbTxmOFHgmTukCypNjVUrjsCr3ChMyP6eA4mlNPcn3lYlv6dguA+dCUnwtavt80R
835ojClPjkDXs6n6JT4wbAuYr1TGdOTaUGPlVbBcH5tq73CQqa1e6kNE16yY+Bm2pEyI9Fc0ElRL
HxdbFNk32rx2XVQyee1gomB54U7jgOS8htLElhyQ1WbszhWzYUPQhK3Pu3ahK0BYGxj5/vplN7KL
V1OCmH5DMrAK6g+JPokqfWZUpWIiAiAh86NNy8KaOMgMtEcfEvV282nQgdr9547tUqjl4nxEUdT5
EEd5+tTb5enMHXzpuWOHCFBNiMJynCwDLbERvON/GY1fGmeAivviL8AHkI1nDxlQRptPo13NGZo1
R/QQkIHFHuCJzAmZ5LwpLvTygCxE+4JM2oeFXiVv6ml5IkL4XrasErpH1FCENU1i4zwEzkzU7dp0
NcxDOgT/15JuWbwR62N313V9d/LZMDvVlbvQEf72tegprKccU6hXmNRiflr7UXCve7cOwzFSuoZO
cYyHfPI8QY6EkWRO54ZNbv3f923rXN4Jtu+x+iVRcOmAxKBKBSNPVM7t5t80kF4avmaBr890tqq0
mx5z5eyLbfPjYwmNNXjhZIoRkKEPoOxvhbtf/1GnQRcos8+t8cjmfah+2adSzVAdcoR5m7zTe9mE
we+DVPbwkuwe/85yxT8/U1V0WjoYoL4UEjAsEA82D5PrEJG5bIkxKRjzvg3bJf8ON4FMuOJY3rmI
tfpHhovYd2tE2pf4xhUKUdKCLQxPtqrz1CfQfNLvBhct6tSD63aJTMr+3KnA4jtOePSJA9n3qpXd
Nxg2a08mRYwKm101XftDNhji0deOPAysgh1mkvHn4ouXosOsWqfaKnVwc9BZXDrJdYh+t7WZ5YZN
zTgH8L29TNz3VzK9zI67uzlJ3TF+UOMlD6WZP/wDlwOWIshogauQIB4k8qNClOWhIdZcmYBvVvJf
SNsh3q+lfUItUAmbQOK1AQCUpv1Vg/F3mWlfOgFvnEb5bMer8jEZoQjX7FPEDad2Ijn8slIN/9qJ
0Lro+IEepyv2OAkbe+6IahxI2JdqiCsftrXrFFXRGkmhg/GVNL5bxDqKlhuREnkklnZsZmLFzB1E
KrdceLO3tWQMM0dNxXReHlEHGhMSj+g8XB3fzlV8OiDhH7XvmX1B79i0rE3mlq7/gDGonbIFREV7
kJNEoFlaljmI+Yn878TAYcXiby6Dinflw5HwTU7ZrflDAba+6hDUwcsV6NTbryCMDcXPVb/z62it
++M5clgba+BD0bc+EuWwvYBwzPV0zWttR+iTrIn6SlIpnKsJWWtGW9/W5AHBRpVgSlnIxyL3m9Cp
Ge3DouEWaZYAMhdiPdE0UjxaDEr1d05hjqDx58IAkozVssT2U6F2qGHxX7PZERZm3VNjKBUyHh4g
FFMbCRRCqyTaiRESTK4b57x+qh07tJtlqNmQMHTZGQBB69xkX+tPQ6ELmlZBC+3dQg34mXwUSE5m
iEp8STybwGebkOxVPpiWmg+g4Q7hwZww8q/qYsQDE2pYolX/eEDE44E3BVDwizdor7FOphBJeVYQ
qma21As/Kz3U6MXNC6Tz6t4jT8uPGxayCl6wqKEtWtHpWYmDzto62wCcGnR3oCGfNza92ELUC3Bj
fXzNirVjkD7wH6i+siRmHHtvHyrhcKR0gDPsC2n7SlU9Sl0Fe5NaaNr1rAEiz3v9TJDzjN85pBY8
srkNoPgZaCpYBNH/dHaMbsXjv7gCwOBD9UACTLjoGe3yqI0ZX3C9Pslq0mNZg2Xa70U34GBA8RUP
d3F4UCInCeECywDhXNuvyucSMQRkxpIq3F8QQfqFo8YJBBx4ngGR/m7TYZmzqH9ZuD5w7ZwhuG78
AWyXgyEkQ6mEpKErrIHr0MN/Lkv+LBym1hd50dQEpMlV1ewphPoTwc0qYXVExYr4Y94SUw0pS5Jy
WIk9q7C3DTkYYRg44EoopxV6nmmUZhJzOngoniHcQbd6zb1e0+BYzmdDhDZc8G9kYVEXGf5RI+CW
wUoFKe6VJHA1QDTkTC86ccnTo2hoiNqn2bGZZZvk0PH4Yq6PRgrCJbH9JEyp0Z5CFp8q/baDYyug
4NvXOsdOGioEMxjhVmqcylgqzhc+3+40zwicgHs1Uq8YSNytFSW17Xz5A8k9q5hRVcJdrEI0Ha5R
d8+tjHp2mMg8n0Oj19Iq3lrPmArWWdHuihMWzE8wlp71/HsVjaSbU9BZfrPWt4vU5//Pv+DS/LB8
Ns9gWBZ08SYnIkMcdibMpdwXUtxsVHFW3loytkN6s2jAyOIBvP9eF1MBYWCOg0gqRdvu+CzQF9Un
/qCtICOBclX/RRYu8XiQAJqdyALBylKKWu/yv0d/BcLb1HyvyFvZCuZVmeSfeGfjP3bssBSa1EI5
CdSiyaPvvSEfnxFpmSECfRhFYeD0P0E06T+7RU3a9M9LJE2NEMP9Jp9ijX87/UBhafWlxhSNbvXf
drm/ce4Ox1LKXa08oD/WPPg+jKFxDugSLIbYKHiTdtcQALQUnxoAsIFxmWdxtKHFn6KbxdeY50dk
S8MpGD/dfzKcvNqom+YrPksDNrCpHtZxAl0He5u/GS+URDJNBwUXoffxCsInSIU2HJPpLfw0TVlN
/dn1Hyh0+EMUIDxJz+kzw/35fe9krhtOmWjM4Y6OZxaAT4CsaTbbCesfiTUMnSGXXI6NJGQQ6n+G
DwFz64Z6mJ4k4OxQCk9cCQSvU3kYEAA7fxSyPUFCqUmIk8ZS4d23/EDIlByvO/eNquvvoISE1WkX
6JbNOHmapPpjYXwx4EoEk4JZGYupTJQ5Z24Z+wiTL8IA/SR9WH4y9TXruyTI/ZlLfg4RYPHx//Uk
TS4ll7oKb4lRGrnzhfaMYcls2D3O1V4vrGbEEneiQw/kweW7DOdj0wD4fp+YNJpxzQuzgunGlGY3
BB9E2Vr7TiWtZmE18zZOIUEIcYjzh9FLCzK0NZyWVSlMVC/bJUfF/1G5Tk5U40Hv4+SpLI/9f4n3
k2Seww/y9nHmn8/8Dj0vBpKtyi3jA4MrStk4OrjhKLwzbEUk3h193ec2cuaOmkmKhS2xkCL6QIsH
3PdMkn5Ng2KHKRJv3OemzWFGeqKhPBRiZpjyJB4h5yPH3R3JQp7JkMPXzp6Yl0whNSWLP5zwakUm
YQGi4D3qSzwXkppLVIo57NSEEk1mOoQkY4WjNgLjHnynQWGyDedrRhW0LKvvmZfOtzv9+IsWfElT
sUrMEtvgt4g3FVoRAm72RwDRzrO0+iymlz+7at94x+nD4cR5C198so6IX66rvM0xDm1jbmEvIgD3
eyWr2QK0qRmAskC624dLgMai8YyD/xvZN0s2NClxeiHclVqi8b7dJPszutfBjKJXWybYWeAsbhDY
Gq/U4LE0k0zP9v93/PsUBQjkXRl0+kefJFjADmexbhATh8J9XU29H45CovHmXlZVafZ9bNpvrPzs
E/Zt1KY/lrKBpMtQU7fGftdU+NxXHpXm0B3V2Cax6PN6xJU5XytHrjx4HoQK3Jh0iXel1uUlKhEK
luRtkoXtcc3fse1+mbufeSFCGLOblOK/JKPE1UlJzVgCeDCwD5K3HAN4Fxv6V6VErZCM5TSV/2tk
wOSVbrz/enV7For/Ios+SYaIg1VnTzN5+jTrKFOlav9Fxh0dHJ5DTseUaj+z69EVxxyIZqVwzKVu
kw1eZ/dTth6YsR/DWEl+nBFKxSfFUZjqOpE7fyURgK/O9JG3qzFmbhqAvX9N3aNjoPR2oBHHTWns
Vi9bttg5ZJVZ5gEJ4xtrwlz5ZlcRqqJS/mn5k0TeOHYyVgsODSF4o5ZHCETgxfRKujACswvUE1Lj
1TaFUkgEVnAtB56ULay1fy0FrEiRaS/zJR0bwX9w6BjLNcRm7leigZwzc/8pfWpCba7IuXvtHeyu
IFO9AVcvnkRAjjVH46yBtVmSV0MKAvSGk7aaHTAhdpEDQAOd5CdECgwSkVyXZMAHFCLSKSmtNPyj
g6KpDT3ucni+O+HWulzwHvTkYXZMcFlMZj2QSLPuqWirVk9BHK5emmgDQgqnrcWc3XxkTPeT+hdb
gl0MDeFAKOatnNuzrJnBdWsktuwgFJCqEDut7STeM3LWi71xuQgmGn7r5J0jXRp8hVcqLEmBJ6aA
4sfxqH3q1TgCM/L/eu9ogepMMcsnH9adgShb2UPRYK++hAm0L8hVBBtriUA8f8rsypJHvs6Ey1XG
JY30oxvzf2whyZlMeEcknEs+ICDKqs6BKf6N0W7WIja8CRuFhhVN2QFEeZv9XQ1bpTo8oXY9lhXF
3bBKM/7wgq832vMS+oEkKUxDve9JOOIJnzkBKOZuV/ZCc8blEeZXvRuArgVsrR7aKjFkW1E58TGV
KGdnv8AxLn1oMa4UtjRorbsG2AdGHB+FoInJJwS03LP+KwTMVn4yhUwcQonDT3v0rTarr0ZFjBSx
C3UQa392XKNgW3mxIKs6I9G79GoAaWE8KVssf53k706Dy/O0Y6DwPvk+GDfCRccMqTJi0qxskXk5
gxpoXEsAGcDLsXZa1JrzJf5zg6ynIVjTtHCAwREpszDIoDpfxr1wphSJzReeuWgpfGnIJBc+QpGf
AGpyQGNtrK+FsH7AOjaWmVgY520bCfnjOOeastEOSlB1+cwmQHy+Po+p117wUE6jFiejpAgUkQ5h
huWw8nagb35mZSKYYyq9d1sCaV4dYTXV74ZlEhxhzsPMIBR4T+ZKfO3wlqM6QnoIJQuNKs+g9I/F
1a0x/bqRKMe6jOAH3eCyQOUAsYJ3STm9HCf2s0gPMZTykDoJIjSFnc23IVEGEiHJeTrzcrZp65rL
/u7KoPGDK27r4/2DpeZgyhyvgRRJScXi4pXQu0OxGcEMkA32AqwY5i5x5nctGHK0br2sx1QLIuLS
JvSdYuq9sIxJpArP/rqYuvbLwRjdB5SWANHlzhCSPKO+kDGKYqHfA/ayYvjpkSZz4u2eP6DUJ8j9
PtedaQ8FYXBvjdGvBug+8G5do4TQeHNDCuworpBqzbi4Ls0JvRh3Z2pB8qaquXOiDgKPpu0pnl9g
QzCsb0Pqyj3bKTzhspQzgOv3gbuZ4OTge6gcYWDsOZfxnkdWEUbkBkg+LD4dsPH3+B8GXoghlZyq
GdOKLzfcf7DQUSubepFCRhuAIXaxoW8f0A2YE9SsWfRJlDZdMAusMDyIwWCUk9ERe1yXdPx5oInV
PkH+2/49xZtUmG/OKyDa6yA9aqABQXm7n0wf9MM7LPEZBdQW3Qb2AUcaGLvOqVTKRXEcoqwVUwlT
YY0FM6iK3ZdaljrZ79gf8wmZTINMB3fZJcCCH+uBHCcHTcPSvdfCpYpy8AweeRDDEw1xcnQxMKA/
C+zrzKB7p/MrwtQOEJtn+xaCbZ01J2WDbKYq2dTKaABy2rOcv89G8+v7w3Q/DhVkYkG4qXtLb2V3
A4r4eenAZPp0xCzMUMXW2v/wUbxBSVq+i/kvY8QAnXSKd0PQAAHuTirr5DRmJ1nI2U7p/3QCS7z1
uDnN0hl+Ex7lWDwVyiFQUzi/gtYXWijPsTQdF/sDpNC9J2gxuAfSmPEKkJAMfQ4v6c8/MzK9Xfn6
OOQrZk5OcH4Fvmk4pUSXxE5qFfQRNKwCtepN8zVx4/tOQhQub+UkHwBbQhwM35ai3VgnelhmZCDw
wm08bi3cNJsEu8tt/XtbAd4YA1lphDAewjsRcj8ErSp+rUXc8nMDsZcdIVn6RFnJ/fAsPyRX9Txw
GL3jPEfJ9fYbnVr9GykEpViTcgwnRX3ExAmk3xAt8SN0BWQjoVR5JbGl6LDDKYzkbq7y0b2spuog
mw3TS6lH9iK9BHF3IoiSvpx/RTU2qiUs6XV3vf8UpgdJZQ0lnu/Rc+UubPon/Jw2YUKsV5m5bxgF
e+M6WfhVuYa9wQeSVNPDi3hXgOtMJSuqLYGQwfTI1dbjFMC0qYiizJ0BVJVrhUYmtKqVYx3Lxygo
dXWUS2s6oUFm1hH6xB91bdmdCOkwki852hPOgqU8NIEA3FBWYSH8i0sUUG7TEuZ04Sk2uPpJEed1
Ih7DY0HERFAQS6ZlWEEdbQRZuujR96LQeWHtzRxPAqWeik0eePEt3mheEiE9nPmYtCfC/4jslZgH
RMfM4XZq2+Dbt8ZabcjF45sIKG9jCy6/M5E1KD0jF0nvzsaIGO/UlUZSarbfY2pDnLGrh6kwTMDM
MnCpJJnULqaaqzzZu2R4d1KsrF+Im09FobRbi0wNWIWb8FH+Qr6NVizhqUC1k6tL5jg5pM2vHNW+
85nS35NGQlZbm+WQMvqYKdtSqxHfBJt+YYMrIGGYYZdYEo5hYCddipaCsvYTtAYwkqVpp2cQjDte
e5XE1OsGVU4FzTO93ArxrsNJ5TF+7B/wOLZQuu52bm/HXmBRj7hG3oG2+SsN1HgeL+8Zs7u82qoJ
/yEaf+pCPHaL12UYBwGJN6jOHGxVOv0AMMoIGGVU02fTma2Ljy+0pZWM8NgC2iBg2vJvC7XSNMWa
xeu/U8MgfVbqI9h1gLhU5PITQXoI0PJ28KN5GCIQkw//7xIOcX6ZJMzbEZIQXDLJlcyngss0dR3b
3Ef9uomateTHIx04D4B4Io+v6ul5rIkuFOD+xakb5er81M7sRL/9Na695/wAZDKOLyfRm1SMm1h4
uaOBK0F0TaBCNKF4WAcnp5Duio0tzfGTDCy5VKFpovc1z2dHjlwh9kfZZaXUbS1BuwsbvkEAm05Q
Gv6xU/a53A6YpU31uUP/3Y+zLCwMWEjw1Yh11PWCZlH1ugswSiZCaabo2LuYot637f+HUngfkNOR
8wM/8BWyBStgN0vf1GfQ7dSbgx/zobAHC8kjJr08Q2m8Iv9/nTWRHaHjHJEQHAn31mtQ+kG60YwF
kmoxnlREfSgUcFyxk8p+gAC0SoRcQCbqm72B397xTrtgSGFh4Vg4k0ETWAfKITl5EOkV7ouwaEC8
LCfyXu52GWDxwCJsmJPp7ltIFh+Z1RRtxoQK4YISBmVscP+DpA8GUGK08U7CyygREjsYDq0b+ugX
iMF5q4s1o6IYQ6R+G69MSaCxzkzXlMWdaGApKjuwUDPeAgEmvorwkZhmzPkxXgRzDx3QexMXd1Bf
kDkOogaVqwTJzx0u6UT0r+20+FEeAwChrghsRzwscWJlmUdUUlYI/1uOnroj5QMwg43MZ1P62LAb
peoGyM9oLYUta8RVBA5Kv2QcdGHLcL+Xmn6y2xyUw0N/dPeW99E3hmwq7fFG4G6WnCzMB4ApVE2M
W9Z5xOvYm2zQM9lL2QY9QdHauwRnQE+3RglY+fskUOHOKNUd5GyrkfCLWsPGRdnXE+c8Iuv87wvH
VuiRj9CCxUYDYDk5HO2o9gmsCU7f0aE46aYC6APJXBfCKFHvw9+h+qduAptSj5TNczpWIdEaFoW2
1/4ZjszGJHFQpYTDndAIzBgNeqxwmYoSsYHu56ZZNBk3AWIUUSbkVc+9HdqbrRNgq7zGIiwqnXEq
4Fghb3y+GC8D6DwAcYxbi6HvKUuMY1wBKU//OjLlk63D5dP79ouLLgY+mqW101onGwC9pd/rZOHA
M4oRMeI6EmNurBpLlw9P23k9K3IqP5dxWLvhUZZdTGf+y39PS8ID/XybOZs/Z1J82HMkKbJ/JgYm
jGU7PjaXW68p418RpVibkD4O+oU/J5+NlkMqcz/wIPjVMgi4et4xmPR+eC4UaRA9eiC7PUQLnoG5
o9wXgDDRLCsbORLkPPjttIZq4KFxKEK3t5qMBAOSN8W7mStsf+pByt30QVdOQRLLz4yqWneFUUZP
eTjh943w80B0MMEVUFfQByafH2diae3ppHM0CBRFp0zxwCMBS/dGDUnxyCtko9TF3Trc34SOPOPX
adsmyVqZ19MikYKVDf3ALyWjpCGnhu0H9dQ6I5MpnkrE82999ATAF/TeNCI1Dpl7ZyIXaiqpiH8a
fD2Y1X4YMx15fqfIkPVqUHx8IIHVOM/nQrZeMaO3eAfR0gOvkIGODEYVAsb7f55kfpadVtjOCCyQ
tyLTv8TltEvS4Vm+2rSLt1uvpjEU0tHAgqX6g6JTLZX47z2DtuwHnKzKIXSmFauRpp/4mEdrMgg8
AVFUl+iH7TghUVef1WStOpSakCRICd3B4KvqW0yJf1tvASxFItbnJqLRPxOkwu6PrsjtEFdILkhQ
E59q9ex0hlUF+nMxbH+2nINd7HpgmTY4rsyVmuj2GRQqcpUAFTRqxAXeB0QgoAFv5iGWLBy8Tep8
YHzpbwuiX2PROYhovM0a5VLmA8qH+4dRoZeGSibrCEu0giauDNp1H3Nl8qhoUTVzYKs9CMytWgmR
v9H/2g0bFSgPkTDYI4m1INxvQZ5rsr8HI7aY/3J4nJrvF3C8a7YsBZ7dX3Dox+DP3yKwJAkglyem
5PQRQ6Nauaw1MCVfIlg5XwjRm+4Pa8Xza/bJohFH4OV4LoX1n4agJfS5iBm5SNh99VF0FWfeSinC
S8zSomdQ9lTz8EYlZhQD4IZeRQE2HWjq6PxmGppKjyRzES0086yqRRVbYcIQqr4aILpEt3N/MZfk
WVUq1CxXJb68jG3nT/vU4dNMAqx5emz31JjtMuuYA1TIfiNXqODHIkweUTosespTx4M+BImu76ay
zhNAqz2Z5hO/Nw9UosDzfFTc0gwmlwikHZySjbtyfXmQY1TJo9HjqQxnwb+lAP/FdRwyM9WMktpb
xCdf89/MoHU7Pnj7gA2wlpst8fwgACUWmci5IfyH+zj4YBsNBSEJSc08VOBp0EffxI5lWvxrCOG9
OeJI56pXRpFbd1vtz1zY0PtV+UTdMdj8Rhn+8DjLqjrHiUL5RjrJNQuzucZUOjNUrnmspproIYw4
z0b4avQi7ZeqwD7Txvu+JkEaDgy+CeAljPG6gAJ9c1Tut+5sRD6R12DzRUMRXdasZuzO/FqKDwXZ
CynaU4Ec81oIkb2pJb0uCvC9PxIhirsym3tOexeAKM72WZn2n0FtMqkgMzo5d4cDCCW6uMpGt6v4
A61grls5zmcqWSEVw3JIoJ9a3t0OCJTMkxHTjgKUT6MI1cji9LQM0t8gFeiMaeFf21QWVxFqMEav
sugT0R42peSn1J4CdKYnV7BJbAiVNk324akwfbVu0vUZHjSKy09gQ/qx9y35f82BdYYIJrgUNugd
J1oRVUA9l2N/4K2BUQFtk480784pp0pjMX8Is3K0kif16tVjvsTKywfAw8TXOD1UppPC/KesVFQS
XdcxRFEpZKHqH2tE7QjkMuEuVDIlNun7F46L3y1aTq9Zg5nTWFfcvuEvnhBY6vee0oeZGwqjjRSF
yVMlOCSIIaw8dNBTaPnUsJXsb/0NQz+f8SZtqTK8d0kNNQIghGsvkfsydYMlpoNoGsskXjSkYdvZ
glYnIxAoFrT70t/uxFTEE7QTDJ3O2NdBJdtIFFnemKJQRx3b3BQLOwrJRZWUH98IqF7bf1UHisgX
s+7IJpQhuJ+qJzuDdO/R6d9opFcTd2GM+U7cPkCX9HhKcKu6mNXOR8+KdIbVfEwCGsr1N0aRUp0F
E6JaIwopjkBjjKFCRX4Z7icb8QDD6Y0Nd066MtaNOiWOOww/SIgwJU9m+X5+goMJgNKs+UbNYQAn
lHsdzG9uXK3oQRqOM/bTnNFfAmDlfcy1t1buhte8V38f3JbxkgjfnAQZNZNRlcKnWjcV/u5dxYlt
2ol0hhBNwr0lGMwsCcpn5aaNGEinKl6Kbu2FyuSteIELDtNbufbRFusJio+vjOX2SKJUAQhGASzu
KFKZIvsTov+Sjnk9UVJubhx8y/eEFB9RD6L4zQ08IvZQZNliSSW4ktw2jfyBbb5PVfubxFQaeHHj
qTMLIiwynf716cpzrdKp+G8WZPCbuw3q4ovg8B7LX3QDK9T1zbGpIVPlkPRuqxJvrpb1CDKfeFR7
WK1Ne7ztXNkvPRx9BS0AV6YmlYwWFu1c9HHuIgzB4IU5FZznDU29HDpNUSWT2TU4yfyqb7i1eEaK
g9vLE1r/iOzh57A8tu0KX3CfJgFd8G/AzTDlh9tOefoIG+DxGngVj3C6vjgdMfw7qOQkZechi+HN
fd9X4Zkmpds+PV0PXHBQRh8A5WF3YFuBI2NBzXTykOx/xYPm9304xnfU9usSXfX2MW8u4e56BEnA
fCNH7Y3P1WY+/Wv3hcoMIWuM1K7OZ99mnjVMYqCVJvEIL9i9GGvt+piDEsrFH4NafV/5rJGqDFJ9
ErnC3o+tdj6PUkgnscYjzLoOE0rmQKZgaAHY5x/C6YO7EwHzd61p9KzGnII3Vl0PG4DT+SLYyIjF
11b09wP/qfMcRqdSnje5ZLXaT051Zh2t7FHCuBiCKue1sv02GMgKA7sFHLvbi3QcxSS405VwQWfN
HQen+FO/47QxfLwjPC7u9FXANSaUbveVKly+pKaon6s8Kqse8h5PYAqtZH2bvT+BPj1THAwDRRQS
bF454MzqrrJ1n1pzD5fs9e+wOTYF0h+hp70Ahug1vkx7baoxVS/2wnq7fWtxC/cZ9nfq2w759he4
hsebKj7gXifX5DNRTEaY/R3HRFdSqxwwGV7Qlu8lNbVNXzV7TWJBw4/nVboHMavROGJlBxmqitVK
Z0CTTeTuF+PYezNA9FXtFHMREGfqUg0ze30mvJF9e5YapegRK/xDk8sQy4Xxjro4AJrAkmCagxdU
kXxsKwsh4jxTGcmkXWxrCzEl+gN1swrxRhwHm/2MgJ/kdR0REl0hmqunCaDPVHPhA1LqlfjkT5L3
U0R1KTIL1VMJcs1AMpjeWx1Jg7L44YHQMGEd16x++bLUIndlkbHHLla7N+mXoiatDjCk+k+9TYCN
GrREOsKSnely5ItWZ4zoLfOxWnl7DA7viyH8q3/TcxxbB73CZ9KqVV7m79yBvnzFwMJwvFXObqmt
+0AIK97x6Zs3pgL76V0Lnb3ugfdmUuti3Uswu6194QYHlsj5PJOZNt6rbkFGMrfNVRC3iQar8Dl2
baVvNJ6wOQ3MqoQm9exm/OXh9pVAUQrJLkGJdlfaqYPZ7JSfQKnFiaSjMSRfaCREpczuktUUpeXH
DSbKiq524Rirrr1czD+igLqswmBg+ROqH07WyyewDaR+3EpyaSnIrhIYDNrrKDSgpU9Od82Q040r
W0TnPduw4PpiWXHDTdOP9jlmEbF5+ZVTe4tFLAyysjFkVLTAhbRrdgdQD2P9d6r4Q59IFyAfJYYw
QgwSLKs4nNs31tgnFb7xb4AX1PUFmWfYDtqH65Axh9AoI00hxtnCHDGdBxC0q/T3xjtxK0IUYTG1
M/kYAcZaipYEsjdU/vKTfKHXCmVAL9Wf7Sm932DFLukeQxBA4+kv8YZdPR/pqson70XVOMqkyG4l
U2bjcTFJ1UwY7ZHpvyRfRVPAbo9TDboxtjQJXinYwG13KZzBNnRdSM6Hi2FGpvnkNVXT87ap8uim
AKAhThvZ1NbvPKqHqphWKuy16Nv9IzjNgTVypS0hF8ssviHpeIXxbFCUHwWjOc4OdBXPqrJrsUFu
0gH/lmm12P3gQpdtpJbfrS5R3WDvURbXzREWuIXPLqwniMHTN6dTOK18fY89VPEeFqtdbTn2cmGw
y+jlapC6zMx+37hfRhSdkmSM9ckQCW6QyrZQYWVEBsUzh9T+zPR9QsbbrQXseyEwYTDDeeF0ch1i
tPl6VJKw0h+liuV8MvviREOxrADWbdL6cBn4RWgNkHSRm0P66uIwt/FIsQkSScVV3nkk+yoakygt
3XQq63jyFtWEWE8T4q1oljYgbrWkluXebbXXwa7ICVRf+dl3aA10ZHRshWEYhr/A54bZX4qme/fk
pcvdh24AdAgfll/Jpa5ZpA5Ki9qWAlpxddSkIV+vYl3lr4AICV0i7S50eDgx8b5g2CNNYjkFQ4C/
39D38CtpuOPyrWlNOFvSqIe7qBn/Qn5fYtiP6mnXN69pSnZseTARDz2uJN5Oiiue4ZQC/ukS5YVG
E6wQwbCdeUUs0Jgx+NFsqWFwiOAXiTCgUEt8HORH0jXYrW4VNSdlZJsyW2CQpYRA1sX3q0FGPb9K
V2fPTICMaadkPA09Gnx9TdvkX+i9bNqSX0dXbEOUPHZqWfw2vBR424gyMQa/dPnq9mIZE1DqkDti
lzTfQ853HcbBIYymo4fvcEYiHYhxsv5WLQLnZ7s/Ev+ITNjHw+q1px6LD2iu7IGDm4w7xugy19EN
dUy0G7OtK8AjjzAmVz9M5BI4tVyviW/f6b8q2Xn4QJ2rCMik0qrOKbsPbiAuhXQ04Ip7+h/0q6yC
epDU2EGg+ZnWplyiGH5x49bE30o1+VLtU/d/I/7dUiBrak/Ewzj07csCqMLd5ysWGX9Li/ypwf8j
uodp4SVaaHmhJCRyIOtQSAMuG2y7NI5y61z74nkEBeZ2z0E7JC2WVetNmhvLmsesdAt5tta5cBO1
Xr2hTdCSc6cCc7qHW+ocHAyRkOy9gDNWM/MvkAKwd9GWEwE8hdTqrZjtJ5pZFnb4aoTT1V0n7jzJ
c5OKKZaaYjNhZN71YeBq2yb3ZfWiP3A2M3rHPbBXv/+D8LjKk+/Epz/IZ2YA0uvb+a1s86lhAq3s
UV9SY9P8j3hTOx3bORi0Id66gSrSNVP9ry4Uaw+kKF9WvU0AXAycYcYsnVrQj34ApHH+P51DAsJQ
PMRNSRujhr9NU+G5H7tJj68UBdO6P9aXJ7umkVfdS8fzXN8rbKFGKO4ZPAxi8/K1c8mA0RyQmIIb
Cy26Xi/Ql5r1wwwLDLV4GBhMUSOxPwBgIzaO1ze1whJSUZfobs71T5XxpEKBF47hLHQrqratvIzE
kecXOf5A5GEwYmC/McWDijReXINUpzNPTdzeZ8KTmhXb/a+NJiSOsqfbKwN5gD9QFMGqQJmgpLcu
/dhvttBp6P/w4XOCyRlYRDs527yiGb4AtA5QSAHVGqchqG2X32xTbUP9shnfpMF3omnOOC55FoeV
Qt/DQYNngp4jnprwxmu6LldTstNqP+llgs00l5eQ3XLWWT8sDoVhMGNhM07+Y2EcXPyEUwPLx2N+
vpMsQ94kJ1TA+yLlmtWNbVOybhq8vBr0Y3AhUKnIu9amV0jAzzWGxNCZImQtLluAQPdw2y/rOsPt
X5wAIXwO6GKZXhiP5MyVAqpU+CAMjLnUECYgIshrrzYqMRjNlourEhXdcqD+qsiprtm/Q3B9i9yU
rIE4ImpbpDphB6zEL4K6n5fwmlEcQonUtpbhz9Js+eiHw5HwYRm4/Ru8AsMGHm+/RzzRKh3n3jMh
uP4lqRAJJpYqvEg9UqputLWxw8EzMJ6Z32IEBvAbURBAmc/qdQplYJ9Bw/rpL01OdgdE2Pkdr6hm
7fLssFxJh/mquYRUekr2HWt6j7qMFydd3W4LE2wGaLtsB+jSqg0NAuunrtf6LqQEJboqO5Qmp7Ip
7Ed0mK784Pa3znTKcWlN053YBn1htLQgkX0tawiDIMJdppIoZWBLrseZLpawFLpL2LqbfbLdXuhB
nxcWkj63i1zkcAS3BfVFQ+WYhhg5HS6HsvPPJay7QqGO14sAqffNyFeX1s2yZOriOxXjQKJk+4qm
XGCbDOwJQYoUXg9C53biVcy8ub5z1RGfIX4iagOUXREx+BN/j319Rd1mdN7Rs9mC9x6z7+YeYEGn
Q+rL/rtOHf+OXuy4sAGdGpg9QfHg1yiFQouZPf23neAke5iExxnvd9KdJVBB3fbtg8ItPbEPRBU4
h6Hwc7DJIVSDWDTkRDSfP+gGi3lqw88w34FdyNX4QlPTRPnt1BgAb6PVKEE63wck9JnGhmOL7qtj
OPhXYc7NPQuB1wiqAiRQZDwRh31QMYWxekppdZO1AAMKnHUlvo9Aa5kkjo3hm6ziHbaGP2rh+PAV
OZL5pZxIE5t7xCkc4wcSuAnhYHtTT6JW8uKHWZCMzkVZ781W93OIBBHX173NcmfvVg05m6fKHPIx
NjyZvvGzjHHZ9IasoKl4thAhI61uux4lKjp6ft9Oja0/6ILi9cR04EOvvNyo20794F8FfwC7ExGj
LF3n58xdGzSH/cDvB9NgHObeNwxrU7hI0YtcWbaHhdq9Z9AKXO5kDw3AZgE+tKhuwCLi0u1Xf6zM
bBXvguT+IpgTdohO/EfqsF6/yTNO0p8QL3b0GKbQinHyRKGueNlaRra5CrRjhZD6Li5oJYZ/udw7
GO2rL0LodRlCC2JD7KtDOJvVcyKIdqGQzCvHVh95SDTpzwWCuNHcSUHhnrJhGxt0GjTN4vvLW1p0
AiN1ugF7focx6NTNETFLaWdRFnjgKHPBzSCBrJeeGgeXpqMnq0Yw+Rdw2eirz7s+pvztrzv+obW1
rwXlCFvr3KFvK6HA7RtM1sgRTmB0cL0HZH9+BEtjris++NC3/wRtuW+vVTdGfnHOoHrwLpKcLfIH
HFGHbfQHIuT430X08jTQz3yxKIaOnBofIDpH+73whj8dJY7R+XdPutRb9dQDLN3MdCXk1FeypqIf
WNPPqFOQtwHUq2pqwF/0yApT9HlofcsP/SVfFHy5X9mahHcc8HRP8YFJj4dkanZ3IA4bRZl40SFt
hD/ELhnqJxHwsJAMSNjEO32X7Hv4BvN2WclZyHa6nUykGiZ6+tWaGdvDGXjIWGqS09a64MGzzUHm
QQFBiCrP1ZoI0TKR7jLfBu4FJUmzd3nScAJEfyBqj88xPBY5xIY0RhZzi2SghA+QBRyoDosfujZ0
f4m1fnWAAWPrCRwCiDwOLZ/AM57IDG0qAO5T6qq2u50yaMGSc2n654SwSMyu4UURnRQiiHD32h5g
5/UVrdDxbzFKw0JVCcevrf6+mau4II3khNgPPH4Cp2auXuEHmjkG+sZG/FqJw0j6J8z5JXg3SyOl
AknAHR0MHGRU2LiglARNkvfHbQ2sPiDjmSD+V0Ty1+Dq+Fk7DUVn9QZC88+6KsA2RWjlMn0P0XVh
PE2DX+x3ldDaL7l8rWgp3spwedcvBKSGNpLNOsH3dG7oOZ/6I6h7+hphNRq0/aYHnHG3eJWXHHb0
OR9Ew8r7FB1RyCjC7pe4O7dcG9WVFJKI//cUs2jCmPrGC0sJNBtOUelNjuRyWmjPngn0lZW6/F9r
AAduoE2y1THG+3sRJthIQsgpQ9fRaypE3k8X4F3Ikk651AbLCzYTig9jZhH9oEx88Z2vnyr39vYF
9P49l5iR6hcO41FL2pNMlBifxpoLhOaS0ArCvrS12d9xTPKbCOpyMMI5v4G2iypymBYIl3oUiw+0
59VjjxUVo0qjVahAMKLNwsWikqHCW9Jk5m4Nvc/GRxOna5KK+UumWykqDzyiqT9Wj0PNv2boIo3j
9+vYXtvK/BfSqdI5rNQqw+pXORZt03nZVC315TBTuWQcceK33m+5kERPHtYaKE5rafv5lrr8y8cv
pJf/aU+z2ahuZjmT8lx0r8GJXJ+yAVQpWVlXe3sk8f+vn4gt4+vQFY034uXjHNcRLeD+04zGGJyv
rIKyWXTxY7VerC3TFSTMEQv9lzdTmDLNBaD7iDXwCuFqfgw4XzzAOlNZr3mb++ACva+KXiGaw/pm
GHv0DRDJjNNpDitNPKsiuJIEgd0gnS0d5IY2omyTzSDxMe21mjcQtZYaSj1hxVx/x3iu+tJKAtfA
5sZRLYOeADn8BqiL/iXjDS54i90PvD9v5/HO4O4Ap20PtphIHYyGEYO2zeU3r14vlhymq5AfEKUI
by3fqZbR4PYYnBdx3m7CEAu3N/yEkvSN6HkRMM5VjU2VUqEHX0eFQPNu5IeaZJCHKk5/aToOQaDi
/OxHy/uTcKYJVPTjqMOFkEoIPZmtYyo+F/9U8HBnTKMX8cSqSe2PwIsQbg3UGxXkiSxfxMB3mBI0
X8J1cBTUvYfpALezUuyshoIR/JQAOJxJjcT6ubPsFN3vk0tjosSiasf3KZ898hF/doYw3BaCznnh
lOUJ1pp0WXnXf+fZV7Yz6dtAi3AXVH0H/k3K8dOpDGbxpnstTE3uCAQydS+p6nAiTdEqZCj8KMOY
Dt2WBf58kJZri6k5KFJ/UCQAc7sp2PcL/2vDuBV86Ylj3dWCVWrWNeHvhZwHqRQQc0NLfWjbrV/Z
RPXwxu5AQBSfqPdcj2IAVhy/shpER8oOrGoJQCRIN378nKL7T8WS+Lah9oBppKY3qfYU12d033HW
oj6Ok40GArP0IZqcDhaWrC0XN/YyExw6KC4Rx4fpoT4lZdSjetcEmZLr1xlPhpplSy6LR1Hku0DR
2bmk/dGzdnUJj/1w2nRZQlfmpIQ61diNsym27hbw7QGBh0E2zmDqCg9wLttKkgZZTA5qPU/PhXM3
iVeHULCkoRxLadPzLP/JfwmQ1F7FZUYF2gVYhKVAnzS30mQGpiKkHIKAZdIUR29FAqJ1Cg7qWP6g
/ADIAwxu/RZAvjgdHqYp7S6ylr2KPgd7ed2ErDNDumeNri1UrZs2YPflUIaaxh/w/WKBBb9/5gi2
TWiYNdaZ000jP+CoUwJrUBsKcdSIfd03jXf2Lm0m/4J5E67ANzPCpNbzRbAvM58+SZfK0Brk+hbQ
sdlG1FtyKxsMar0SSVfTGL4iUlRBwBpJuPKQU9lwZr7NT13+VqrZd1OaE1B/Z9rPJCiQDaocbzWG
dW2J3E27I8Mf+ft0WbTPJNoMp2xG053xkMXqDE/HPiD1dTW2+jLhsQYhk5NIn7pj+YEHDwj+Hs9v
44ZgjBiU8NL5AQr1LFBZCVLR/5l5kOAiU2OooqIsRsToVt8zdmw1fgy+HFsUpSMsE3R2goN8y0kV
XqULKGeQPNs6hkPlsIQxr/m9cfUxh5QN7mJ6RowE+EOJCboLY4d5ISYPY0TD/bcv6AnnNUpkca1I
3bqAcIys8cyjE/19YlkX+IXPF5LdpY0Bo2g5iGR2bdUxNu1QUEOxLHUg+ekvxxTe4TdSPzmmEpJX
BTr0MUb/eMlf/Osw+1o3g8osiL1DM6j71oemolqvz6GAfbCbh5lAvrHaZ4fV5jpRneypLRaTyP20
NBqM4TVCeqzOYLKEEyr8WBbMG/wghtX1PKmFeh6y1NQy1uVZWydF73KSPUm6QIjn4M+yDwVE9KgJ
NuvEWgSS0aqM/b9N2IEHuJXAipy6ouy9kryfPAT+Wo7ElCaaIOp7FLAcfdFrWYCXi+a+ljXPFMkL
Cj8GNKOBggHgfNRVraFqPF030sJiT2J0kEoEvtqOZkBcyA+2dapgXv1z8VLESuSMVAUCj1JCRa0G
trVTQd4cBT8bJKtVZWWlxbFCAhGp0qAQW5veJcwEQhTFjLXqttwNARb8fkNvr+zyA2NmxVjTDYm1
x2gzYo4Pu3GPjlwY22VL6x5Kaj2ofxdrLHgoH3QRQmxS/SZWAP3zT1AjKs+8P/qPXsGUMizVXtDb
n0LZ/UPpcguBf1bsQERpM81bMAf7j8889I8HaVgsTRSkWbiBYfSODFm0/w7OJgfrH2tyNnzMPavo
7FurXMbHvyiAakaynOz3MdOdwtIX5QqvLdLJ4QK6BLzn5gWhgFZCXx9jHAbkD8QkxfiSEg71Nr/a
fYeizLS3+BmDmlj2zYLstZsS4XvNspfuyutqihmjNloLzqkh4kaQyQK6aWUKwu2MVc5mlsrmoNHA
YQzrCVv79qt3UtV1QwaTO0l9pFh7Am8EliR1LGwBkDTcdsLGAdNSe+mdr1H4kyHKzAnDkSfsLqRo
WCqRpwMVGJQUqKmeg1lgbjD0GzLUs2j8aY7qHvto3kgyrTRIMDAta8Bz2M1c98gKuHFZDiuWNeOR
mvt18NOASaOedm1nTZPUJU6252tgcSz/fM38yyYev9gQdEGnZe0T7AIPNAMTMn64Do4l5U1usSCx
JZ6JN3n/tvJtDlJNur1mdopEs35Yni4evtVu0GZM7puAHNVluDPLd6i+m85s0m0Bj5/PsMhKBTNS
TNVSxi56abCmhb31oj0K7EmPENDBGBJruuanufybZtBnwRtN7fNzhWuy0yGctiTU1LZYNkfBrjGX
xVxcOptKT/ks5/+itGVYvm3CYG9EQt5sPcM42brJi69tb2of0ee7sBDj9feJ5fg0X+GzL0h/zMKA
qnAwCwQa6qSs/fp5zUlqmsRVT8hIsO2NhMw+cit9JaCAw5FG1Caepdv/8vjHGgK6hKYElzdbHEIV
Z5qf+KnMagvNeyGnsQ/C4+G/qgCInzCXh+o2dDLEV/dhYr5zC+lK9vQoLYMz2xz96QjSWMdn0cNW
JuzmPG5hFORejCK614b81IyAwQlIme1DhZ2yK+2vC2hIi5Hd1NYksdhZuuFsL12trODoXi3bIV3M
R7q9mcvOPRieh2hbDa/ZXleMRHM7AMNtTWWdshpAB29QAiHVkfFVqLzSSN6GKMUOBNWtI0arNgyI
fsFdxhKKJUK08bGfppOkL2aWjgv6cnQ6vdwfbIMH0F9l2DbwJqX7IqiZS/30v0hzF7J3uhNaLp/H
7EdUHsUxrwigivRF9UOVjrbStv9u0OpI++as65bgXa7Ba7Sgf4Uo05bfFi3eUvNKz1x9TKSrrPU6
9A/sMQxkzl/ge7WD7TIX4f2F+5jBNGK2KHVQHWUEMyalieA8NkE+3Uf8cmYHKSVF9I7knP3K1HNP
veFg7f95Vegy3xvE9ze5t3Y4ufDxuY0dRUQz2o4JAz3PFiGyimFbvD7VX3eMYcokJwwRoHr4m60H
j7jyARUpg5qdaEUEEmXOzCPxTWgc3NiDyIbOfuuRPq1zdlhqRNiMay3U+SnCfDExX193ao/Dh+m+
t63RaRxfdTm+oRR89PVif+foIgEz5Oq+2NhSJQEyZ2ecN7iVxl+FU578xKThxINMYP4B5nTUNFy7
GP0b23iHRT0CdhcoDz0/M8EoGjchTVhIHcPgAJkB/1Sd5OIuLqc4iQUbigkKyZeCnAb9Rvg+zV8M
k3HvP+6ph1V+X7lYWrEVFfXHxLVn13WG5lLguPKVwr/SkqkhqvSmjDPaHBLGqsxBYR4+BJkHnqoG
bkEkKx47SeZnKEuMrbZpKsq2GCGM2Yms2GUFReF/jAfMLRgnLUgwXV0NHKTBC/ETobD7zAf+f+wn
bMMFz67Vrf1ZWFc3JATQaWdkptiFi/ADdHSlGY3brCG+MDOh2BnEA1njcSj64DzPb+STHugIQULd
QbFzP3A7O9CgrMTLV6BcoMkzbVEFyoz+xvx49v8tLPtCQSl5PF0RQwL76pAVCRZSuzWICB/S25Ez
g7mv3Xc3VX4q/LUe67ucT4oDnkuUCJbrdvSG295jsMzXYfYQHyx/QHyPz5wB72RTYDjAAckq4s9y
l4zG3TZGk13Iyak2fXk8QgepSaYak+RadJHskWgoOvOeMZaTy9RIXY/VAXt203YTQa6DMAj2FoBM
yIuCqPhuVVRpwm7u8fUeXQsfNwYHZ/N6nPVt/s3+CoSXbwdL76oIKpy7fg0h8HGDGVf3TuZqjQ/R
6nMqjijFVcqoXdfoJYPrlOv0cXYuTEs+PKwx93qStkMPAyhqb0AxZaAOhAvOVWj4riktdUSr2GJM
BRzM165f34HanaYXk4bJ9OSma18+HMBu4Y9bULfOFWbtHT9HEWXpfJ05WguM1gDndWrKirBLH0ph
kub3WlpK7g7EmPCo7lfnTR7AgIsTFPtL4NcikfJwk6/PMG3WUsInF3zPHJNhJRBYTxC26nk+Ln6S
mmQsM0HUmc5yJSPNYFaFZgFU9NlkIeIYZ5ldcCgJoIoUCW2yXI+J5colc9FR+IW0di5GPKUUlWzJ
WoRu2hkzsjjSFnOAS9y4uVKYfRTqwdYT7egiO2tqIVepQ+RfxgvNZBGqNqhUd99k8VKitKtj5HYE
/R0hDFooc9u2Xaze7NiNgxf+7jXdwPEJzd9NuF3YWx5Pfl4aqpPNy14sPnJGtL8kjKqNNjnnCFTl
oJojC23rSDQHFD1/fCI8H27prECKQOYwLatEvQQeh+pjlltyvz0YebncUPzZk6Jx9wjNTeRuGGGh
nqzc9veOKtN/vHGrBk7sCMAkF6/55WkJT7WYrvyXCB6Je/BY9q2fu55QcxjqYsLbRdBUyGEKvztJ
ECyQwVEXQJ321shsqEFjx0JL4CF2sdIIYaNDs0SoUTEzMS7arTfqY/ShMUmlwzkUr7Q2zn7GeCzF
YFxNj8QUA6BWL6cN8HRQRJkpZxs1OAaXJIBy+ZuXZoWUIk+UIGebT3Og9PIU+FTlInYqIsHndej1
S9E67+3W+ZG1oEMn12u4QatIXWPVKZc6Dry5xvadjQ5s19mTb0x4l6J+EMAUe1b/vn+YDyP+/Qz/
x89/ty8nOah50pc2yvoHmgooX7ZOE2BeLnKfwT8WwXz3y38r/wXTcQIKk6h8ZZ4zW4Kx67cgM0sq
a1+bV0nUtgeEyaspo+1nRtECaHOmR9Ce7HMiaDQQDduQ60+uxDz5jlswBo/CwHBhrpCfv2q2mg2w
95KgaKG/mrHDuhROh0KR6A+RaR4T4erZq1ZX1za/XMrADedpkgNuSEDqwh4vEP0sLQukSWJ1d9Sd
PCfRbElHkBuJRtnFDlSJjdoU0ZDoQvItNCje+6m86BNKVqFzMiaayLnFKUZ+lG0eyHJSiM2EwRYS
BvQZk6q7g09VhLKQ2cB8hiZAGXYeTUrqZJv3S77ZvDWamh1yeCwjA2spNm6ixL2K11uYLT6kcjQk
FJmygGHCelXcA5PAJKKuLkZysoY5kLbzYteHdlHERjmxNS7r3NN4laRHYefd2D3xlnoLbwfUFnW7
9DmX8pu6WeniLNtKBv709qg0Lwh+buBv/f1poq0RpPIxqjb1LSJmS30UT0c/L4F1gY6B7XNZFgdM
/29kzz2TrWD+4LzcbV+5vy2Us+VgvEOpVQnMSlPMVzmaA4uaDu4KrKWMbl5W4pOpcSREmjO1oDEp
DijZ7uA6O/9M11+brAyInAiQYbeMUn6k/187r8hfcErrMoTSqdSSn+AEVdiQnx2uwgqSyEaCqaWp
VfG2PeYukke7y4CCN0ngjGDK212Ks06fPaP0/gYlJB2DQ5j040HIVbfl28TcAJLvbn7f62puhRnC
blqxZ7tg/zvrHLBJZNfk+zAb5F4TuDyKTf8GLJQUvtymuO0BTqb16LUTYDCqbXANjAqjWdCrG/1t
hMMkKi8sQn101P0gAKcEcsqWEVm/q6+FGfx1ecrmNjDk2KNCe/VeeDAErIC49NCE+7lSWikmY/yx
3uvkLbRczCghTsZ+PxrV1OJCCEijIBlmvJ7WhnK4Tg+ZlidcYDu2DMCrTkJAYvJox1onl6Lpzgdw
rbF5FJ8MWdviwfmydb39AqyHygAdlZW7mdQ1++Wrb12WoRY3Gmfv3e52anpYWEuBzhpVXAcFEa5P
Y18lOfK8XeSjlaKoDh08qH1qVc2vkatSPCeDUxBkJrHjWsgVPrtQn7YgBZ89qPBzibrVPjfuQpJK
CQtb2YJG+9qiIbDIvcqfBdABqdwTclOlH/wwuG9shLlup+N7RFKdnOo9AHW8gsFBxwoTcHDDuxOn
01O4ODXGM1//OKDp8kwHl6dJDhPrrZLNZGk9LLyqwZdi1RE2Rgz9HX4OojLcEiVQsMagoRnfkoHf
LoFW/Bjw199pe9PGVlnZ5eWHaDtgNeMdhUS2wdrH4dwtG6liPtGil287Eum5RQcHFQZ5EYxY3NmZ
18YXFheykcmTAeJ12Ykn/l3P4hccgY1Tn4gWNDkz2T0P9cWg5dwuvlPGs+LflEqrVh+4/QujjKba
O6JeQAPMy5qJ114yPqg1buTSC5m4oRT6zQCO79K4OphTVm8CCsYEj2EtgjOXBqOKgiJ26znmIoSg
Fw2gtt8cX4VkxolgKUhea3WsgWgL69zGBeG9d+tEnRBr8Nn4gKLNzyRzURg8lQdo+E84CT0HgAYk
y07yGN5JDGEb4bmrkCeMedxjxiFxMWakjoKPFBpcKTLAyrCIq41uUX3J2vbZUO7jUwEjYloKBO6g
so9Q1DrKkdFYCjms/R6M+A2ceBjP6GQUTYrG+VCyta02J+J+M6r7QKQd7ZG90rjF9cICZv36tWJS
B+5mFwrQYnmN1prF7CAot6SIk2lzciRdwmmuSOyw54gfDmwKKBcqlBS8myn6fw4WAlTtw1tCbibu
L1HqvE3jECp1PuMyK3OREfIYSdODr/R1I0jA62f2hNI+FGDIwhQk8RdN0uJSFvCDNJ2edBhXioFT
gbtMQJszMV+Y3XgyRV9m+6P3ErnGqkImh3no85FycFZVAgOoBbqXQoeg/AHlJKNw2KtQCWjWHBDy
zr1k56RDzCU6/aX7tEUe0O9qI5f8NeStenGUrPo32o6vQuYJvINzCslkP3SgQAfVHBRvxvgpgUU5
5RXixAxC52XHa/ejbvIJzeOB+FVxAuRmVGEgcu2ij/wU2vUF3QKgdCocNuEI1VHu7d4cEKn7oaRn
jd3IVw00v2pL5ePxZ6griRFFP/3lBRQ53Z2PTC2z+JwRgmNJAMe/WGUVwTJerjR+8sY4YIGpHw++
tfhsJ1GMqZSO79OhUBbi7LSe72zEQDnnkloFXjay41z7INY1jYKovGTjGqk+ZxOQg6kCR7jmY9/I
yxkDWg1P5PJNgEmykMkvXET8oS4PVdH4PX1+lDATLUS5Pof+8LeGZwHpKKXJ1PQlMxcu0hATzrXG
VpStq2WtGHv4IAK1GtSvOxqq5yhGLXUmc9L3h38cvgB4rlGo8GcGFlMpmpLz2UwdpQ2Luz/pd0Re
LYpaO38zxZe6QSqYXpQQeN9tQKDVX3n/76q0SfJSt/ABKX78oF2qGYQb539GYP2Ws/LjQPtN0PCF
VCrY3EpY1xufqO0SJtfJ80WaYFNHmu9xwv8tk+JNprMEf7Od40bIioZ5eHsf3aE43LZN7FD9Bc3u
wNlP6sT7wg7HxlMTcLkf2680brmKrTV0E4pyRKIAPdYM0RZhSpvNApX9LUy4GpgAsw1NKoKgq8nJ
uQSDY8Z+aND/F/ERz18zisq4q9fFWdHLnaW6z7CAedZO7gd8onYJDYvA9ApmoXzJKlgMifPOHYom
H2qQ0amJ1U5bPtlCKzzLxlyc9P2zkf8OVTfihEyz4wT0dGTMd8GM6Ji/Cxbd5RlYbhEEe+fTflha
xO3n2eR/7ZM6b7eJwwfwAUoyfM0tpqzzCYXUhy83cOupU/0m31vYWJDNhKPrg58+DRrfNx77d7Me
z2V2fFRBrXAFdNEZqXxh8tLNbq7pgay1iMsO4diQfg79Fnk2uNDaoHEcTPWugLYlmKokfaDEhQ4t
Ac4dw1L8ACMgjkdv1jgYZtLk/Ux2w9yF0TxMcS8V+LtEiNO1IaPMBCbXWqa5A93yziEx50RXZSL8
13/kFzq7DBLN77OOYxfjLcIqeGAGcSSZiFGxf6+jM5ZprKSnZGijl8ZBuqdzZ7+AKrziiluP3oDe
NbkHIIgAbpwtvXnzdAUrhx3si2DKZz4IaHmmExchn06wzuiLU7L1SzAg+Lt19sbi6Iyr3l6VNntE
7tw9hPuQ/Q+vKNID5xYFCyJO0GAQDAMX3ZoBKk9lAjH8la2ef+/IDdW1bhV/8/jIuaewkwOSFkpS
WOWx/InVShXyIWKbklv0ESNnzJhaJ8LycvhW2jihgLHadNQH8gkBW7bQfgNylC9Mlqt8wVjkIHYz
mcLrDZXTp0wsE2LYMfn7kSsicRVvXKIqNOohiDlKQ7hzdsSy0A/O/H8hEYKZV1uG4PHwTnFpmqfY
R5/bn153ceMN/BY8xExEe50prjDi36dh4JAgeyMI3+isNlTWvXaeF7NhyrSgUxkD5ik7zkKtTIb8
9RW+o08q5ArlVw1I/NE3RoLNAtznVZOCPb1QVLjsaymSVZjNK8dgdYlwxqgt2w1y59SLfjGXME8d
8dmSUAZDXzP7AaeJp1/a34Vhgkl3K+qpy4NeOSBEv2wcCVwH/puV2pxqW3RukDWRs+SvoFPncF5u
Z/64zSvTYZBvt5xxAjkgR2Jd2y6oYll9l/ZZ/MXuVpOoBpdvIJbtlnSb2225DhZDhEWQD9GURFXa
BgAVJqg4Tezg6IMGXd4p/a9Z2o8IDplTgYD6oHxK/dSWU5zwrD9HzczfwWrwaj70b6FYPuoHRmZ/
DeW2oiyG3dygsOrPLDfDujfAvU7uzxX4tgraGvuOFx8e/shhA5PRVPXzdJxuYbYO9eCrWo3kS1n6
D0pN6R88n45Zex1coMHHmZv2JqdlNGWc83/aminiGgEQZeIxgIWGX1C7uAcxZgxo0BYVKfzmaz41
y7Z14axjp9CAJB2ZijY0Y3QO/ZHeXkjJwXvPosXtfG4439OYDkQtKJ1lGpQVeRWZQRSluhHsHmnO
ArgokptkXzCKcFpXgjedcY6/xI6mHIPnxHgNBZtupizpynBsTHB5xoAYDhsipMA1CPziQHFYJxJW
EmDoXB6H6jiiZdpfMtfCXCDROLtJgnVLrvW1Voyyp29O2hHw6IZG/+sOV2oa3OT34Vma4VO9sNYC
sSgbKmyfM2UM2W+b94BS1IsYbt9paKoqNHcQrliIxxjnRt2wUqQkh8pR9OZ0v419qwUh8D4k7NgF
pPnAuvqa1bGXmbrYyd9iyWzkMcRmuhyMvgrsTuWHQ6V06Ru1JUt3KAHgRtUhxDrr2HgTYLcuXjFM
AwbFFzrlPIUSeAZXglIiY0JsDzKalf79R8RL2W7TNnZfVxbKz7xSgqx1DsMHFroPVqHpVQkwPshU
+e9lmFJztWqjweCAZBts6twvVmeqDjWJAsGefptBIAS3FXqytoqDxvmgh8oLEyyvo4edW4vAwbg0
NbedPz4Biv7Gw4D+clC1C9q5aOHhgTDLPawZwOuqe6JJHyniXHaHwjvITGH4BWGM25G3JC/e/q8c
04vFdTgtTMWhbzgxWG2T3Ri5BPPfe8DB4hFllocXc+jC8OffQjnR7mf2T7wNZ4wMtID39zXcf7GN
pWOzTfV4pSW0yvloVYnlnJHIiVujiczYKQgNCL9uJ7wKXmERQftabKEYIUYPy5I2vTYZjSAax+WU
YeetCW0qvpIf5+Koe3m5L72C56hu0Btp6vu88PwOSgU7JNe40zjxfb+9ffwKgH22nxboxuWKklMb
Zob87VWZI9TSXwaKUzRYcx5cgHHKmdTaiLyt/hwZhI+hJTFKoqzP43RRo1ejjaNaJvc0dSlqTipL
dpBKxalVykse36CsSB++hfOiIYUZwTGf2BhaWjZQjXNGidxxXN7cNYvz5rmrhSTrzFdb2CUDMctf
GhUgT0rpM6LKuCMZGLoMT7Mui/noE6WqnXOnYFkpQUfT3Zt2lcDbjjfNkM7LjC3fX6UX8i2tqNss
m3UxQbBEJntp39kPnhEs9fZdjLmBnwEBtJ8HWXHd6b2+J1fTNqixHl+xHpDadja+YQOxWNrMddLg
d6e1qGQpyzT/XnokHa+BUCKNTsRjlfQl6MKBn7No80Ymdq9Fam0m0dWvsFWpNZvBIuwH35prKxIe
mDCFBjvpTIakeoe/nNTRmxAuTc8DhAKHWI5vL6IhDsfHwVLqg1hNIHAWZWsX9iGWU1YpTVIVrqz0
Lwz8nVWlgfKJtuO0TcsVEg3727vIrpHPZg/+70kMO8AR/yYR4cWNFzeLGvSyWLGmU92xPoTApPvd
iulgZCDHIqTDhGx/JhyR9klbQsr6Op3TL+vM51kYXo+VMI4QZejCzKUp41cg5KpPfXrpWkwS09mw
Fah+F8z8WcVqJFt+KvTUHTvRN/X28BDSHdpA2Ykvne6SZWK8DetaZdyBbAX0LZnHbjnIgNOX76i8
9il/u4+cT+i4bYPPQcSS9WTnt3ltQ+P9HfvwNGatA5Z6SAOovW1n7czUQQxGOfDHDzkaYe9BEMA/
UmL80Y3BVlkIgATAW2FV520iNxpvErSr7ow6Gf75YXjH6b1PdXmJBRcMDa06fhvmXxYwR+PTlT4/
lO/2IDskHZQcj6wMmnBpwPQTz6GDATU3fPrh1ufUNsid/Kf3aw5l23mZ6QfgR6k6mFlS0sgWyXCe
O1BThM/RAcEjbdDpygGK1RevgqcOV0lq7kZFXBhD2tLIZwXlgOgGc2nkKezjYqCBgOOpQotd2lXw
6kFH0tqxira/luh9eFV+xUMNJC4NjnyYufXkfNBCmvl4O5/YBoS1CVxOv/9YLGNW0wMyfrUz2R4m
5t3+GwZwUSx0vcxcfLyPRrgOZ/rgbQDhvDBA3u/OKqMyyIna6JxoLRR75oAr5nkvVe95wJiQJ+vZ
tOHZOl2vE9NKuivrcismF9gZGDRTv14sqcmkcnSywuioe0wpT6Qk1Ph6Z7c3k327JyXrfy/ACWIQ
G06a/xj9WqkHsYBpJsjaHGbJS0R3m5GET+/LA7+ll06ir8QtjTD9MBCQEGUh1LO5mOAmx6l6mkrU
5BJt0+Z2LJoACK3hUV4uMqdFLjy6k6YEbk5wEtLQTbX6X/3FBby2MH40WkbuwftKUZQNJsNnVdsQ
lm7djt2Bvcc1vqCls4OdalWYn/uQL+3gMNhmHvUucaGoF4e5yFPTxEwRGe/ogjssg2Z2PL0Kb+Pu
hmALTlJ8Hg1/eyOd/g8eKnw7cb2m3XrWHifngdP/gNvJ5X4pFnerv9tABgvaRoOi44lO6OKn0q6E
9ohahWa3lXjmgdxPkO+d/6C1oIt5yg3qusv07rW7jyLkMh/ZqQhCMcnjtBS/RSlfpPdT5U4M6LLm
AvTYuhdp5uFYETwa+nNIMq6QRbRU43eL9rXsR9JTmcpbegCTppbgXDubrjLQ+7JYrhR5aDLJKO5g
uyCRPeV44fiC6opkbhr+V1qJZq25XumJ67cxh2GAto78sIEkqepNMfnT3EeTI3KjX76LDYs/0U5k
9V5uYCZAUL2uAI1+6Kk5C13pdobuxH+Qx+rjb0Q5UrtHnEfQHjA3FqkemrITWBwZTVpH8JgMnOqq
r08fRI5wL37LN1ZQwd0FohkixjSmphmq8akKnT3zYGMEfGbn92/xT4o82rwYZZxefsEA+l2nztcc
HOcH7oKlNEiSKgfAl1z8O7hMjIgX016PyJQ8bTN20RXRmKwrj/AwsDUWIMYpxdKc19Oy89vhM3CT
0fPWNjoO/nOfuc+XRgxEcDdEbMrHQVQIhw7mhmboe29Wph1M06yDuwrEzWd+Wg7xFHJs5Q/yqytH
NvYgeeAAMIU0kARbZo/8tEtdVIOTH6gDBBB1FKnelMRMrOMpqDE0l0ol6GgsgwQlFYeS/h4gI2QM
teALerM6uU+5sBTZd2wXTZkyhJqW07bfxsX2tnRPE06BixAKaNO4hj53lEwoVNN9YCrVZ1DOIQG3
1dJF1mR41kB6k4sUX8xU6UcgN9F9SqxxMmDyMay7F8Z1Bo8+6WiOt5dvA2symOLVMQKVCNrSHGUk
58pO4xLiWp4yaJuww/OA0NxNpFbBZNyP0FrYB32/p1YDB4qJWqtS/5GjgZFFhl15ycjTMkyJCQVG
q2OHD1Z0kDDcWUOuIPqwOSzPiesohrk8XIqAlNoDwZe1tx2HPYelgGP8GzugjVq57GytPkdG1DsQ
OHjq0fep+cZt1uunyljhk9/ejMDXQ5XnJEyl3OU/B+mg4e0gAUUNkW++PS2Q6weCKT+SgTPiW8hp
chtaRMuIobITOnmlovwDHL3YfDoY6lU73SSRqNJUSBMbpcvwomSnPYCyJ5x/+3O8gUjJOavd7aeT
5rLz93YbY51GxpWaXmpD6cqZ3q7fplMRxTu8KXYy7UztIhaDnfoVlDGbeytNnRx2l8GIeRT6gBT1
kyr4kjDdpMnEgzU/KQ312sxWEOCyOi99/XVtPFR8wRBCuP/8wtxyZJ6Q3HZHGzZDZYIOVouCCdgB
eP0iQvsGR6vVVmElfszQ+K1meA3Qm1Le4A+MTQnEoiupkSH3KNQ9KPaE6k/TcjlnmWkm+XI2N4lZ
qK6s1N6igeAtOADwUA/zDFUyI0kkDqVQnFTtBMh/++uFPzgQ2jcDAue9HTnK4OvUIH8mR3qU5uQ8
DKlNaS+klG4YpYMzcl0taJKakZOCw6nrZWsXfoxXs/brfuaMvpct3Hhn3fPbJc7/dFQwqP45r65S
Sht5xdkJlSapTxPWB8uRWpQ3CtRFhK+9+XHMe7pt/M8Bc28Rcx+nznDszC8WuJi0NR9yUWyZ7wQp
8ilszU3Gr2pMxyL432fvVZ20Jw5Ll/UINhkOWZTdkf9TROUb1jasnD+nJrggayKXMPMZdGV5C6LT
Mwb9H90IImRTNr7oYl+AoX6Wvm9BVNBctvAwCSVr1Muc7TqIjyuk651xOt/qtMgIffXzadsHCvWo
jzFan6+gVgHS9tqPG666wOELMxNLoEfx2pzMvKIt5cQbUKMk1fwcYp4D0L45ro/JisJQVFpxPhG3
KuXNXLZCIg8mNgKrbcwl7u0Pmy/0QgV4wfcONwWEHfNeFkDAHVRXKzSAa5L7KzBcw4i77BTVuAXO
5GUQlSFiPr60T91m8G79+vOxqmaHCnehcy/zpmMX2/Aiqpno5B/sach1dw3pRoPIX+s+quAfPjzs
nu7iGrFgx8x0keGj5nm/QmO7PR7gVxDprGvCfeY2rg8iPz1113zpy3UXOGzWKm3/Jvk4w5UxCupP
Y0zMfjSnJOeVPxqpkBcBaveGRKq3j7gnrFeLGwl09V7fUOCRrUlsLffdFfR5Ehr0E3K/uLIQ0Kz6
CKoUqLuch6AgeysFWot4wgCd+dd72mSJgCyBDcflnfB3j/fJolCQEBklFJm9J9hy43kx63FeHle4
YTf1mt2OkFEMyIw3wUMqILXh4z0mvDz6vybc402yjiryBB//AHtnMDMdPHXMPUW/IyOubUb2bwIC
PB2woJKRsw10rDMRBBhwDHt6lUql5hmrlHR62clT/Gc/kTgOyZrb5O3JbynB7sHBsshuh6BDuBDp
ku3G1qzFjyC+Z37BzrkMQjqAhmxI9EdGqhphLP2AIUnLpxiX88Nv14uJz3mgXksZ2mwoeJNKvLB7
21G7ofxtcrPSjBNaqVRcIMAmhZOYwxLXm5Bzo1GiGW9Snt/HH1El9JkdR0o1jpo40K9B1MFuZqjH
1+8SPPSEs5abFOY6qQRMdjOBO0kVEIL3DZmZczIv+j/73S8YuV91Q16Kknu83otlJItbI9bPICzM
n9bAWTXE/npVZ3SiTGOgGovKQTXKzjhxXMgucZaNs2SgcV9A/pWu9DUZ+JSs4+7jwe66aRCNFaA3
hePNlWgIonFpBWvPsfHwmCwV/C1Zza09Cns2iJIcLlANsMTLQoTtDV63aiKARYLHRNrBJLTQC/U2
30I69bgxJD4HA732/mq58kGDLCAkm1KR4D36gqAc2ba8nGZR+ARFPZ7D7O06qOUIYk0eVVfyiDLt
aWsyB6czOd9e9aNOglx7ktyeO8zHbKP8aT8NAEfwkG+6HS+Ko492YZOWN27X2MhwKuHib1PG/SOK
AA0fxIzSmh9ic7W0QJMEzyVtRTHUfZ+jX61zUN8aOaDTPg4fTS6pNiHAnEdIaBQJ8UubH44lMc65
UW35N58fYg+wVTZspaH0PoxzuVuhRQaOBtQwn43TSax5fWpS3Y+dpXUDITJ6yASyunuDUWTQu+jN
AEV2HBU8uvS9z1zUzymQWJeVpolLPYfcYDQjLcDNJCeFYi+7OWHgd0Wf0xPKj9B3an8wCh2HKgot
eOmtTSS02zqSRDX8O/Eb13bl5AkwTUTelqHr1zbfXVX39qQRMPeZXP6MaV7Qu7jMNcDSWy2x2tXt
fZc9+QuqSuIIYQc91q90aRmPgyMiXDfB5trlpm7umeZsTG+tAyp1tW9k9Sga2/XBGgWUd+0XAPOO
2rflsZm27bxFivJSWgR5g2eiTgIUNMfeQvivg0j+F3wSkQZRnkZORyw9WO4Hitym3XR/GM3Y6jgt
R3L3WsHbwXoRjdbF0KrOHXXxXT/UCIGkpDymhuJB7l1XAQtyMECrNqkyDNeKd3QJH5wkPaiI/Vpx
AeX1g8OGIx0ET+5Oywxzs6LNFTG5GWbUJDiP89ur9zYCqFYM/PnXFeKiCoGE6cvUMjiCjcp/A6ON
2lea+3WGvwHBM7pBSiRZzsnO0XxiPEte0n2LGUkWftwgHmJ54GmwcWZ9bhpquQB41BAyO+ovpDnT
mwRr9HEv1Gs1Y18vwoq74BB4PeZISxKEcE7PSUCKbsQgUKHHnHqRRyC8aHWbG9J430NSpIZxe1O+
cY6DtJ7mCgZ3zkJl9CtLMHEDJddZCzioGWdQznEUhZVXmb7YwXIG1rqOwaNdkVIu8T6Xd6eW6jz3
a2MgLb3V6F18gVhz4AS6FukFatxWXRA9Ikll1UR9jXEsYUZy5pdGA2eT261VSMyJo9mxQK6HgWzW
N3tsfg5s4ZfHIq9E0cdFw48ENtwtzJGAb8Fd48D3jQjZin2QaEFJIbFZjHpjNM1kROcZp9sEu5dJ
hM3mZix2Yvx9cXOQCS9p/Y5l7y8imA/NIMrWoZnVSIzJhicnuLRvZ1x77+aRIY86A1YUPtpeYpSp
YVg+Etr7mZ2GPQkqEq5REaSSyi4ZNO2DDaAyzi/RT3kdz/KeF54oRRSJRaAGvsNd9vWSmiI1Plkl
rsCRezhGbkBYowuFd+xG0ftpSZyMQL7RenpsN0vLkOughWCtNO142P3R/dpxuq4gNr0oHtmIgOaJ
I+evlXKPd6u6Sn0Oo17/LP0X7Yscf1nS6LtmND1f2FdLX0Xh3gjhcpLwsti59N/Z6j2t6lpHi6sk
G8OEyuCIRGz579qd8xmb4iNH2sWtht2T9ewG+tV3tBZD8v5CbtHj/tZDPIDqsWsxi8GEpx6wnql3
A4b/fH+oV0+S8XyFjHlX4kbQ/hWqG/1h9Djr9M3iWkq6TgESJW2F3yLKZzghV8hH5TzX5Or8ylGm
BXx264K/X6rgjAAS8FecK6ZkbaQnLJn1a1Ar/9opM/iskfHJVoU4rRlJMgIi+h25DaNYwQuVOI/n
x9DSkCs7iO9oTdHipqDsftza9LqK9/ysHTpsNDBQ4Wg4XQxtDWISWPvtq16hpa3/Tjcuz4JVozzy
X+HdC4nH7wOuFwkkYGH74AcGI3CJ2ja+uLcDGNTyja7Ug2pnGDgP/K6aFbkYZrnDZGVseOWPgy/e
w7o2tlXvJlVzJxcPQOTU/poU9KNLuf9UFkd+sWhKA5tXXP1MFdX6JgfuRJbvJNlUizKHFUYKgUWQ
DgxmmX0CtWWqgDYCP8N/23wsssH8JndnMUNelJi/IE7344RVeWK2Y6rT6aS78MWY4moJV0Bn+5oI
grDncTDODfNw8hSLmwLGgReRHvPVTWpojWJs9ZgtRDVOy8/7PjbLD2grnBWbYyZgB0p5Syb8DbIE
NnhbqKdsfikIOcBiwaTcLedc7Ose03HtqqMlSUbtBZGEgcaqtLiX34tyR7N2rAREz6INivMEU49F
WHbRUqq1E0UQzH3JhfWoTuKY5YwUGKJPkBNrgjp3/cfjYEaSijr1cE3uS+TF4n0ohSLYvp3wpty5
5sMy4wTv9Zl2qtZccZX/SSgfzuLbKGmh7J/Cdt8KRCxyaKu+WK56ehxMfevPgcOrWGbz4G9rOZDp
PXHeMzcLvFpIqn03ThE88HBuLvu7N0dQYEnJaVvlqChtctINqpsBXB8hVdCuDepA60LtdElp6hpt
bvzJUc2z5N8zvjbfcf5gfqxPd9GSWPCwNvSg5RigD/ttbPkvTpDHuwoAKJAGb2IcbqQ9EIFJoIn+
vFY9wbJueQ3tamPIw7KUoiNjbkIVaKwmfjAwFSY3PoJJdWwA8T9tWL9MFqDwrvt4sDesXW20TRXu
93TMlI025CtYBqLdMo812PdeBz74N+iNEK3F//sy+oE930MKNZs5+sm74cY+pz0VitkrR+1WkpSf
vq7XC0afng/qz5QVtOFDxZjlGSPbfnGzyRmmg8wMJ+1zVOlA4LIdCTbVfJg+yzkXUWVoaTLw71a5
gasogpNrdSurV/kSURrK0w38OPG/vWHY2XPUb8Nnh6Op3ycn7XCoEc9IFdR0qzyZ9KNsEPV+w+JI
cATjWQma8wB2hBbuEzS+dpi6T/aZvFwDb30UHCSC2ZyZCaz1HyGBa0JvAyTcKWuEsJAjDfm0PB9d
Hl+ThOFvl34Phug7NVIWuHiR0pbeOrfxCshM93ymXVdry/ysJ3zAU8vSqc/nO1/+51nMOahSK8Uo
5T/WaG2ZjBEcfRcX78fLHwgPT6dTSpAb0i6HeP4hXPWPKvK+XdK+cMkj0upIih2ceNnEiwpxuxpQ
+D2zq9LlVR9BY0NhGYKoSOWal2exD0tPyMTWWdJlY0pTJkSMbyAEokzDwokbn4NhsOX10y0Uqbx/
kiIJdGvZSR9EB7t/mpmVmqPyCQS9xoJ/Wqyh+Vak3+jXAkStri315s6CmFmpNnFkVVt2s4mPv26v
unr7Okt2QPERoR3WwA19ScHJ4ZO+QgCQy38rGK3tTEFo0kpSSmR36Ki6ooGLWBd1nYhb+u040ivt
p4YraOut9AT15/Q65Dk0JrxEP2NEPatdm2nB4foO6REIpUcvYjWOCZxpIKpIJbbFDI7PqdgJOcvd
K+5jNb2fAlQfAW1nFhP8jP9THutZGCNW0GZmD7Omy7/PlU+D3FnYu8sO8nkFgB/qaOmZwHLheY5j
3DWNoHbdjSy6wbCB49/TwQgbN6D5m64BcGk4CVmvtTJ/PTc3NobSO2mGho76/XWFCu9PB5boJyS/
D/egpX7O6KL5VT8QCNFJdwhvkA0zUBSAZPwBwvu1AmryP46sb3FodMy0RcBEiI7BrO7oCdf0eH5f
lp0M7orWnxmSpY8g+3Ucuxh5XIZ1jFKTMAG1C41XnaxjC0g+/93GucaNaRoy4k5dVZ5LLaBWzx4F
u+jLSJyOGy1WbEHytxsbEjTWzoST9ZkJoQO2aqygLrYLCHjHw+FaFgxCI6FxIbE9csmRV8GeJLmm
lBgXmYp/+aSqGmlO6HZfX0x+lVXe358+Nk5Ceoax/TogYqE8Gzwzmq6LTJ//ZkFOaxhi+PSSBr/R
TFSxy1Aib7VN+y/ZoU50XCTIk1temhqu9qPDf9pqFTVD3mRQgWYKr0l9+auNYYvEEkxzf5kuVB0h
bb7x76Nd9Hta3HAME8n+Cm/Fw/UZsCoEB/OKIfseh4Hxn3KBMMRlkcajWAHpSOKa5kmsw5ZAwrf8
z+9NamdCIQDv/7PziSl9BE5BinoPZ+BF2m1v6/M093kHyG0SYg/4oNUj81NBhe4W34tt9poFwvCk
Z8glO86umkq0pm/7fTaRIchVXDf7Z01xNLu+niBno02g6J4AIXPYa/3HVKPG+gq6CQwJorikaSRe
J6aOEp8Am3i6BIJWrBW7Mr2tHtNihpXidCr50NSYjanNQyh064RPKOOSwCxzoMxPnf8vVjTzp1xW
v9/65Se1dBVKzXa/cjDliuarnLcuPWte3EYH6VI1NmhT+SVj2K31yQlvVmQ/IG7wDuR41GHb3zlO
uOeEh2o7OM7c3dZMjQ1ruffIggoy/VOMMwjMF9MzVubMhBZOJ6a8ot1nQC+U5va7Gyo+PSEslkov
64dam5yARjkLxavgr2l6cv6HjjL+HGYedpBWALgOTCJxDzmhAl6FcYt8/G2ywcH2xHqBPudkYq3L
jl4pa09UKXkWKGzv3WThImb/cI8Am7iDp7DPhzkmS0VN54Swvh9ZesJ0npAONBoTHZUbkOqhJ+My
ezfuxRu3IE8wnN3RlSynV/zEsGBguwoob2JAevQ0hptPK3tWMpxNwgsYzed5WfpkAsNKcmvhIiBo
i9Ok9IfjBO/Y/jKL8iPjFWtTAA5eAHoJ9KdJals4c/b2JU3FqElUbjPEe7y6KNYjx9CaZRoZBr9L
yG2TQ+NYy4FNkSpndLdsztJDs3fIxpeop9a48sh3v6DJ9SNh2lyv6/G+FvKrzGs9zOcDLSVf4+4A
17mhX7loglMSXO+OYyjDYR6egaBQzjHghzK/fSHztJFePvQWCmwIiVD1dqnhasD6ca8O8lW0+N9r
xRtg0vSlKxC0+5r+WMrlKpkOwaJ4Uykz3eo/m9+lv7wHdrBL7Z90YoFH3cr94v2OPZ+dJnuwPp0h
A5kdktz+bFL7EGUnk5xXkvH9AKMB9xGCUWSGcVM6caNEtLa7HuCxPj7xvG5e5DpX3JPAOQqE0F/i
4Pu1Bsgn1sB06ek5VLeBjJVrWOVg9wfb96A7k31T+Y5+/1NYyAyxy8vN2ycqooMzeNb3263544yJ
N9l+cskS77VRisEGHIpvI6oC/RRLbGH3ElWXiucD6E5LsjSD1p8TG9spjyNsXgdOP1HRUpnA56CE
q6s7bO/30Uh9naFWGDdpDbJaWFfmkf3Mqjs4CyrNh7rdw8sclK+zf3xnVzKBERqw6GCtL7oWMezH
jxbkjU8ka5BdBHa85CxAcF7tmV/OQtmCJPxrfEPVOlqVUuDqOzVz4Wwr8xZTqG9vZfjn3mDme9Mo
pTzavmG3mAEJwf0nfEBsSG3UO+hR97h8GVmosYewQ2RewYiNu+WOabo2cYotRojMbkinY+ubPU/O
Q7Awscf3yLBl465Cn2HG4HLPkmEABWzRQgsabZL9gzTtLirEWqZ4pjWHhToGt0jWaw18nyjQJP7f
JWJzhH/CIxXrIn428Pf/RVTeqjjZGCiU8t2HKevrM2NrmiLrt1m3d4hMykhGnLFip535XbI9Ue1G
sIyWo41WhySMYk2qBqKZidupSzXFNKGbIhEHKZ+vT+eAad2qI8QgufXgSotICs/xb0g7lUK3MYU2
YfOgPkQogdzQ57zJY9J1SWEt6fsKo4UBUSL0zn4nnWVGROmvLuoQMs1+/hd235vr9nm6wJVSZQC6
b3+GZW07XLBWOsE9vNTttGju3GskcnXnkZWWyVG9gcsM8zLgSa186pTJsovswdzXHlWVfQxCKMX/
6ZcX82d85VQswtrzcU53ttIuF3uoL3dHXOQdRaxnULxVOzgWwJJBnYKYp/wqtSeJpDkyqJ/wylFo
6t8PWLOxdOyN9zlwSaE2R13uQg2MFXDA66DvySZBFpp5X/8OxmvVkhY/r8uhIVg5uTRjRO4I+rJb
+41/hCmMcKYNteJY8tC2BGX1YxvhKz1EAzOyDvb5Kcm/We0lkJGuT4R/pTQc1Ct9xI2qgaE6pe9I
JwKDTh+7cVYwU1izrsPH7yvoEnqgXQ7hlkRyhjOE79rWOF1EPLdB3bqBiiz2CSYd3vbN/RvT/rBz
UfjrEXKKLvS7wyZdT7Zm8vQ3uGH0wAk7WAIv4fVz4hj6JA+p7v1V370t3UEh+Difepzv3iBLt0xr
io9+BXn31qnw8nG1W4WlM9JXSG6QXA9FGvrgotbxk6RI4NV9xQK9QHmJs3rR8abCXGn2m94Rzb2y
OqE7327QNt5EDPsC3kcaZYyualDUpWt6uQ9n2HfSoSkcYffuGzlx7CsY/pntEoDeWB/Hcokqrmcm
MF4dYThojGTR688qVRNceRtXILwZij7XHiSr+9biZAErgSqpcpgwjiyJNUWOxs5fc+av2vId/Szc
FynLWv3yBjXIaVeWw23hAkokJ47xaiGlXe09xnTsFqzutJFLCvgPv4ypwV4175N4eb/t4WjG+jPg
9G6CDFMJobmljZyigZE8/a5EXvPSIPCr72Co1JI6Y1r8GbOLtkILu01fqBN1yynJ5wXiPpnW8Vi7
tycTkHsAz/oZxH7usDMs1c/3fw+bUm8a3V7kvbg+HdGhgvNk9S8qADFCBwZPMK4qoM9KclF+OEpI
bZ+w8eA+zvN0ZYrCXbQSJXSBLXR7MiyYqA/uZztuAH5OntGCpxVIjPNIDvr2VsezkhHn+sHWvBBD
fc74QmvIc18iCsNv/XmJqgun3csVHgcIiWhi7kg6RIERLUqfvfGidm2UbuEhUav63quRIr6gow4N
nhZ87Ur0Iliw1GvMm0uamuFQRC1+QhIV2hAzruxxA8FT8kvqBzkMziM64EAp9li+QpY1mrpVQzvr
i4vHcSeoWqacJgpy9paFjt7QQ9tSf8jXILK3uLgKxgbXlhpSkpMP1DyLfXGy3355RxvSkl2uybsX
TWGV+aGCWenj3b2Z3E0NSsiDHGztiXXTwwNWhaRtTYBmvXVTlaIdF2H7FdzWGiEVPDNOPRSMXDjr
oUsqMxEEOYESfujyVPB6eKhqfVLRqboDeyQZ+y94DuSOX8fRQzJVcI/qPyXAbfWa1Wsy5j36QGi2
P8mzN1xhg0WHfUiVT0qHcq0lTtQuYrlhWTraVfV+BXJq3C3l7mETmn2qkYFFIF98jQ9q58Dr2140
yhV7NQfNaJ+3mWaDllrMYW80WFWr6dMGYw+0bVXBCi+RLD7mHdOi7FUJMlxYWFX2tarrALNz1Hyj
jOzpcu3NeRkqfmboTFTVZ/ryMUrYCzcWJ+OOagtHu29rdEsQXVgKbXOqaY+ob6n4cy7CifBm1kCc
Y6/uexmQNHJif6q1MYs5MvCvZBtXqxsFi/9N30VYGKZg5tw9OKaK/5R7q6mkw6mA6OdYC1i8bjuy
u9FKjmbgAs+wliItSiTHXhODQiLQWnI7G4mo56iqLid7UyanQBE02dSa6hizP24X2QL0v+GGJGkF
yUg6Niz6lRe/O7oAyqHnKVrat96WzwzXTDVztB6DCM97BlsBDksJ/pb9htYuah8cFkZ0/NaKTLdm
ekpTBHbvUGWrCgibjcT08N2cQOFgwYniybdY0xbRHxcpzcGpwQvTKiHOHTC5P3MPpcBj969QvR7m
1M3mEvGy0XRIwNvN87R1NcZYiHamU+lh6QqO9NgxvAWUzjxe4Gl1W/DgJMGQ0nR+oJaXZOBJkYbA
3iRc9e6NQGmoJyleLEaLUOqZEJQmMU2OMhf488Lssq/zAFBETXmnbXtCnWBcWz7IqqZ9pwBxz/6K
Eik7OPvuKcqWGxQvycDhxizaCbCdMp5Ga+ZVjkF1eD6uqN2i0Sl18qnLK0COWmtY2UdUsAj45p9k
UTw0uKNrlzfTfrsEVPN3n+plYUgGvAdfw8n99cXogWCXrkqwXfJhgYKrAjV1JZWaK+IZdvq0zf0j
I7TiVa7CmJ29o3AT8pOPuTSCUXSGFO1M4tq2u3sWUZpmZPoNbE0toN8Y1A3h7KHzbK/6YnlK9EWV
U0C17g10egFEgjxGhBuQia1qUo3jE8Reh3f6p0+a4iVFFafwUYUD9QOwS/W9a/0w/NxRJr2Xnf1L
8jBNo/488zXD4JjgOKcOObD5+BYOlc1Zj3xwV1EwXbvfCi6VHuHrBcQzIMZvljK9v5M1ltn1gYwU
zhXnkoToBkPXVoRCxr3E6wyoD2QpeGH22rhRaADpwLPoh6SBZ2IEFHItTW3rRFMN8YP1V90YS+Ms
ledrFYvP4bpWmwK5qjOM5OXdEKDmlZDnJT1usm2xcdejb7RGtImPsSXcViRllwTWB47Txttgp+Y8
/XRMn1MPWr3R+eSpZEVlo1qtGlYrtiwgKcOC29HaEoCIN93dKOL7T3/IfPYKXIK0dtYGND/URhvL
Az7Oz1+PSu3+/f7b7l5bZJQZoK+ipxhBocoCQEWNxGhdr5JtsUa2eu2fWiZfILSZReTlMv7NpU8y
mn5SjJt9YfkrFwL6O4gCQaT4yOGmDx0/yDI595/4TgiUN7NO3UOH8N0XQXLM25+PAim2XRKw2dQd
6ANeXTRwIF8NWw88ie8T2fuZVvQoegKM9Uzw6m/Z1nsEToBSWmF+dDjUHzq3YMbQolr7WXq3M2Qz
4jCbbOmjIEOdQOqDCObkO1nyj90zen9fnXrnSX0vUzD3f8OcB/xXdiAjBppzf1CeZG+Jxn3ueg4H
Mp4c801gcY2FfOz9Ee2HmpuXXd09bTVcXIZOYute9f2tMSAZ1gD5icwIZhl7tjIj37eeKkfnKhsr
ee9r+xSdfqknTN4ff7yCP/GVvF2WGwEhYmMFHRpQkLOdoP7P6qE2h3nH47cmxBjtDNy3l6gJWdYZ
qywc557Nkwmvdvl4PFmyMm9Dw8rvCoHqC8DdCI/x/JxVR+xqdWXB1QjaJIy/EUG7+57+TD5B2j8X
4ONw25B8u4ncTrdwUQxoN6BE3LY0sk+EBpVn48ToTRqLFgYDieM8yAsE5/oubjYBnoK2jA3P17h5
5riZj3Xp5uJzwBn2wVK+fWTA2w8iboSaxYm9A8euYIRfabv/hm+uQ+G62F6jHcDSdCtZY88Z6xJ7
ayhqLa6yvHTDPPHziVSCrEOEnAFnQIXrfNsE5U+shjmyFLftmi3f2odfM5yqc4KiqflBBHrlpsID
BVZ532Qu6zic2qsokJwaQZYawS8bHXxlqcD/5qWHlLNSFxDaWfS1s2etZcIppHEy4z0aZHI1G47R
BHP9jlPfj/KfhSZTkJihS/klFO/zsYU0x+boMC63d/JZDnvAe6Kfm7fWemK632K45MdWlNQI/evd
ADE65gYAhnJQsxJeKtF8T8XTpnQoLFrnAr7+/+Le2IIJHhvhynVuHcsNuUl5JiQ7c5Wv0lKtKwb8
TyXVmieJl71ieHBu6Yb57yj+3uQSKRgOvE/YFeDaBJIaHBtG0facLpDjM3EiE5Zn1P/feXBFEVwk
pOCQkxFkg4leNTwSP2TqHN3/VLh04VInVRaz11P+fvt39f0EgCD+ih39pQTHiNMM/eWyJKR5oYH5
g7aXaANoTSEgDuLfaG8ri4+f74tZ+EPMWzu3ddh5p/Q2lsafCem2inzL9z5m3b+QdfU6/O2+ano9
c/lHThK98ZSDGka9TE+quq/08hvERu28iGn8E10A+UsLaqleM/uomi38QXARcXU1Gi+Q24pGUlpl
lylA/CF18ObeWNpsr/tjwOC44TxazYo3XjV2u2sQB1qJJie8B4PzU6uXi9OtWZWP+gYquJfVCF06
ETPH8EZPK66Ov8sxRpFqxe7rNN/2BHMnz4khnqve74DQ5MxtvWCEW2EkUa/KY6UPwLtp8/ECUQ5E
n6txtvGZ9RnZz2hOFFWuTxQ4Z4kvljcDM7wxgKfeROTT7cJnImg5OyHvUcm1XWTI13d4XIWWGQjC
bzDNKalIjGVvf3ySQdUudgUCyEo0F1a1l0Y2OHYHE8OBSWCC1vdzEzd9Vt29JFD2wNPh7t1yRNkH
jzmrUG6/rsNbeaIr3kqPKeWzSRf6ZYSRZtkHudfKnLLC1+ya9DrpnOzJaMbX7In/akaBbT2sTHOD
hK0NY/Yc9JjrgNrQCqt5TBajnNGvcqCcKo/F8Zx4+9CPpqZkl2fdMld2uBoe8iliAU1hwnvwFRnG
kjojM02PCzO2UFqdHq1hYiFcJUISS69uZeWf38iCih2OuJon/wLpiVWjZKwWqTDiAwh053h+3mup
7LWdZCWx1smmHXdEkXabo8XOd9NJ5RuVmwZJylVAa0J2kOjbd+SBKWaHT/qne8M4aiC4xEcM8ir0
pMf0Li1TNBzqao0JT8jYtD9uR/Nrer4rNK6xsSOumNj/+UFCG40Fpo7mBQ3Aw861ebAaVa3Psv8t
mA35i2696e8yZjWK+je3gbNHSzr+Z7ZOZ2lC4MRtNrxH40pprF3C4gSxKbFz+fClivKdEFWVpGEc
GOhXf4lMmO8PYrOwrw9rKeu9r4K6SHMPRl4/Mk8ERmTPgKLWc0b2JlyFiPc451YP2+ez34yj/0ou
NArm+PcsW6n8ywF4cmtgyk7hAFduOXs1RMrp5N3/Zc1qFV/q5GWLWgqylPfqERdpVv28/9yvFpEb
QR025EKmKa9djZUUc73LISaOqp+LobszgwfkCsp+xDIhatWgZ51BWKgL2+xwL8hnbnEVNYITZV3t
k+1hrE7bRE16TlOLcY4AgJZNX1a+Um9hDf2ezvz60pZbbgsjDusU+bfW4Ukdgfse6r00JqMITFyu
XGGoq45LQyMdWuT8iOP5P7CyrIR89P2K2gvEy1FaKLCC8RMaIXuYKWzzQRg+1+Uc/P1IP42UiqvD
aJ+Da5+i6ju/S8GLc77x3TzyeusBrtKh4Y5TwblROy3sp7fmsKp7fA/337jeg7IWt60c2h813q+e
AbSUhxIW9fynERbcZXWJ9ANXvNJslYp1faMTT9iwY7pT14FlZTR3S32AIp2/v1adE/P5/Et5u9un
XMUnz/4qOtb0S4Hh4oXZLbMdfbjxznPbT33qzvRn3HD43ctAMK9LRoTrjuF2tJXpFaeH3SyVA7nN
1g1MuPbNXWD1s3BpjlOTELO4YChm3SUpVPxi/oL+MC2vKZb+i1eXbsPlGTSqFj2Y4XW0D6GvVg3p
fvYlBlzAuiE+NzN6JJhS5XeOib3UmSAOlc0/zp5xVSdHiaX6GY5DbRxf0idiIUnIx7wG9y3UV1kd
J8Kye9eIaHR3m5h0Vw2QWxcIW4fnqS/f7VAgdyYH2TIk1wboOMXtSx9JdOTo9Pu62tsFwb9dZFS0
5JU30lUpCGKrYI1mJfXq9Ux3LT0vOcNVVrah9kC6sXqB+UVT8dgmqTLZYyXUmSlcQPdpAEc1pEUN
gANmv5GhNA6ACZjD+NZedOhjaRyrzaR8E+EMSHFIuRqSOo9fAepMn7yN32vJFJR8wjzfqrXDxFOk
7pYLXP2hj1B14jtfWGIc6hrcjki39cjlt4xClMvmh+gCUKoHi/Jp9EAAmseEZFkKKae+UXSaSmnf
4q1XFQHUImbddOPDOyuDqHfzXcpHsMHqNdO9TEuQTFgYiP9yDgdYXf1crGZaQRCiQWzQmXzg0412
jWUOwBdI0Sot6A1lcdnrQ+bbLf39njUGJIBDW2oYWsPxp8BmSiyzkddeIjIXiROh7jLjZ4P4GhQs
ChXuoQ4pMtUP/4ftx42JBJ7e9EHO9Gi7jnkr8rXz6y7lKd11IWAMKsLH6gIXxmjJ+p/vJITAO7Ny
mcsWUwJpwFQYwIHPnPzhLYB8fqBSeuRvI8tIsyqVk1jydxxVtHGObgwAXZiy2o4ny3XmbVPn+l8M
RtEvNUpG1fie7WXX+C89Jns55G4btE3ndIuSStZQMVYPJoRqpKBd08N/0Z1dpReWHshO068KIWIA
3pwCDseOpqelrJylVDvnb129uXO38XEhUQSu8HTqcwa7EjjWzVvfldEplKAwtuQ0qjXadVh7v7Ea
OITefQ6MG6GNyLCxngNBU1PFL4Iw7VKKS+MNGsifbWip05Obcfs+UuZoP5URCstNjfv/g2dQfCr2
ih5qlqIvXc3x0y9+SFX897anq5JbRmaIqdQRV1EZHCae9KxkXMlQAYCmAYKL8QbnpR7PRIOorVlS
d/BZc1u366iabAFgw9j6a7+K/FInd/FPUMQz8Ci+ULUwjOFxV7xjMJDzApWHDuZCgx/UghKgBE1p
JuauhD7a3qUFIAnjBT9OB9lIM/o2n9U+J/6o1ardILbP9TWiUCyhcg1GTYWnLFeqxn5HEr9uFI5X
DwkfD1IF1b6fhTBnYFJagWL9BbSdO72G5OcItMrx9iGBfudRlHBqiBbVzTY5i2S0WRC2sPy/GIks
Nz41uOs6oGi0cFr2Nl2pCbpmPLXAXC3Pjy2j0X+3YntjUIQULtgY4Soc23wOiMgbzZgWxUlHscPb
IV7QByXmaPAgCb5OfEhN6CzhW6Hqinx1uF5ipfWBiwptSLxRoC+QgdKGQyGPNj5K3XjnmtrJoHqd
90iL2kzExmJorlyq/yp/i5Oh+jwFnirNT/OEkfnvCooU0PDTVWvlXwGeH7M5JrvIIvJKxVcqUdJz
3Lr6QKyd0JnFB6Ohkh1HuMje4z8iNy3Xft9gPqsUdU+q60N7m4ifazQfDCFtnVb+oBYFM042gGVY
Y3uVJbQVkiYUsCXC4/JkouyQ0m9RJmMt4mj3nVZGEHUN4qH+gd345+TroWWTvO2/tKeBHCcKw2Hd
SyeSiSJJH9PAF7A2h4VF5pCNfBTPqiIw+43TQMN7/W4GmuDyr9dYr/rq7Z9QOAfXOIJWdGmlCPdx
3JLR3QKQ/FeUBXQJL3SnAXulrrtD3gnOna3TKewhqBBLQ2ut+pQLboDEz4dsLITtSTJgicyDmMrW
J/eOExIFwXCjZmvWLx9WF4UJNwRrfb2LKmAxjUQQBNDunKRki71RNZWDdvb3DqGuIGzEU40H/Lr1
toogKIqCx2a5WPh7APaz1Fcqk3eLT3qq5Xz26HUcuux7/W9xq68efFGKbYDRzLhSdmqJ2Vy28M5/
UGIgN9MTvvjnEiE+6u0MRv3Ywph67Lr9DCvkgEwH5JNfq6Vc9zvYRIwhRBZE/vgV/0eYiAsiDYor
P9HPhnKPDk91BYPP5qv3NF87YXVGEzxVhGx9GfBeNigWIcItkHnCrA0YNTnu7kcZdN0FK4K+sMUc
BdOJ0hEBv5rTnorycn96NcOaOloiw5XrPT+vTuAcT/rQFy7dfZbHmxcJo9PiozchQONoG2ZRcQwi
IVCZCVQ3vmwwf08Yer0+tHZSqlFvzLg3Hx/5NWxN+9lUcmcc8knl+DOgtBgUCAX0zl97KyuP10Uh
IlfHFIeHGgbw2hjy4EMBESF1kYkFrTIyjtFlY7N7xrcrh2XK5V7TxZQ+eBy70RVMQPekC+zi7VOB
FrQtuoH6nL6CvZLX7YgRi8SrGTv5r0S1JV5YGbbH6mzfVk4lrnHfyVRSUudy5PFMknIfHM8moX9A
6y0cli7qPlqs13PZRUzqNSCbI2+F4UI5yAi/yqpD8jAxp29Yh9ALkdkD3oMy8g2L0NECBawF0F8m
iOxyPXQptxbs09ujT5TtS9FC7AfcQuzuwKxKoKNuTe3AgS/J3PeiVR1b7MzG+EQRrnuJ+4U1Mxxr
vI6JtvonvY9+0SXLHzwG1POGa1+UGFFvSVaIhbT4cv7WIbkuY4gXYUN8LWo0XeN/K41ioneSomhQ
SfOWp4GN559QMdalmGrYLCK4tKq4YccQg4b1NtArOZaDdZmS/CZrJU8gU8y7+o/2HMazNRM/r+Vi
+0YAXz9Cz7nWJYE51C6MAsDGDSte8HAeN5nJPH9t5eijXGoZv/U6ElFaYqrNlui220koyTuNFqUr
a1ZYa2lJyXbnv8To24QN8H6SAB25tA6u5E/NQIlcQy2FZBMvvuLniloAj8BoCRk117XYrnMAS9Fx
pL7EO17ZyIjrx9FMSuqzqupxb6BKQhdRBMR8dwLpGk8SZABLG1x/j/T4ijO1UDq7Hbvi2rvVE5+Q
80mmKjAb7jz24M4RhAszk9aHqAa6CWT/UERW2UjakdfT1VW5rELG+/lttE5pkZLqA1Ekbr4F4y/J
AI4RUS6CesQ14iWDR9XQhyMVA/ggghExSH6U9qPA2MoBfVI0a70/Ql7KU86G/uebo9ABQY2NEw0n
atRhYahVLkhjNWo7nlKNTTEeSicG8yTvmOkcD+FyQXu6nD6v0t4Znev3Y4OjXYUJ7xZwDd72qWEg
VXHQOp2decvYKjhYV7PmHs6fzhHe9rsuONqn4HCPMhMnfXfJ4oVSioOXbvhBKBs5P4U3BFeyhW8+
g5vyzKsTHZzWxisKo18y2ZWpszN9dJk992hXhR/VBezvNRO3G5niiooKSDXphBmInPFRfAvLzWe5
1evlq3WRQrgjun/rZUv1eusDIRfJJ9xyHr+sJK8eyfGeT6rgI/CmA3L7gZBJbZ3FDEQQIhzBAA5t
DqGW+FtGV92+rOMA9TsiuMaFUzqit9pJHfVB1AJxKDrBGDk+zLNJmDEz0MTMaBLtO2NchBOQ6tEu
Ay6BVdxW/L+BLOLIMUnr4ikx3ZNm6PAImFXIK3xjwAw7Q7qn6WVpL4kxbmwt5GNHFd2CHa9bpWNW
Hkjl9N7uGMP6PCi1SOtaYYDptwmDixzXeuG553F6heVkKBIvfvRgwSL38zdUUFknOtj9ZBysp2GK
wiG0PvhSx4JIJd4dKDjNYEbvxZHmZBKzws0CjJQLupfXll5V3oFR+31SfejDxKkEAZcwlwAqhSLH
JGO27fl2AUavwW7OeftSGgSn/XHpjWY/AWTvM4lGRkDZGRPv2KPu2YHBVFYRVg1WM2fYVb4hunAe
ADtidhyb4qLA6FhqJHN6VcFZaPuNGCKA0z/kTQ0jNgqYiwaFiwCN9zifCjeOolAzYcqd3DoYAC83
r60h4hy4OJSTpDtmawYMccDydiK9cg0jT4SqFb1cIq2KkslbBZgdOkVsCWSBdm6lmwEXVAUr2TYR
CuV8FDe3EZqSt1foF0gIMEePastH3AGM2+lYLs6l9Xg+XPF6UdYqUXc24cCVJpdKr68zy+aoYjGK
chD7nhhSi7rMla22NYfsZ6S0Mz9FGwxf/SkzwchFf9xcaGaSJ73VfFgi3b5WtwflSHwdaJRAw36w
Gp3Sf33//0z/dX3fe7OwFU6DCtMMsSZv7B2ptrpHckHgcnCICwolXZNQaJlUrtjA2g7IlFM3XyQM
L2jozsbBzGUKqCXvkb0i2Hie5S4+fXokLK6FqUY4XQA5Ft5fBHudl9OQCUXQTZ9U3RQsVEtANt1b
4EJJjvb/3HDy5YryKvBaQZCEesOY81bonEMtM1e3T32QDcNzgFbjg7d+At8eCheHnYTBKucGhZlI
C1ADRO9Z+OHNqBHOBi8SPpK8LrA3mBzdep0T58A5Goc5P+SGsQcfMXaA4P3MmVLqudrFO0LMHeV0
lKKBwODBHE2LOeqdgfy3REQfrl14phF1yttUK7oCdi49FxjchNhmdlT7ytdndLRUK1uXFaSUi5TI
stM1Q9TgtWef3necpP+REIqZvmGeM8EGMRhcbPWT82nLqZYdu0SduNeRZcp5ObquQTMaNxiag7a0
E3qWO/8CxCKukujccEUEt2KCCd9YYkS/HIQ6jS6KtASYDO2ODz5G6cUzBr8ZYWMQYaeQIZtj6zSH
axq/CmkUtZl2pGbTOfLiMRhKDrR924XpK0JHexacREzPDmNWgd6v2xmt1+AR587/PBP5PQt0V14l
oKaSQYBRl4iYWkpW9AUBN4y3BgCl5qL+iKXIx45GwHvqHDlw2PUPdZdkRR1docD3IIskyxy4a5Qz
z2bIC9JJ7vSlSzFXr8bFW8gjucy+kK1Cwdne/7qsQqvIAx583ARc3i/0mNsCjGIA0vDiLfe0yTxe
2jfIL8OAF9lRMNdGpBzCrdIJuZcZZELuUGauyGpJpgw2PSGAgjm1puToFXEIPaHaII+BPAoyX+Ms
6vdDB46Ef7Flv74czYTC1sVI5/fX6sOBTQ7ui5QAnana7QmMu5CLxVBt3Ut8Bumb5jSzU8J5Jhcz
gLnDxnM91j6cW9RvTNjFKpOH0HeCCrnBI4+a1PjC2FDXe3Cp2JBXy4yAaXVnetn6VGIX+KPPK8I0
ofVPO3p8P32blJmngKWiEjJjD7eQZOIfSmDBIAZqe126iw+zqwLpfcGQhxnhCjFoLzpwAeNbGaW/
z7rXY1jIsKWWOlKUenMWc6gjhRFsJJFh+0qlMUG20K/LDmNPgPYm98B9QRPMx+b5FyjA2Kgr0nx8
s/QiXes+yDBphSxJbxktfuGHVi4Ph1meFE3EpeY7Ni7fjvtC1K9jvYbmmMlauwdo0yoboJuE1kMu
LgFN4eoz+EPuC42mgrnbXc5vDftMilgFR6atLRrIYJK6DqTYKST/XvhJaI8tXc3D+bv3qUqeyKv2
UJr3KbviQSUlBs41vCxCCxDu3p+qURqF/i6FQAmkDf3CH01NGY7DMwd2E0POVhNVeXCXsuX5cdRX
lGYVy7iwzKujIKQorVe1fphe3PM7FlnYdEdd4DKCWyqV3/63IpXFSDS9LCPA4N3pmXgIYQ+l2kwf
oGDSdZzQ2W8eojPuYCP8JDfZEvcLLtJI3j/S/tCmchF9A96rxvpRk7p8az2jctZqyIm7QrAaxg2+
XRBT9kJ2tfBSq/K1HHdMIRP5bdDwz8JA955QVaLrerFtVUokX6YERPrderWebghWiTvg6UpgJchX
m3h1xMRuKucNyl8yhkhVx3ML+FWko7s6j0cpzTTDT/XUyTkkDath2P9sGIIE3PBS/rVkRaBvgOYx
sAB38Wb6lc9+WXcEtxYpbPti18SDPnSg5bXR6UHYuc7DFq1SWIuHaZsf3Z91CE/k3t2DSgBOWah7
0MnTFZitamj7ZLpiFpeRjxDs3RVyvzTrG0ZJcBJx3/+1u9dxCzp1AswJfVXEVTu4R4wyk77WIwfX
aumHrHZD9rW/K6kwOaneLylOHd4tWAsxpeS6xHTbryBZ3hH81NyiLOQHXLofOvUn5a2Ck8edC58k
poOO2dw1Ox2gQqRSUhDUHCUqG6ipzbofWU1Q7y8UVLqdRRlw82u2uKB4xEASpY0px+W09ueRA86c
Xt6T02vEOYUuiD0ZolLS8Ju5HQZyCZh4Zi6l295+vJYYXxMx9oNbyekmqHLPz/oDJkpIMuNrZhCN
EMyfL1ltFqrC7yWrDiqsstsVnoB3oXSmzObqppbbTreYeojuQxUiV8amkVxAVCwnp8zewhSeWETF
jy+P6lcg1U9mH4xBtaJGfm3DzEwEPy2CTKeKTqqDSQ8yH4/+FigcXLK/1GzuyhKJ0nZMRsOmQ7Xa
4L7MLkwJm5zO8I8k38vFqQDC0nNeHRfMBR761TuRd4x89tcb7c0YVNGz8QQTqcpTHBlePcySLTqi
++A/3UC4L/Orjk0NVmxY2ye5S9sCFO/Ed2gs4ZqlMlfLZzb0UH5ZNRa9vnreAvXsAyqO81SiOOJT
YxfWQfDChDOiq6f6mPkXlkO1ZnWYmWBrJBXvDXy1xiAJ2ndmuSIaSuKY/Yq0UseQRJv/ULmHb+bs
lQscqd53FgMevkx6OJ1pE3tnnMSQHX43JgbVdP1QrE8xGwmnpSYXFyo6HaG49NzM67/vVqjHdakW
RdjzutNqrhVZmRc26uSgWcnDj1agS6mb+qDld/vSDTCGqo92w7bZpqhS539smKcwu0euAUVrj1Vh
oExfKc8eR4t17/xHEvIzwuzeBIa9O+/G4MRTTeBP38KtfHSUrvhk9E0s4YlysWLbhJ8+ZEHteuFx
r9iU1pLd2nDnLMPS3CDfJqKrtGydY+NlMvLmFlqKqxsElQHYnBica90zN2nm1xdsNt5ehhE9IS7V
DPOqKL0P7DUudE541cS7jgaIXUIwRk8+ctspcoIkxg5lr+4mecrRyLXafsAz70az3V4aoOVYKAFC
U39siwXVfEsMYMhzo3nfXLJCpxi39ojTB9sBQ5xPjb7jUxWO1khSl0q8USwXTBGBdnrGTONWftSU
OEqBdk+1ZmokkEX4v5XYTBFT+Y/t0WACEMyz6RymUGUEorjm7drH50wU/+qFDOlu1j2KC9v2WITy
iRtpSSN48rsgG0ulXGNGy8Y0cnQxmPP42KXZkn0Whm55pKsGjoYlnVtUcRCJ6K1+rst3BFAPI8Qe
LFhkS8rAKbEuXSvxcNNjZT2mKp3JuJL0V7yAgu0wG5IF6rjY2lMHEI1GITk/ybarn8j7E3uXzoRl
rp/6OHQ3we4ZnxvOv86FmvxSiTucQK5+t7dzxdmuHPtXkesVg5aUhOBPZGaZa/kbr30YxdTfo7Z1
zZSGUAY/E3jgdv5JB0Ezo5kcMKv8mN34e91qNu/61J8qNbhhahCjm4dLR46FNtOqAmLk5pGuidjE
/725182t9BmlZyK3XlV7KSRtJPhSn8CKLgKI6Io/IezP4zuHQ4ia2vvyHiBQ9iDU1N6fRtVboRU4
zv3tCs6ZSLq+JKaYdrH1JZ22u+F35kSQi+YHkpXbslY+1xar7lJvBJjYTm7uUApy9AiPacyOE+SH
Fi+s4mKGvQv7r4jBHTEhO4oXyEkkVWw/ZbU1+9RSJqiKkPqJ3ud0BUkbJOrLEezplxaKATo4mlRx
6C/ED3KDd94O+QAziPZxlIy2v4HV7nPyeeC8YHJQtrBkJrEY1U1/aZSBnvs8ElJuZT/ZyiTRhh6C
4INzAiTz4y9pNzVayh3xoseClxE+2ITCF41VNhhsm19F0Tsw6CL6v4ctcojLor06n6szUbDoAPKI
hmVTOsAz4FqBkGWVaFiIHbKMSAzWDK4uIbpiiWQCsvfnqVUVvlJEn6iCpzD2EdoQgXLT6ChoeNUX
/gZMcDwI3MjzQMfvE95Zh/BjXJaDNzDssx+vFiOVw6fIZ4rl972TODfDV1WsTxdP8EUGMBTQuMCY
1c70qgZwy/RsHg3C9SmoURt51/lg34rgVhQBCetGsjWq/h2YYDwn1jnXedq6zBAQWQlWIlS4woY6
971pRERRIYatowUZMDbC5pJpXpv4b04bCa7FKsef4SZ/JFDXWEPnLBrb2PlItUeWAWAX05cO+3rR
YGCl4n79Kl722yJO84grr8a+0YtMZVjBO0K4QnytZxRpG1h5GGQKgknaqCQ7pGF3irLmgNIyJFPX
Brr8dX7ZQrbT4wcKu3o9HUCfNmCZulYcjwGbPDC/EVcqASZtrq8FWAZhVP+j9yN2lqT3HeeoaPVD
4L35tqYJyRtmuWceq6WhCQEyc4v9GGaCjT8b7ohfW9s5chdXk8aNrhv9HArnEPekNinShXPdlQYn
JkTXlOW3PRic9nkJRpPJMcRlybjbkI9noPfnq/sbAxmMjaBVHBzfb+nBkOHg9yy4XH/YX8w/uzF1
X3Yu6/PNtn0a+eHxIs3fyNl4/gGJTFHZmubmXymNBiXZbn3OReY7Ui4Cgmz6qHyMAKaLGPSeFmh5
hcZGeJWgBqmLCr2f4Gb7gOCy148ona4oJTxP2ce1ao7M8c3W4an4L4b1YKTPYdHy8bzxh8n4KNk4
RjpKylIcMp1gEaj6kQ38ydVvAAcvoOo+kBoZdWZLhwNQsMAxKrYY/I7U7PPF+MSZ6GgbGKkMgq0E
kN8vbdk3I7MYy6i1cz5a+inaULDoXSg3SEAwtUplFfltmnQOaRu4K5LNpB0zbTFt7reE4Qe3fSzl
iMGBGz3gx48LjzeePGoySMK7iqoxeQ+94SCtYZygtgJW5EMacblFUVUn5VkqfCjys0FS8UHdyBbV
LyR1QHhfLu7WVphduuUBr2S+GPdqQl24h6naNnu5ardCBpk+XS/hF0jvSReDBL5lkJq4k7r70N+f
MIYcXzQBXuwmtsLlYTh65ZdeJ8zQn2tm9A0iQPnBw0oEbA3Wl+YBrLxz734DX0a0/OoqGIYPHscC
ZF0JPMkqCwGHkyhJBTZgBit3gY1SKCisEzjQT3/9auhWmQKyD92fqecU0q1DfrICLQcT/GOT3L3b
HqFAFvUYuuuysdcaVf/9TnpuCRBNVmMyNZ9qItwixxMtkvIuw98HuWHADe6sBS3WFL9Sjk7abrlP
V+HUCNYQ/+z02HpcCoM3EYMCtLifKgSEyKjOcMnSnkz1BZ6uZGu2f75jrAAnoo5ZNKy4ojpjIbRM
bjB/v4YjiMi4Ydm5qXuJvPjU00E5MK8x/nz6KjstQLyDuoJiDVnUicS6YLt5a2vNNZKZzV1pgHow
Zt15T0OVUfXrDZ5yUpHLQHUBBihrBQbAHh/Yx9VmjLMIbDU6mQ5zv5090gZdSwS5aYjWRH4zRhAQ
a5B5bKKto5F/7QPOuBfZX8ZXfP0uTT3Ngr4KlEn9PAThaEOxDGgHNrTXN6t/JD8gUORr3LaaXzLL
BJkUiwS47XDNBvwWxgzgeP/8AHzBq5RuivEKJZA+jjFw1s2wXHfzHaQHSrX61VmkjNl7ILHXJLwA
ySTmrw3SAoZ2HmnNIPpOitjS6Yr5yy9lHX7/fSn2tEeOavp6IG7U3ctHHiUfKTnvIwUwzxu+CldU
78EVBmZphjdNIn9ZvUdXhFH3DOb7+6fgh+2HUWrCa0mWJVt2pjUeegFAx2X6S5rIAF8Y5nuTCYZz
WjZt9wwm0xgYe2d1EcwzvDy1Oo5g+640ZUM8qsqaEgrEW87cv+u4C7nezPUHX0m+vO5QKDM+AFDS
Ma2fohxxYYtHKitjzxhJcshEoZsEnE+gPQyU2q1jFDh2ZaT//SAwTN6f+KiQvKnjMXQvPUiGCqic
EdYED4I69JJ8c3v7q1sesP4eCvpXU+bsibbKC6b2mtLerezwEcTE5df/ppcQL8bJTXQ95GQQ3R10
l1Xw68am/k+pIsOfySrxld2sfuD41ibQMfFusiUyIV3pUv8y9ErBuQmrciIqZ9AqDtxYGya6+RXI
9OsaX+kcuiD6hSbsoe86DjW/UvLgN1058idJRJnSSmg6ZCxaDUjOwxOqvRnqCJ/gxP6II2fwqSp1
C/oJOP58nLdqx/xdVQRkahsCGMTXn7N7OUpXNOX3MqkXXHkkKtLYE2LpgKo9cun256r1Q3NnVqae
9Kjvc2whGU0reWXAYZPVEfA/cR0Gb7TweWGalN6bJCj3Z+ynoTnVKPG8CQjToptpbb6wH7hePXPL
HNubiobp/YP3jaFGqpkUtYdVJ4L9a47X6JCh/uP+/nCEhQdR18+jYBGxfEGsyhlpTZruohDL2/lJ
Y876pmWKfgFjtPisnAllZ5wge0AQyjbonNigyI2bUC/q66oR8HFVHOTqN8qxjLi7gw6s+BR8yieN
fXOCxjFjHrukZkO5cwpGemiQUHtpLv0O7ZZuiUW5YO73PwsnEsPR9MTbS0OKwhANO3GrNJu67aJ1
Yq6i+TlYohxu3Xi33KkdkWVaigJUZpYgOWpxsL3bFU6QzXulEpQKnWzJx7SokdmEo3bVH6U/Z4Nm
gpIxVqWMkwihPcKiDDIUOT/nA+eh2wjglmSyEIGwr67R888sEIlQjFYs40E3y7fa3Fst29RivliC
FlHDdZ7BTTaOQ6IymYxBeoQsRx4/+w7nWpy4l7NnQr/4ZZt165mr9uhE1RXlsHfjmQI60CGIoRhm
Z/MPfibbZzvQrbRKxVaiKN+gHMEb2oSCpBPNofQqv2m8XRG8oxlqBds7Ua9RnWPb0m8xWk+Z0QAf
J2g6lu8+JKjD5I3YZZOs8HCq/3BrwemgAfcuqZRySV2ZYRg0J014mQjp7cPLBXok5r1byBESBT79
7GsVWgH0DX55cj8oDRqOnrgRUKFaY95Z8/PqI4KwNnkUjzvIpmqZDGIkLInj/SGEvl9p9Un9m0Mu
L117ydTXGGjuBVvKrPiUGXU+IWzr8VEu9/m0YSbeYJUFmSIigewGF6ih+Orcgpc4U9XKU2KpvAHo
0wudbCuX8WYkwc0m9k8fQI0OlpImsz6OCseBDCyCG6sibI3YzuID/HG5IX7mf+lBaQmz3ubGxoEW
PhPVj8S9KbJZslHdfipQD8qntYwip2/9rqB9kM6hiANCOooaReubzcE0OFtj4xVkD1sWUfK9LuaY
M/bN5GprUqhNMsa4VblXpjFT0l30uaGCWK7m4vBLKyQwMCHVD3zJ5YPJHOnV7fwZMUrvoZ22/gYV
/616vdydUjOUSIzKhAMUhbPKV9v33xODZJlj4Qt/fSeDw1j84Aj+9wVW36sJg1485EjhYutRkEwx
TK7anMmjjOs04hgcyPImaC+CtHh8CcYB+kYpksvsCsvsyXzHzdyD8Zug7U7i/+7KKFrqT519YrtG
OjRtYtvn1X4JiQeIaeqQBD7WzZNA5SG1Qano2yv1JabkPAWdeWVZuVN3d7PWvBseq9SmerOVZf92
snrA42tROR1FYOC2G2EZGG0B8r+aejQMNBMzAZgZKLrzHyicp/gdObQ/A7WFyaiWrD/yiIbxS1i+
A2xtFh/D/g9R+Qk6FbZ70B7aMiel4S2QqhbhsRmW9TXZgARhpQZLIIqbWRP0gzyRNAEKFDCJtFTT
jEfw1y4iav9koWppwM+sX6oV3kwAubVxGP8lo3SHPpChO9gVRZODYncP0st8UMAIj0XdZPo4+2SX
cHuRiLqF885tiUKTRE/2OR6HCZlEVdJgktmdFTnZp9f4njnI7zARLD4hTY9NzVCsJU69RCwvj+qj
HEjDWfobxscs0FygJjOVbbmo6gAx0D9XIK3gYr0L4AAhWZhDht6N54L67p1zj1xYIOUve0aLbutv
08RyHrK5RcqQ1NcBXiLkLPx4cvFXGHIOe0EPr/iUIf8fnz/oQXo1hFPl7vmR40RFphozWvpg6IN4
D1rTA5SOXWK5xGBz4xdwWG/keTHxrPr//kocgaDbJw5JaST9WxZEbA3guAeLTLhs911y/V+vltwP
tjGu8aa9KYEiArVJ1YQ/X7QRi5pHV9CdpwCG90srV/PeWUGz2lLBg7ALbuICt+shMLL+7SyhAlTA
DJQVnOMu423CZP9vroOpuSJBNpN6dkhrhrVnaYpaAyTcNukldVr+Ha1a2aCrQBqJrQvAjSpnzqUR
pMBcNIkgTCjzyEivXnJDRo/f8OcN6Pchypo+R5Q2VhMHmkitG9jR1Ys/gYDfe/J0DjEEFnmhEoKv
my/5DlknOckc6NeRxxjCgiYMoriM+1ETWFw8jS6pMcTVB7lKHDKvsgmSTXku+ORN8M8aTXA4td4d
f3lj/ypxWyjaSMh1mbzpjIeKMrFwCcTPLGK3YIEFQongJykbvVEou7T1ESjsraWFibRKa3fH7bhS
o5WC2+wlwtVf8Mku89I3UI+mjg0OR4SbYrW33/7s1nqvygiyMsOyl1IkRdNkjzNiIYTi+ZpnqBzJ
Vy0+aHoA7Do1I0dsFbk+Vzs7pbdKkWvT2MQAqZ+mZzbcwKgPt4KFuKlRijXUyU4m70h/LJBBTQ+L
/IhBNYsMoN4jcAZJHO8FXxn0vNmCftHsFVpls7HnOKaDyHeTPwlud6bIvmYg5CJD1hxntW7YiQKa
OD5qRNcnCnwc7GSrIX7waxKF4Q0IQWmUxXWt/HJKAStzE2zhBDpN2jvr1upjrUdJLmuwBZ/Md6Ac
5cqBQTgSo+4MPxdxSS26AgfXAoWTdNOi8Q7Anc9qzvN5L4nY8SLQyQlWAPKyYZYaN4/IZQh6lLdB
aSOwBUxltZvp4OfmYLUzGF+f2rVM/Y5napiG9tZ6Vu/jjPeFEwYpJYOW7FnCZ5ieicTcIpL+9Wvu
MmlQ74d/d8vq5zsxvw/Ef/WFC3bT8lKQ9WeNesds9H7r0E8W2jsBrIbvEunndGzMQbrdRdKhwRlO
BGxGF+r82inFti479rmVbAwgk6OZa7orfOUIKryr2989gMnKMcIe956oSMj7/0izf8nIqNYbPoRn
lmKagbaQfvWlrr6LdJQTTMoHbhR0TQ0kBObZOxmHQshCceLWukkLLAW61JW4/ksnc8KyJaZxAXWl
RyAWC/9xL/Ne3h3syS2EGMphhXDs2ZE/Lq97jkbJbt9kAKdIQ4k5lbwrxrO3BNdzOPu7va5LOEyx
83KT1BemApL/pegVaiCYWqkSX7hstNHY1KTXkdJDyJXb3ysPubQ8hv66hIjWse99+UGsAhjr5PBh
RoWd/Uq2U1TkYD6BKSz6gApzlCsijyv8MXgD3yzVF0Y4nw+HW1TnST2Qc4fSqu7YbMGOURWMQuzs
bcX/Psrll5vZQfJ/NQOmP7YHeuxCaecDayKVQ/yU5STc0Pajvv0Yg61PPwhp9HczSQ286+WbXDTO
g88ddZb+ho+hdtt6J3mhmLBHoWuULYXvvCfcn5SJ9V2xdcK0phUAjX16MudxiYeqxwIT/cDvM1OR
z3reXEOqM8AvGUvIqSWUEAYOwF70Ix0am/5/uXx+UAWlYm9dys+IGMBgHdDRB/PhjGJbgVVFskX6
AjsPCWBtMVq7mKkOQgZm6Wcs3/qqaRaPSULMnfMFpTEHkgjyGKmdkyLGprSSsq6AGxyfpKaF0slS
zKmO1w9ZRYvK0fbNXDayCcoabJsHjDs1jOyXyJJC7nYQCMX2/EItrjgobU2WIVCgsYu3p5QELTlk
h5GxamJWz3vyfqfqyntyPqQLSmvpTlEuOi/3wiSvdcca9ggVTVh3/M4Po6U/yaGM0WsUlB6uhHgg
kQDZWXUB7OB3sOXC0S9n5VNJcrQzabx16CCInIp2J/bCi7frRE8hu4tuMWHn2WUUE2bJM1qnSOec
sEL+iNQTGW6uTmKTiNjraxuujKhxu1k63hay+68YOjRAuzcVceZiqQyXVXn6FSvGILEM/CPgKpnZ
262MJvXfVvKHU4Ev6MkqgDBGdH9sYY5ROmTVfsiX3g1T78D0bhBtVY5L40ddXC6K9sWVT65TfuXX
IGlNwERfJahD3l8N0+TjmMZJsLpXaxVREmC/JJhKaiXjMnjaFKbcKkGSVNyg32bVv5XWfpoVwE5/
22PYk5D69U74Lv+d12B5NGf1h/QAco8ioVZkYwfnlf5ApowJ9SjZpA+UJHWvTnlV0nqf5yqN4yb3
OS+b4DPcYlMxN2dhd3y7pqNcLtj4FbSmuIDP/ERiiVhWV57FETX7zOhFcyIuqtW7lBhDJpr5UffU
hc0tTygvmghzQKXDChTLWqu0bBjhMLXmh5+rMUv2IG3kLOBsSX710SsDwMjbp889cEsLvyFaddAS
VvJInFFL/97DndO/Z1tg/II/ZYhTcN2eskef/WJgzXGpBlpYZaWWh0eqD/FWGu+6RSTeRdzneYYk
wzb28IrmY2Ms1GJixK4kPFNn1c3SXJe2fI1X09jATIngZU7yF3z/tuZWIf77kUFkBG09qNOb4wbJ
X3IfbH06wWtpJQw4SA/PjO7u5Yl53VJUahsBaybN4kBDhAcT5LDDz6+T4ca/8HWSIb34psV9QfJt
nCyaC5PThxg+0ftTHZFnkj/XTNk2uwZn0h9XafCvsMyagDeucwAq3VoCHmL79SMvTQQQV8/ANVmN
3irfyTp7A8aLy8Ux5WEkNg3O/6co5z+HcPyKw+0dx60r7YShUQbCd49Ro3bEbLQxFnysSv2NYecy
qmcP0ax5e3xAr9tjHnJARWOYdS16FiFqzZ6qTF/FsO6rucIJ1qHjDEoUvu0SOLtYX5pm+QriXUhU
iOX+990vuXx/NWyEFXZ51mvnC3Kc0cC2lsOjEoid2LPXkHjVBwksnwBWudDPlAcNohgO52QaMvl8
YYHtzNkrTNC4s4jt59SPTjuMyE9gGlE9ITa/wGSg1r3IbhbJILxoK8DT5qj31dd+XfpleMKzygZn
75S3iaRCre4Nb/4yjJ7Ii11+a9SbzYyKqfIPW/ipdiRtrXBD5HSmQTyS5OJk7CpOc/SMRah72HtN
EC9gR8hhLR9uAhaoiDuRq87YKqm4Y5EOWLKAgYd8Z2EDwwpLphHefMfWHhbnkRbeRUYbIShNFd1i
RACVIkIJl++7aHtWWLF3yd7PyD+zuvbLRNPfhOv8e5zFT6nLspWZadbHDd2llaYH13uV66GVrWFZ
p9Hty7Uc3ISRWjxqbdicHwZjTYQjebIBFTZa7YwCjlQ25b2BS4PhWJAGESzE43eI8tzbDK808viH
8n+vIe54JjaPDEXIa5b2q60AVPUf22n9reCBexykxjpT/ev7RRDsi/X9ib6dw9SMoPp85Ppwen83
GuHGfbxVvEcz35wLDwlITr1R/Jb1q6FPvy55IaHK9C8Wv6wHswwQwTYE+uVckMFBGMp6Lnluk1cU
WYLsrw9Q1gMeVKnSlg29zIOVfPACZZikdPa9WnFfs8G98wlKqu7oaalyWdIG22assucoYXlKIyyX
V66ko/Rw4MHhtY0t8ThFRJEpv5PpfsWl/PhV59s+EFKsEjxitmcE/nuwbXHDeKWcIOJAYzk1R32c
AGy8Y8ZqXJW4xn6PUFDo2ixb9n9x/4CP6Y1aKOaWMovsMAx/ace5q+rkXWfSDCGNfU8BZduZiolM
24LINCO1scSqynCJiZffFuhwiUOFCyjK9D55//zXfkj67yNMj+YBhkk3AwZjVbxnmE+/Re4UN+2B
RfUyFeXJ7QUW5kE+4ncLdce3ONxCDbFee/d3/+chXQqfOq9k4TMXOfYcR3vs2D3aQOblKehZR9V8
YnFxqPIHWpW25V9kIZzA3k8OSTvghkcYZbaFyyfEFkxuC8Q+NPOJ3Ap6dXYSPGJUKg/bAM7iX3Pz
5e3gS5UfZmZHYCkT9NFssXaOvKYJ/IPWPVDSnRQZIYzTWBjBQZ0NxMxbD4pbUkIxVRQlkr8MOjFO
zZX7NiWVaAj/S7tAcUV1PQ2fE7DsuiCS+dQQoi5W5B101q8LUVDxk9/8/pyCdhURGITUd7nR89pB
dmZItj32GxQ4N8fwrHca3JmRr6NZPlKm/PZeYfooV4bnjFtDxbPnk1jHx3fDe3j7WWRi0D6dPbfi
CtUBEDJRgBI6RSyMWF7XI5iTzRUyGpk6BoRn5qjn/J13tKr1NSuuEoJfePJoCllruggsRAGBYyV9
BC522zjW2D5k8NkM3HVoois1PTOFTLUMok4ffKELtbKaI7t2GDxPH7y0XYzLPRypuViMVuog/2Uh
mLTFjLdQFy9z8aO4XvO0OWR+UmY5mXaI3n3t4idPSR1N0JkMQZ+p65fAVg8S8ElHWuLv4MK33rEt
3NeR+++PQmGg2+IfZXbF8NsijeZgU+UrQrJUcXyDBiGREkFi7kamCaFbNL4hIpaFV6abtVNRP4CP
Q1dySkvlcQB0UlTeIzKrhNWa7uPNi3LsdDrriCo2LSMNO7MbM5QjcxWzFCRpF4D5nu7dLMIFvgn0
QxqLFk17pVNwV7qMKiSky+koAHV4Pwe4u8eHg6FxwE9y/OR0f4csy+/IUQihPwOiQJkpeI20rJMY
TYyL1uydr+DIQYxHqxGTMbHzGxIxCuQO8YW3fp9KYWrHvlQ9BG2tlB4MdGKXOlrTl6tqdb3SLiGV
+ml3BKTqWmpIO5L9x7jCACvwrlb78FnoJMdcjxy8lpj3B4tRbdhS2OorCwmGzdbaBamBKA98vakp
5XduoJwX+X/JL3JcmkwswL3P2FXIJzPdjbsrsWr+s2j+Ljpm/8ZY0dhMxGFdfMiI5/lET8nTDjsS
EasnoEv/9/V/InQ2cL6OES8fj5m2uTL/HLs0vq4YdYFfzhUnTQBuB6MLVSVDhRpPNLNwbKUfreNL
G9TF9NHeFYy0NRp8uC3N9DguNYd7GUhBgDLXOTqv/AP0sz6BspMZAEOWFFn3DOrEWU/DEiTgt6B7
v0uikTdPcl2ZJw0lYUTD5WytcfqXOAHPmDABvRTd5KvQwuqKxrVfj4MErkdJs7McCccURhju3tMF
LLuSY7CQwA3vigW51XyZDY3rk6qn4WCNDHzKnmgngl+FOJEyufkfONSkUzzWhP8dB9md165C+qgn
SvRBPnSZvWb3rDnLAty3nDKEAkn7Aysbi7WCvEu5gK3tfeGitU/WUOkcRi3oShOCT1e9b3vNUFgM
6j1vQ1mbVL1405uMGJX1kXfZE833AbaRtGXnuui0KtDx6KoqCrMQ2SqTNDxnB7DGUe7lSOFALEiu
jWbVEa9aXAIGIHKAJKqrsnISAtdkxBJwZSy71v3Prmcn5wp5iUhzpzBiSEii8hMNdNbML5jyV7wl
menvmZKpxcxIBX7zfkT04Jnz/4MFgigN1ndhU3huMT7+rDWDkHjn2pRqSPwot2pN0X1QnN8otCbW
cVHrk8PZWG2oUaPS/BrSF84rBkZZP+sTvuOrZNugI4DGBVk+LT1cc7iCWxQbtWKMQjLG1YeFpl6H
SmUn6eVExzUEqTBfCIjdHhlgBRsgcNk38FHqY0/lDlVZGxZyL1dwr44VZNUhrGT1RpF6EtAomhB0
wLgz/UeZmVPxjKsIp+qk8BcaO79XYoOMY7sCbChKJBvXM8gHBka/h162Xi9IfxhIWvGdBXqk3yc4
zRrJNGQpFZub8hU2HYGAvFh16m0CTlKyyulyLGI1Iw2eGD2AXsRVxRwX+uzGaLgdeUBAgLmqjVUX
EIN8c6HAKFw9TVbslc9fZF40vG+6pQmNylZZfjUDFEQDvzVyRX8rpoObrJjZs9NUQfFoNoZ6vCPc
GroWoeilnzatwghjMiebJig1aJgv7FsVXPFj3jo6K9/5IU2r13QCGVkjJxu/N4Tu7siSd6ZfdEvE
LvBH648bcwi1UxZm2fR8QTM+d7zHKKQMFBf1zQ6zTHw3f6k2LUYIOd8ABMn4D216qq8P5Y3p6I02
cCJ9IM8obLmwxm57vWaFpciU5kuN3WzM3bhbEv20SBd3X5nEXGN+TOQteSWfKEGyn5CiF1wWFSgV
J+NxwBhySFIGBT0F6UJ3z0j/dj3bHLRn2uJVQVJuVhp7+mOfREowL+WlnrbI78GAHLkQrXMZ7j93
ehl34aJob0FZPfzAvp99pnEvh4phw8XXmCpwhyWV6CJ/D8nakU63HwzxQfHhHzTUO055YYwtGyIU
eCLBNQmRXOFayDiTsaesjReM5uHHthj90Gh5kQhFk00YJWdK259h/E7UGuf7UUdLw8wWvjhy5wN/
kV5ga3BXreBCzl9WFTJqngK0HVGu2ZPcJEMO7KesOv/pfs3WjsMyZut2+sXSi0y/5rnmX+GS+5kA
dxRb2Rbw5IZCqyGbST8lTT09wu6IzvpjBEusVNXAeGqEijYDrWGw56yQAfB0/hvW1I9ssLZoMxDF
GLeThE3VLNRKOzKPj37Iqu7aqUDJ4Go8kPNMCN9q4ZbUPhPWh3u8AkAdu9ZWAaNIZIE9mD6JKcVn
iKvZRIGj3b0tmQQySbAoNI0Exj/4drIr/urFEtHVByDKEechSGxxdia0cFXF0UXXdp+GvX6FQZE/
DfmzChAk+Oc3ISSRGmC5ZZA2X7gQRNBb7H00FlDd9+do4o0oe+Wit/YqjneKGQh19JneGOyrmhyc
XvqzQp1juKMswdwFMd487BBBkmIIEes8Zhxw/WiI+Uj7k1A/F4J/m5MGXBjkuKQIWgQjB0KA9qn5
Jj05fLzCGNMednv3sCo8Xmur6LQyP00Uyml021ymkv9Zb2gtjj3C2LN6LqSMa/eMlUL9Uv8gL+6y
Cl29liBb9l5xwSEWPt8W5DDG9MoUmB0lbBfkaB2gU5e2bzXctsVBHoylBOUOJNkIpir2gCCmGhh8
HgcWLncZn5yGiDwR58sB4dxDXQbABKQ2rvWoP0Qi32nJKd9M65APVxyv7yn0hHkHaHA9GrE0ZhCo
HGtBDniwbcL1H4kgWGIYMmDdE6R+BK+uuWxB5jtKaXtBmOqiWImMw+9s3hAeQ2Vym7TEvcuv8RST
x9sQuKz5rRBTVIc/qxxJ2aUrwg12yDB8DgeI4fNFPHfJEDkJ5rBUAXk6AtfTddddLzB97n6vd/Ng
QqF0undSJ0s3tXEseVbGiG79AVkpyj/f1UJ/HLULKvBQVE/OpKhiyZUiEp6MzFfX57OJ8QnegGGZ
kYc6hU52G3HLHr6eGchbuTmyQ4uM7GVnpu04ZRMvuMVxva98fhPYGlDJQZRARJsDAddTIbAVXViF
VmhwjNd475kvAOpPTMqNMCHBj5Zj0sh63LBKtZSSnkZWPhhJNCc8/Wqa07tNuM7eT3wT7l4UC7vq
Fg0iKTDJC/Knlp1ok5rjJCPtxf5xf5IGMhsEXTwlUEA1Yz3ueIGtNcquFFmyKg/A29JQNcAZUN2J
umEnbZHDLA+kpbtMFGJBDU5+HHG5inBD6YgCcZ4czVnsgc0+Ebemyk/tjbfT5jU2yfp25vhD1qBp
9iKERDIlKk9xUfDJN+lP+BjkJ3gBODJ9wuA4u7A13tbkci+tolQtbwh5Zzyu6VkWmairRmfmkfdx
BY1fnaxFb1WjfVx8xykBLVLk5/O3Xy8vY5QK/2q9OqlG/h4cAPrmm9H2ZY62NrCvfQv/XhGdnuM6
f73zwkTkf9FPjbu1rNZzzuUmb+96kHL4fPgzruQHDceVU9zBemFaQn7cmVeHgK77UJSEFWZXUz7f
aUUsbUxpaEEEKvJlxttqWWwMqld5p4DzY2MbyXFCe+hL5au3e+3kuEJM6ekPwA+UXLCL6zPou4ce
2M5TpM3IdTstLX0JbVrczZedp3c/3oVh+JD1hk45KH1jq0o1nSK3Tfv0wKd4V1Lq1CAWFHpRpuHk
dy+5FGqZ4Fcv+fUKJweHSHTXdyec+PHGpg+yC9thn0if0A7fGNi3opmW7b0p29rA5LyfUwpmZ9Ts
7DJ2AHcpxavtncuKTUBKXpjydKmeDGGXu6vL9I4RPviej/kqrkWOTwATrG6j/rqympz+mWMqCJBf
lJpUwUK+rHWeBW5VF5Br5LwnN8q6ezXNS8u3Ac/prZhpkkwSBdeaMyHy/EJpDbuDL0DwVf0zxGeG
0G7E3TEaz/1VhUvVg+QF4Ms6bLbLJjbrL5Qx5ggu+HNlAZuU0+qaaJX31gvsNmtuZGVw/TNoWDTv
qI3zvFAhVGWSMPbW8eg7Yr6KgswZbf+SOVHJRYAu4hfDIZYvW8PMD+4KdeUw22IsiQFcaO8B7u02
2X+qhxOLqF8TNkY/2OpToRDE8miYFUpTDWg1+y1WcxaOymikfusDPtn0XBn8GpZxXGSmYBQlqXa9
ONPAs2kPCBW8SmCPPni62dAqoT4YVks9KvMiks5pNZ2VMVl/XwgLqRaLrSt6J455rQ5Ddi9atbmp
l2OWkwWA17FJkP1wTIeM/EZZm3MuZCIl/1KU8Yly53qJCDd4dyzRN9fS/4roc/X7IXMAu/um7b5S
mC7Kc1ylrdQOkUWrblm9+Ifi9xm5Idwf+gfoXeih06peBeDoMVKuYbcvys+3XDaQ8cHvEkCQ2l1k
3U3xFBtQMZdEcww9znlhzGhUoGKTrSfvSq1Y6a+AGLKt+LVKxWI6fnYJI3g6qGmr4hN8zVBwp72T
6hWJHjmAFrIZzv1awDEl2y4NGkaj97k7cwcEy3uWJ9gPF32IrqOVjDr9WZ48DGEuTpTzXqo3s2Bb
MD5cO6DHEUHM38uErCnFZvO/FFofmmTpsNiJc/SioE5hHzhMEc/EdVofEHj1h5WTr5wsFUI+A2Yr
nsLRzZKN9zU9btBx3GzFU3FFxzND8Q5gdz2eV+A34kO9mA8J31ge8WagPl1TjVQJNchkUDkXS4Ng
nQzxiWqy2Dffc5t/RSgpsLVVFoRjw8d7y4WWbXJ+es2mBD28bVu0pjFS5r522p/2FxMFZb7lOJid
CImZo65nVlPUDPA44fjXtQDSqVJ6xDf199Acjsa2a2QCp5R8v7R+W+cMKi6kiwsSX5k+V6jNj1Hn
iJAp9Rfz6b1DBo1G0Pqnxpkr/04Ok8XSYFm8MGTlvE4ylXoN3NxceSn2ORsPPgXuGrMrB1sMCo2o
XpWfsKwoVo5lFLQcQy5RtsphZvSER0oYPbe35YB71QBL0cC5bFjFKRPiufikhjRsp5+6ZtSXmo+Z
Uqy8m+2jtm3N9+gyLLEptE3vGMw984pH1y+kiM7BSUCxqcnPzRQmDjdaz1ReitjFyuMPfI1TwpZz
sVzZvQJJBa5etXsIEm3kHOwwNEFF/BijKZPjc1CkRUF4ukPGkk0tTOgVsuUwqqlnxAzyydVXpBzX
XKT9+k+r0Lt3tl1USZOOYi2z7iQlIgNU1O4NnbcbUtxLem03xR3DxTXuudhfkM6+/n2L+qOw0iB+
bI+a9cxBmFEjK5RCwunS0QwyK9KX6hMl+sXdkEe+i3mmsNMBN4fSAY1FX/rHa16b4nsy95p7ib1G
ipagWQBoAb9xGtSqg40GClZPWN+69I3xMojuwOX9CMkVoSNRmTmdidLarewxYn3EOcctFLD81DtP
RazhyJtC38naUNcxmkuibezT4lik/udyOPmUKwfzfs9sPkju7hJtsZllnlzEppwLSBoVyyj2juqX
/vcUPR8rZSxLDkJYlfmF0KUUQl4ueyjGpnbl4yKVw+KZJZdcJ7lYK8bb0zvFnOnqDtzEHSA9mWE9
rQZhZMpGdtd27je9M462Z+S26NLYGdTn62oh8Tmv1h9D0mULgo/qhpWvCkssQpcH+p48/3U+gpCj
En27bO3fmwjg1/m0iv5Jfd70ZYIqUcnLYFqrvpLBlLPjcQahldZgdIR3kTO4BN17xzpVNCF3hTXb
TTtreb1sq3lwbAb+DO5hQtzbeIzs4BSBjq8kBOGU7rVzukJsYWw2w5f43s4/vvsSLNkzucZBmrPe
qU3n2asU9fl4oeuE60VtA8pVim82XSwLewXVGCrcskGTFzkETmCjRTWGESltdGepimxO0Kyzs2nL
Q2wwBj9VCk2cXxPzbPMeTc/H4paPQirNjcmhEVxZNCck+JNEA5bfw+POgaj0asisZRVQoPOFz3jt
HfxzgZimxRPd+XOvOunKQvtCrBbJOUvj9GgPcD8Iuiu87IiGmX5sQXj0wnwESg3IWF7TG3dTVKKx
LU5fdPu21BOUKSnaQNhl+lYeflTGs3uDzJQIS5TmHkdQuT/LUIosOLeDQXQnemkUfoiz1vZLDcei
heL1ng53008gZQ/1yYwjEKcFZC3TPKrGKww1XRqKms3hrOD8CiDSkUo0oi60NFAkY4ce43E6lqxv
xiXp8NglefUKb+qLky+VGk1S71lDANXlyBDnikQL3n9I4nsRJ7lKaNe1LozXwi8ZfL7Vc6NeljdW
6p9T4GDezbQmL3w85RMq4pOh5DcWmeA2R72VgYF0/A3p4IhDCIDLyLRxV7XIKYtgkvUmCNLr3j9A
nIoQLJ5T5ItjxqWwNXW91UZpFQRW5rgLy+rpEB/ua86Brgg6w1Y1KTiLKec/uCdLwBVCrnayao14
SbwoX/8jb87fOm6KiGGhF7zNl9teEanRFwDlmLX4Pj/XJenQtTj2Lfa0++olbUX8A4HXNsb6NhKA
7lCbsxuoUeVPiLUFfACIRkquEEpJHxTYKMW5OGkyuIFEQvFPMl3tlwXLmsxKPvzycsbi2HIos0Ji
2BhEAX6E+z9SG8ddRsR176MYAxteC3P9I0Ed/DlVJGqmAa2pRm3n+mh3cMSaIxFe7DyYmgD7jRAS
PUCElDSKHtSkXUyX7B06+TpJvYNN9/5I9QOCRqGYH0K7BKyioqyyiEZUsKq59k0lNkKRpxCPCdxN
jhstguWgU9Gw9ShThkqVkGtjJHmiuF5zTp4nLlMz/RWh/0bxODUXCkOq9/cOYdE7qCuNrxcUwDRD
LvUJBNKRCIcggOgembecrugkncfmbykP5upS0bAYWF7fS7E8T/ezJOozuXVTAMp8WuyPDLUTOiVb
Pyfw19TECfsf0T7cbEn4oRh3fGINIDddjPJrkat9DeDadkT0OwnBlBOc8aWMX7CH90MlRfxIiDiM
JTrrN7s0KVJ+egLiCXAZmtRAgClStuuPD5fCLs4D8ysvhhDG3Z3ZzZH7WZYAl/IQF1lRmDigSbtf
0FQLRcd5rpbiM48dXmBLztO2K6uVX3TbJMPI+cbPF9gpCd/PJzvz8zlaGLK5Iga7GVGh09PPVFvI
BbLt/ER5Y1klsXb+hIZq8DCZUtng3jZ9cHUHUZadTjE1lDHRxfo3hBjljIqqbKjEXuk7CNQBODlB
C6oKO4X3bq1zP/+0SFbc25ff8sWtdX3v4xdT39+CzV3sBtL4WePCH3N2SE89tOK/NANeizX1rnMw
AJtRjDVM7OXNg3ZvlpyhHscCGzouIVCW8H1HFb6KkF+SrYTsh7UHq8WhcDdOS1urawx37IOGP1ZQ
NFkQqqPhrKnABaRFmCqXNl0g7ZwrNM1+adI9B/CuCdflxOtIh1woU6dQ23GI8rPDZRXUOzVIEaSn
iqBViGG8GBy4Nss5Rg47+9mQp6eKu7nJKw6EJGhILaKSpVXFKH6oaRMsUIXA4vHq2yqFPb/va/K6
gEMgSixAxXyq2fDhW9Y+k/UrSGL+81qwJ3T67P+vR8/+IazLknLklKVNzJMgrl0SRp8zc5koNdvr
aCTAOfQt5+NYtsiDjjqNiYnb8UCKUq54x3dFfdu0YUoqwb/OrXvcckIz5I2rpl5x4J8FGHLExLTY
bzrJ0l6RxskfCJdhH3k8x1ff2Q35dZsvYfiM0o8n1tYgyc0O8FnEA806mt9LhvGZcfcUJZYrubIq
pe37KjeC2rA7JbYiZJRBPeCdYGmVhESJueF/x1aa2vwmlkHKWEXR7dE3wv+284njYS8tuycPjlzq
YxvDnbQTN6vxVh22OxVz8R9mZghrBTh1QRuHNrx/TfC68kJm0OxRwmvr+54VkGVUKNgqbYtl4u0I
71RlJ1BqwDn3fFzKzKuZXzsWvuOtOI5K3R8bDL1cF6Zk1+w6tSIbFuKx2x2suEZMyfFtBER5m4/N
vh5XsxsjJcJx8S6rN1kH7VTrQ29ePGyAm4wub60cxMmajvL/ODh8INRbVqRQ+k2IOSvLr0G5gxA6
aDIw0jrglkjtQXd65DEz0ybmApoKwEuSFpM5NZMf4N8cl3CTZlhkqh6M2L94IJySmZFUt4EuYXqz
pQoIVC+hrOQhSmvjFGEKxQ/Uo3PtEGgeFHXZX6tmJUmGhoM4hu/M1zwwIOYI8W1+JzOCFptk/UUD
JeyuZFcTTW3w7/xOTaD6z+xJQ0rZSn+9I9Le0mJYlZKVLaT2JJ6ZjO9m5bBY0EUl8LAC12KUVdvR
Zunsv9GmcPBjnAt2f7gUKHWM46DMzqBpxxg0ewoN6YVVghmIIWh+b/wNQjgu9YPKdVsU/DLC0/a8
MG+mF++/NIMe/C7CQxe2fLUw1cTwq3a3kFNx0Dq2hXC9p7hfC79wRwVecQkzQnQ/d4uI50suYRO7
SQ7Cy8BazgPgorauiX4hHAaP5bMBVqkAdsa3ZuIgAWq6NIiGsNWZf8HhT8HCNqQaiN3BGphYG7qh
Fnp8QWRMuDlRPAr9cXS7T9PHZqfIMyxsybnMO9jd7yC4cyx5JiUl/cTACZAQNOZ84GCtOQCs4yl0
XHjyaoVzvc0/D1viNW6RFAhj47Y0D6Fdo/ispFAPDxf+jz+a/IPqKBMleiXPu0X5h9hCAwJIqZSv
WBujs6VJk1NdrDQJt9F9TtuIDAvKw+cZdPJyTVF6/rgpWlAR0ZCw0JW7X3sovbwk42HwGr1+/tXd
uTy2XqlfVL68LgISDXJtjalxdbNSUfv6/kZz3ikV0cgpk+NMgcqhaz/GTfDrrDDbrv6TrxL62Kzg
qfODFjclHf6f5kOV7Y6Foi1aSZGfYLMXgTsuuHdOD4xl5oDlEgcomo9GXBzopJRUygac8AfLCawQ
tFf1aVvlpqPsd+e5Z/ioUYyg7c3+OH2q4OUJXiuSFqeAE00nfx3yqRux7JSP2hnlOiFVkb2Z0T0m
H81rOMIineKeAIO1kXeTmI40IbANURk7lKhoMmXg8x65X3PvYLoOu6voff//6LMd/pZSReWknlTj
h3jh26Fbh7g1PyOhxQk6vt4FZjSRMiNv52MbWVozBXcpRzIm8iVyQBQoDd2rAnw55JP+xdl4FxDV
iZC68oj8OY6IEuddW+zc7k/kms00EmaJQziqa6hsT5JxFs2FGdYqf2vrkyZDAE2ju7e+1EpbW17+
KdhU3Nwmi2jDCTbr2qX16RiXnNuGmEbtggSQENe5qty3RrcP2BkRdhrbLDBVAb7afZ1F1noGMPQ/
xRQCfMHLHWw1sV/i3eHM4uIV+y9hjXSPRmS1WpiFRNFAb0qOWAfsPHzeaBZ4a5NXwnBHQUsosY9S
HdP54KL4J6g+Nq/1gF3feQwVKTIa6YHvQwA4TD2hxoXa4UB6ehj0Nw8mTOYPVIkR0tb7MPNu/VGE
UAAN+8RuS5gFIgEd3rRk9wncEAi2mznRqovZAh8J7hw40NBzUz5HyD9XtA+MK4dISh4sD+w0Tiyt
bxPSZ6P4ndf+iN1RxvDXut0U/E1jyd9+0tBUxhsvtcZ6QB9DvoVO5sdQfyDp5HG6qPfxp5yTKYZ5
yfyOgbnM2ndded2sVVeltPlBpt9nlCfJvhGOzY1bnq5SlTcql2no6y2C0mZuZ+lh7HvEXppr5Nf1
T6+53r+lxIW+E7JTwnEAPCPB2RPng0k+j685NaH/BXUU/UFjDdKw1v78tix9BSguumv12egOyc9+
h9sLCqSjN1GzXoXy1nkSwByYvTwcfEPqX1b3Zdxwz/790EPlt/asFWX9KBHdQKF4mkUv4y8xtERf
jTBhR7PEoYEx82SKKEVxmbL0T2/1rbhvRWJ97z/J2IFqxpXwdHvxj6sjL5iwNuVtAX+0Rz76z+pm
Ts7l+fnphB+h+CwR54c3WhSV8sSUQpo0eRfaNi7Ub/usA9SclDrvWOsP7K9R/62D5AdYORlmNsw/
JTK+9Y+9fpKxhgV+G7bqSAdC/tmnGNYFQdXwC1vZiKilk43L1SwohteZtBuCksfUqTe1dmn/FS2Y
OLbi+kKsrqoGpjSoRG+Gd37B+SGc0zkvsYjCV8GpNGx1xUoEXoPtxuMwEkRiJ4ohw2yEMY6KewLD
ufNHfb6Arphsug8L3Ki09MJ6miYqiUp4u2cydTBoN0LNfEGItSsNS9ATrnCyA9z8BRsYzqt0EDAz
bMDDx9j9lJMC0L+8s9bOerYcE0NWrDGO23XjFl7zXpNE4TBiBZ5YYtGimOeAUAikusJCEM71uLw2
2ZSrhjzfySEQL9dwr+SK6ETJHBGqbKn1C/AgQsDsKDNyjPxIJeUWn39OWOfrrVzWwAGV04taSLDO
8+WCYhMy2jRgcPJkBy68LhVuB0uQy5nIS7/an3ACNxoQnhAvvtTvD4kgXE4WTxtWdKMuOmzIezxj
KU9d6ZYVGnjWiJtmYO4MzL95Jh3RUKO2ujubeqaFJExIMFo0ZADvJArP0V3FMJ3u3cbOGCAXuSsy
M30lTEvrnCHPnmlsWKB3nDjtArNDee0b5WYvKi2IsiXgGOSrRSvpUmieOVAx2tafP393nxRdFIrP
er4H9399zgDpPu2I+8X03ADRDY6F0K8y9SuupbRw30lRDmSZq8B2cps2hcj8kvdrn5kq9buTqfQJ
p6dz379MOhg72IhGdnIjslvudm1wXOEE7oTqETpmjFEPlADmJj/b1jZ4WBRV/PK4m43PUj/pzzjn
vnlzkaFE+BFt9R4PQ7Fg5XqeohNnSl4SAvmSB5XVqODqun6VfDxubnS49dvn5D/Ozh2x1JKeq465
2mr/iZLdtNQGr5mTB4M4WZEWKMVzDoerhHXf0QWp0ZWYsBALnvtX1iuu+KaBm5BE6b7Rlrl6K0bH
kXLTeC6Q2bQcZfWuWRo6XAm1h6NL/mllAc8L2eesq0lnmp8Jw45UER3T7h3hsOKGR6hET5e/SHtY
xLKP6dOXjUUdJDz/NqS8UN4BBlmYFTYpLOp0oiOTLl0mI9NjGKO9nNYoJJhgd0/V82NLwUIGIsiA
BNkQFSNX8z4teDBwRjupOxRur055p542m9pfhc6qf4/3wvGkl1bgw+7rDZywblp0j8EwJ2LQtZH+
SIVej7TQAVBEWrfWIxLDAhMHDoIDhzjwp9/YhfMt2bUajEqMn/9vB9qmEO4GX/1GjkVwHwZbEGTD
Tn0EBxwHlsNibajGMA8TI4aw/un3kF5ZqzlpELkvKvWicmGBImhzDDk/jL0YDvEWKCgMeo/UNbxW
x4ThQoSXQNYdJxrBsoiaThrNrTF6iRWSZ2diLHVDHj0fuKAfRfl8BO+cGERZQ/QaRH2PC2VVC/hN
cuYwbmFSAe9GO3QWNGoWTAV6h0LpBhZHpsOz97gbay+dzbyRw6itnQO0ryBLypSjQ5RXKeWJK0Ho
dOuUtDmb3VNLPU7BuO1U42TQrd8xOYu3l0/figd/4S4HLIvus391QB74wztnhly78t1WgncsYLuq
q3VfbMAkucxMgJ0muG30H5vjwWIDjZ56N3u+H38N6dDVbQQ2QNej2P63KuLGvFd7CiVlMhlWINW8
Of+nO2YAkTh+36DkVquSB67eC1266I3nP7QKntax4TtJj8VVxxbRBwbrQdMV4dGlo6byDyAq7Swe
I2TjYDWYPgdapKxgnZg8LifDrsc0nAHqcAjaQxaWvWfnY2uh51sjrsJiriLzNZZxv6TEKwu5IXu9
aZ5r9wv9VFlkiXN8uJSb66b2Uo8Ca8161Y1+ljtMixMB8tUpueLrfB7YKXpN+NQdXhWLdPxkm5Nm
p6Gh91uiCL7u1LfYMQ9pC8wDgxdvZ2WnW05k18qxdRLKHkoIIZmDhtcnMrv5hd1xQGgUB/+fUfMn
+VambTQVv91aRlJJ8nQUR+BnGeTrUhF5edFjpcoh8I3vAw6ySFq/J4jurmp1XiXZmv0KlBRyxzTJ
pxTBy8vaoxlda5LdCKD/hNxP+WwLYiZKvGYkHaZQX5mea+0ay/HS++T7YWfYGH21+VaiFgxhPlbc
kNJALJKd3DB+9CcvRSECrA1Oq/RDR9sBbO4xp9yy35he6aagRZN617n8S/shmKhtktJXl2z8e6Hz
kzGvuizZ0LCkzGfmf94Mypf6EAIVvokb/NsaWi6dbz4FLl64vqN42EBh8615bqtUJFqmSlFJ8ljj
vXctc0XVFnca7gJfD4wLa27BT0SrdI58H0Sd9rfYSG3bCOFP+Nn3CwvQsd7kTmujANFkEOoh1+Ut
oQlH2mvlLI4/Rk94kipbVyVt8sfG2vPXRxQVA+kpqIJxhRh3wCl8MoKIcepPxvSwVUMNOrFSnyTc
YiSGZKWFgzHzwNaYYiEBfdUGWey96JM0j0Z/D5FZFdadGTlz3PPl3mWUylQplstPwQaH58gBas95
pmHiuWWwtFodJFpugYtLNJ4WMlX6NCpnHKsE3pMucQboh30y9kJybtfYpcy3wHAyDuPgy/ZnkuNe
JdiHY62ujUgciy275xeZ0DfPeiHT2ng2GGA3rjJLe3BiysBI7kjgccPjxoE5TsPu9tWjgziajJhV
VAoL2g543KtLQ3M1fE6HnQarrMgRrcYLclee2Ss+8aP/pZSMlzIUjOJuahvre45PkfweHpKIq9FH
1hY6CIp4xfkYjiP490jJA/iEowEkVAel9NuNgJQGEOSz5qnck/D6/xIxdh4N1Mz/vzacxNmmuhaF
W8ec2tNoMm/5esUkRK6fd7lmPnyA06isQHw69guW/c0QhChuDIJhHfzddJJZXN2PqbMoMLUwSlHI
0LvDcT3OH4jO+7b2eeXOfPbT4ue3acBO2w4Kq9rAOTJIvD3L3Pt0+a2Edw8QJo7aB/2YHpwMUnz1
tzNqg1Vj9zgd5SPkxLfjE2Vxrt8v2QZjfNjDfhPnvr0TRpJreMjRe8I/+5wf/mZL7aX9HAoXcEi3
Z9nlIy+UHE6FT7GkTGNZCwf8/fT413smO94JigUuODjfuHTEWb6ySnS6ss9pVSEHe2g7zXyb00eW
lqJ3VFxQ47LBpFg7go022dezZuXXNqNgYlZHiw6M8Ce94oRy1rcPTZC56LtVz2LSqH2meOLr07s3
i7PxmUPUKxYwecKm+4IyFCydm0dk6dysHyacqOeIaoGU5r/o/VeAntUp6f0LnlpH92Nj6fTgd7zG
caRtX1u7rO039Aw6U7Xsp/opddjWyHpz+ujyhoiRieG9pe/qbZZEUFakL4PXArQMZE68MfI4Hzbb
qmxF1TtaYw89RqAkpkck3g+mIcDvFRpSYLaUxeTjj4qrJ8lVT4iAzbyxI2e6QLiOmfVFGe5WaYkC
1h3daR6/dQbkhpgL6ZhYasf/HlCrBL4SQew1/zX57r748E64b7r776niVIkfWcMi0/Wz7MlSwgnl
UehFQbOKUuHyBcR1vEQ0ZM61QuBfxJSfvK2pi+BBPK71AgxH/V+ot72PMVDgCqf5CY1/uu1Wid6Q
dOkP+GrzB4duwN69PV9do42+/ktcytXEYFktMUejTGrbGuXfh8gWwQeyzRbtbpQeMhdKbgYaHcnU
vqlZGTr7hP5NsknpKgq6Da4CsCJq5a8G6CnyjubHAlEmVbD+6MZcCBRYTMrVa98U/9m1kov7OILU
2gnnyFOrL+0/emn3D2PFIS14eU3nsSHSMUklGlsbylTkBkhkYoD16paQQ8lQl8uz+OvOkB2Yh/FH
02zYpwuGaTW/8dylHNiDy12u3gJtSJe81mkgOZwPfsgC6Aad+vuYVIePepO0sBvUkaiIp/ERohKc
XFEG2nOQdm53BOjp1NHXt/erjzsLx+jdz6Wy6c4hn+Ld9TJa3nVrhqaApr2x5fipudhkplPOdzq8
8nDYTnWNEiGFeP9iRo8YK9a+lfmv29HhVxErpJegc6p8jD0mgKQWrDnhAxIUlE11JdVdLftHnExG
iVvwsh8P+DQG2A+efgNYhtdMeIpQoFvU1I6nruFCq4f1GKP3NxA8JI1EZzmDG2J6dVpN0TbDPbvU
BtZEUBzkoi6xJsHg/1vPWu29km2Aov99iwiHiqOi8pNpg+AGZiCmZz69BsvTgZkmTdCnUqys10sa
dV7PAs4msSTfx7Q2PUc1xbk1ADzIUTllMGv8BMTnmb/+4UYBE2K8YE8hCzIkt8JzidwvzGyN6b1Y
Df9B48wzEcjtElDCF+SPFfEQcIG41Y0uKB+XMnP3bIV7wNM9KPNmhVfo3lKu2vE2BpjcsplkktFC
/Ad+vf2mid0a/kJhvdSKAXtY6Yh59ZvXvf1L4VqgmbtPmKuVChyy4naQqmDFPQnVmETh7GHsBLlU
YvEXTiGJF3RPKPE2XxLJy5iyZdYgrhiBsvtg6Gue8HfJqa5z9UQtXFQ+Jm1617Ka72CH1GEdT2sW
3uChHqfI2sZ5Ax4ZP0hJ2nJN5Yp7jzJ8bZ6nrFeE3SeyE70QsKULYL74YCXMBjafQK/Iy99vjGe6
K2eB2rZn8pSH/WgIfuU/pa7dzS3IH+SoY89Xot7cLKCakKOnhETDrrxelUUR+Isj+vljPaQR+DWp
ojFhBa86hrNxi6LvAm0UZj9LrCTV9yxRxilR5N9Ql8gTRiTvEKEawGCszewnSKJ0NfnPRySU81Mt
sv5ehDL2aObxG1Az90AwVoj6GEIW+z2bbXAYexXw2dIXv7D/gWN2ccQhF96trvaiVa68MDRTyWL3
gu2Pg+qmKH3+MSLI2J1FP1jeZpPrxqNs+9m/ibpPsTpYgNVWQcu0Vr8/4n8Oue87CtufN5BNOzcB
zUfbcBeZ66WY4A/yBwbzHt2BoETCCGtZRU4zxgW001d71ChV+kjM9c4HkMvzb/6b6y5+omM5+8gK
Y05/4vX4dYPQ3nMp/y0AvNZgpkcHdq5THi/gV6xA9wXadHv5uh31bn+oZHLwO0BG164smEXhSuuH
88ddRZs6b6TcRH0wV8IVrgI0g1Bmy+qUGJ2Au99mbAniXrXg+Ia/oa0g/Py9RD0madEQeP5HvAVQ
41WaGXF3g2wJmj6705bnGTEPk0xX1UiyWXwp0udmGEKs6YX6tyUCXqKs2wB4OsHXiUshe4SkkpMy
p2j3alQOthx73NWrjL6mka+jH+nzboUZceq3hLenvWsIYMrG66bJMPttNpsrLr6EZ+snsRSgk9vR
Yd4dWZc7Oa1ZzhPVrC/4WyUY6L+omOt22aYProQKWtFcsIShDsufQ8kbeyWzfyV9gqr/ZO8/wSck
C9Jh2LBDafG7Oz6EmBmS9GR0O2HhPxsE3fch3v4z8B2ZGjrXPJhOCQa/zjHOHoxAcrKmwHyP8pF/
gY4ytEfZZwTSDJuJ7DDIcWIp8xA/uVr0qOZrIm4Rpyl01guOWpEybLB9z7RLjLl2vT44PNFRB/Xy
IFpvN6EGVvWSBrfj4fGcHWMkNi1NSl24Q/f2k0jHC6lYRpVFAvPR1zwlvOJKo1Uo1/Rcm6/7BU/z
bqlvEzgt+skzJ/HjCuKdo7PgCWqepn9zjQHNmv+6JxhsExQtmanr9SJzDf/uG+naORA8517QrAYc
ycxdDvtLAuvGMLm4zyT9YHVUy+dsN0YZMEOnLKzT0bmKwPqwPB6uIjuF+au8LrnTFr0rYhwesDIF
+DO1TxxzMEP1Sn54mjh6PDlFPuveEl0J82kIwmVMeqfI99lO744R1sM71wGutDlIQx6nuEX1i3Iy
E5niTDmn5nv0FNOt4XXIv7lh7gLyA8u5UonJ2RNiuy8mZL256LMN4O512DSBnSZ/wC1TEJ5N4Qva
bg053NeXWSH1SHmyG4YejLTqk5imF+MOfHLvz/aa9hf+IheB1x0vhmj7D94RFTxDqg8/1USyusQS
O4I7Z2yBKny21CgrCrYXUywSja1NjfKyxfjnYaVWVKwlvSTn79PiG/DPefkkArTbcz6sju95UBLq
HjX44M8gyZNeeeiCbs0cy7gVYhcd4QJRQr77dhXbnuKkQxB2B/vRQu49xHMXlcklBvqXNUZnqn51
CNqaGDOJQiv/B49abaGqpTTu6fZB5PAcYr+hnlvw5hWdnv7JD87MF+cwORHNmgU+LA+dEtBYmIJf
eBGA459Yy0WW3HPnQvFvp6DApHbCwdglwn6lEuY0wZ0gvrRR6FBvnuzHHmawj5plvoHwFKg1WQaI
4BRj2Pneqdm11eum78qMzp5r4F8yAgBId3NJ8jxFAe+l6S6FDTbWckMF5UilxNIoRmYM4wNSMN1p
mrjXFU2f4M4oSOEWAE+prtaJury1N9Jm36eNPz0UGdpWYNA/iBRZenOCvGY5Y4Zf4ZpM1U3ZHh48
xlbHGjfiMnfxnpN7mogIvd0pE7W5Qga95oc03xbNiI7LEJyOsRIy3O0m/as6ES4WKcGT8irA6hzY
LnLy87ezhHY+1Nq+RsEMBtPwAk+3s7LQMq/V5KPooFHYgfBYCV1n/qVGW/raxeOoLPEPXvoHedKU
YR6wrxk8RsPzjHPtc2e7WgSVMzK1FntfEsUH815NPkNJoi/3cPIX7POtetkQ0KwtmUV3Ji9/1/oB
FHITfwmyavJO2hTcbTl93EREysdSiUdHEihMLbiuU95YVeqqD9Cg+lwHnhLmW+7tVlfupgVvN7SH
gIKjNs7d95kM3Uy+nmLC/osdINZ6AOybNUWtUk8FHIjHauYvLuTbiORjr0Jc3vgjYqtK+DOOmsnJ
oSXO/LeV2a3qYdYsUCEpXwr3IMWX0nhPMnGAiYa67oMpGY4X4YNlWU/dCUSjG+aQUpLoIf7827Ul
rxwut1Nxmv7sFnj8FkdCzC7epHlCrLZBAOVOFuL2Np5/HpPVyvbyrVUF9LCs1k3EPqbfdHh4BHb8
C9hMN/EPKeN9erZNljTO8ydPeB9eA5TjfdEfLazfibTG+ly5mx86vhBq88jZYeKPQOBPkY9Vq7Dp
3IrGo4zwaSMO2XH+gRxXr+LwtG+NO1Yterlf4FTbfhtppnpf6bkQI3nwfOyW4nb8TQA4f4Po7/J4
2V/jE+FsIOlK9APw1E9e+Vvuu9kB31Kgvw8aS8su+HL4vRN9JMvY67yxbD23PYNeMDBRJgHXbuke
VwTS7nRCKbrXN3Pn0BSmL5pkRvEfn/VokXmlRASP9tkptPpuF9sXAYziPuf62Y+oGIgr8gJWUy3s
I0U355tcNl/us+h3pMEvC3xrlr4Gc00bUaq0tjn6ZP3R0FTpr+n1oYnOYZOUs222KQi2WaDTsxs2
wn9MHzKWSU21kHolZ00fSXBB2Iy2I70/tS9i+Jun6BeK5+6v6OiI5RxNgZ1+XoElOzZteRk/vTo+
gHHeuAMwKeJfAoOoZ35zJ3aVngur+5BYMkGyzsiHpIgXGnp4RYdeF7dliMgidvjwiFKQ8SkI5YNC
lXX/dozQ88TGA7B+G6/jRpQxC1OunC+fOJ6S2uU8rMEXzb8L8nN4HJ/xs4bYY90bRkPCiZPE7yLb
3xTTg90wM+vuwUCuvBhSJHqFfUAyYuL7aRO4Cb8jT4m3d5U7jFYeZgcdpWClQhg/58bixYBX34Dk
sWX7fa29kVBVjpgeLGFsIEByFFyP1f7pbxRM7IUaoKXrpVe1OgHqgQQQs/G6ykBpSBczb51rkBLb
ZlVS16N3fLD7nKFUaUupMwtJfG5poI9rspBYzBA15eeA+rmBMNzJoMxNTaeNNTVKHeYn8suehRmw
BJVxmXceeDurMEKpRk3KRvq15gjFND+ooPLX28ybx43I/FJJUC1rhFussDcqvpGSBflrp7XwCVBu
294TwXB+y0JPs24ojEnC7WGanPZ5ktzwl1zidBClZ941ieUHJt4xZAWAFnFiBKKNo5LTLjuOhBBC
cTTpxzaqXumyEqthTsL9AWZhf+OgrJYSzUW9b2HD9Zq2xZLGJutsiUshu1Sfsi8ycGfZQefxsjaX
yyRF+R33pd0ud7NWmvtevBiM8XsWxe/ZGfo5RwfNpqXuelae43rk/wC5pKEEF6i1HfvI5PFocegM
DFmq8EI5BkpVwClAc6e8xXakRxaPpUU7T5YBr1Gv0TOi+9xJc3Oc+JrVf4CL/BFGSajFcEQBs6OA
SPH3VrHJGBwpkFoeGx8rej99/VMWHu5HrZfCdP9nvwsfS1jFf578nsWGPMvlf338yVQQNy0PTCRk
i5eN/gLgklYADDSCCXF0O9gCFtU3xb37Ba44783RII+AN6qZ+r/C5fWukw7PG3vz0TuFI5uP3fPL
uZTek+LXXHre/ZCgthgzYp/9IOW11lHImOJeyp/gAD2hH/FsVGBhJb95/isOf0+dUWOOBOK4g2yd
5DqS5flquNc9lbXSdiUZkf0GK75h/qYlSMsKho6eg/IuNhl3TSdhbqb4vV8mkekRJsuaaK2nA95m
dK6seabbPKIb85ALTBZGXtoLsppXkORsZLbF/exkQuVJnJSnTpM/aNDHXkniuDCqFt0wN2X5RTL9
foCXM/k0gPKgHz/xu4gne7upJJh9gbmPOSQz9oFBitVctBUXcZ2+Q2q3SBjFOtN9+wfzxp5tjnDZ
/glO6sMVoYZ7aA9AtGIaIlC5yRzkOcyif6dFUJq3SuF8b4Mi9axOzk/pn6G+KGx41kypKwtFNFP1
0usCv8PgXoGOqivYeMixwLIANdzRMmBbulDgiHn+XfzVtHD7hJd37tVISlN2tPS/2RbEifRvMc5j
6pELqUW8Iyrc7uMDipR1FdUKhMdFpTtZYrkK9QN33zqYXCn8g2nJWHX199NfaQe30Y211P4neXVz
MkhwfdwGKOcqlBtc23x1CFBlGtxc63MQT5I9Qp58n4vHfsKzAvkkBrD7pqCzN8BTRPWnCpekhbhD
Apx7eoJE7VSzZlT2PdIkzCdghYqReuMhV0XvTwMwnkZrWv9M6mejlay1nlCcpxkjyFxJKX3BZ6+g
ZM1fRYpXWTf4VB39Y67M6jM9ahQN92DKZr9xud4h0VU+FwakCorTv1d+oTpAo1xRc6a8gS4oYccD
yQkyxWa3HMf/88wFc1Zj97XzLv5dCxrOH6MywmQTYmHV5gDVhRW0dKew6xqqOYzD+N4SyyCWeyZz
HAT9TQ+z7jxXzh2NyGVHTvqaGQlhffpQQ33f/H/TtMvoFZKGQPl6QcGVlPlPJ1Ir9NSZ3RQancBt
AFdEwe4XbcSLp6By98qVoU7ETY3zaXs6qo3HH8ZL1xUGsAjg2f0phWmSeSlo4colDSnxyGvx9NH4
2aod6JSnFd31LJTohfjXXWuh95num5nQJoWHkUfe0BkFz4iux6YqI4h4XYtshKonCCfaOXiG2p8L
qWWJii0coQHBoSsgwuw4qnBNXe4qb6H+J6+IqqzLNb3u7ouCOH2M/1lu/l2lb4kfvsz/Xn1OoR4B
FWlL0YmvFvdbeKaUtn1EOIBTfEDGQVciuANjoxY0SoeRsWXa2q4KkkidlWaTfOGmbQagSDAgv5X+
Do59raMeZvrmQKGPpctYCUFdX7iqeOYwpvwvR/JkDM17oyhS6gVtM6gdtEWEmFY+P7AtYh7LIdK9
B5hhcthVwZLSrgIF1tP7uQ5nzEkUOCg1thk3ph9Nt5i6r87F69G8Q3Iw0pP0YL2HQf/KAvOwZzmg
BdaCD8wQ/EUEjhr8Chj/FBwS577jOrBOE877uS2PF1EBVKbeTAVpbcGCFdJP+nSQfuCFOV48AW6y
CkMr8MBra3J6XHrAAOiOJ4yyVIL+v1SekORp9xYPRhqRI5OPmRgdF4P1uJc3JVziMF9otpO8WLO7
fMXCakU5dRTzNu9S+GJChr16OCAI1J4hinnT5TDiEVHK2gdXkCcobj4hpJgopWKPTW3EOuKWxrUQ
jIOCZXtyum8DSbSsBqCgnhLsNbZHsQxpwGjcvrGUZOWaN2e2dvmmhG2A8YmZX1s/1lyH1O85jfA0
PZA5nCwgqTwZW3THWgveZE2YyrDVhv+xwlecA7lFNB24RZr8ciIjAB4sS4B+3UzECgUr/Pq5gI6k
1+LnJPZe+NHEaOecyoGrF5exBxcT2mJUcbn46iAheFfBkEMTvKFB/fm59IbkJ6LcCD/1Cas5tCp9
NehVi6QeLfyQzzKT+K6srjtwJIo9xje/ZzYAD2ERdUd4g6IWKQCnVdqi4QdvnT+IlzHtsA8b/KIl
VUeHhDlHn+G5Ot0O0SCzrQL7KPzhW/LstV/AUqz9QVftxL1eF+ojseU1m96EDmxCwgKARdMJulPA
stSukJclPkbNUeiuna0DEYnz2n1GVB2tPSHgTr3SRRuvY5Xqu2MW/5BB1DNEUPu6c8zL3n8Zy+Rp
P56bKGOSXdk0QWU4Ip7+KGA1eFdgoo/lr57R9Us/3+fvFmjuq7dW4MddllPp7SFfS8aFEmuYgPB9
ieZhpBWRMW34mgcKUaTgm/maR1KA0/9Wul+NFuZURB7FlORmLMQvW+2hYrbD+RXsQ9myhIWVlVF7
/WgmhPb+ErJUA9tbB2MTUZWK/1afy16+4s7Q+9ksZhmb7JpRw5I1xpvV14OyVmYLwLQMitpE1L4P
JT6IApeOSvM7T3nSrPAgJhTFdWr3bQe4e0dICnpshMCynHwVnsvpMXqfbHbGrS8v1VJjDT+5vsSq
7cgCRIzV75aAbwgRInfsLmxypJsplToBGNgFwGUbE7dUoFKPY4zw0W0G33u5OFELrYtNxOlanxjF
gI14Quvg3+lGEto99navkck2EuXGl3UQLEFHoiahduq2HBIM8CMzU0Kvtsxl5JLGFCA9wcph+5Ok
msVziY0+xC/0+RzQNl8qzoU2H3a20xPBL6EhCRM0EU3HfE5SP9nQSYL9wJQaOSoRsEuCYMmZVS6J
Qj63RhLntlDG9zX+uvZQQ8by+YD6knKmktftqbFa31u0T4zHeU1PlN0Qsslk34F5iSOdqyQI5zhq
lCugF8Mk/4i6y8+TJ/RYYLdQBLZpnA6QwKUiY0loCaiYtCennQcrV4tt0R+jG52dyVuNO7Z43Rfr
XSxA4scuke/srup4XsqiHkbqBFkMwROFg8d2Hc3kkLU222OgGjbLLbu9JlIHrUA+dyyRDh9GXdwf
++FYQfYxsvRU4a/M+Uyn6ixBs4AKRlS+psaWx3HNvNOyl79DKRlasXjWGkL6R7wPZq6CaDEwMFts
f67t3fsm31XT0ERI6JuKOUpUU20aFwdEax+GHGAhC5niXfVkxBbRSnN8P8io3KKScj+irst4yB8V
SDBEiD4os/l9nvmkU1gwuxPC/cFk+vo3xs2JHy2wY2BfQqoX9N/SMTARoV81PDaLEuEaMtIqq/zo
f5+AOsu/GDBe0xBvw5A0D0iJLMioFlzOeGLum5QMGRSciOMrsao9lh5o/ZQ4V8yBL2C6Sv8dPi6X
zjR53XHgjQf7bY9+lVLG1GD2gcZ3cTDmHAgHXuPbyGUGawU2GTjOCUQCWiCUaBPRrVw9y53ykTv3
9DACwEBKtGJr/WjpKNHra1BE9nPJ+rwJOm1bz4/IybQJVOCcpAirdasDNdJ9GEgGVE0GCQ+kIv6/
OCNYugDXSLfCycKaZHH+/ole+WsP2GMjDQXOt+CKL9eCEsrRqGjZCBxKTlUsXtROMPYSVUw4qr+o
s6KpzGLunbWZVy2UfFBCmPgY3+fq5on9ErOf6jRV01Ho33kWMIQ/tKF4tchflq61KGSBXfnRuG4A
xCgFJ5gJ9B827In5a5VEegO2abreFtXaSIsbZsp8BEWsj7/1Hy6dyeg7JD9CpQSX23nYCMTitSJq
niXnuJnCQViL5IK2mndgPs4rNAmfe1hxzuXEPFpcOvS9c3+4nzGkLIev3MF9km9IVEp3cKqPOjBx
6+uwR9rODDsa7U2DiOFu+m9o/kZclcNiGeTL6ocnV/92Jzdqrgv7j76pjWOcaM5tJNOu0L3+M48r
byqATeJa3Nf3mbuP3WSPONIpoKaGfmzqw/aIt1b2ev0ztPAKRlpjwgtuWJAX33t3UCVO9ZCizZXi
umQUPf7l+oJcIRiH6jt5J0rMPjWC/o0j5ANXEUKDVA4x5e3/CdE6Hxonmb3ssFRdF7/gPTHN+bTE
8387+/6fkyes1iK+uJhA7zHI69QkBToClaBFWWH4aPPmjbmmxuDpcs3SiDETX3BaIlgXvshoCOZU
/AlcAX1HitqmhRGSmVaBsWI2Nfi9bVBfiY4tH2RlXrUfoe/3t/VsEc/VqN5vuoD3IzhLeOyFQh3y
Vs9POeM3/huCS6Bo+hA9dAFJGqTICAvHgaJp5/wNOoK/NssG1CPvBAPU5ycfGIeNFrL0awowGcNj
R2qPCDQyi8Q0Qkqz0VbfehqxREA9OBZ4ngxrjU/CpT2b7DIbZe1pz7AZns/akfGKLlZfq3C9hj8w
eUTfmEUCZiVXFihk/sv6TBqKLbARxXfHDB0zWBKkj/rIYx/JJM+H1FJm9doVllSvTLwtOumOiIHl
md16Bml1SVIvP1IiYnj0atHKuL9ApoIfw4lxfO1YPhX+dOJzC/PB3yi61lJ6FmJM+ZkPp4l70YOK
Y6EWwY0vRExPy7G8fZYp7g+smUbry7MPqwu6i/jOtjeB3nVYSWRAi+Y/uHZZl6NEB+tzbnu3Z2KM
URABAWvtSk41U4CvcRzVfv5nRE4PNzA9wzjc5EdOwWGlvjIlHM1rByfQCXcK8a2xSYiYjfHiZwYx
xXM7IlGvyYAF2PHboI2PQ3Eun48M2cCbAtQ++ub3igDVtCYqWIMEfWVJZGKVHEIo2e4jMnC5HlMz
maXcge42fSZ9wWolgjsmPDUfdRA8Y6InNJaDIFbnmDMwfRNm7yVZZwFewpeFOyy/MAMp0OI7srP1
VDqr6VYWLWcx6Pe4YDmKt3hs33LvZ9f6NRuFeRi1vSzeQA0imr85qfjQd20c16G+Ca++FPD5LN9p
S7ToVZCdkkaxWEUAVK9og/IZuQWokPsUjID/zXn/QmLE/vvAUwndon4FpWcE+YMq1bpsxVdK/UUg
HZaY+nujV8JfxtQuNAEAwwULTSNgxptGkdM3RtkQrFlv/r701DO3IRDi7N9mbmSDc4BsFN5owvu7
CLp01+Qk+SQQN4gx1rkTbI8xLmgxQ/ZO3sRzXf8XrtBRwySXiceE5YQxK456tGr/RMnvdlr18duq
lFIvzuzyzaLxHlkfGJOv5Gc2JBwSNKC1/Mfzj2dMBEb9WVXN/R9O0kY2r3dSSJF1wXXl1bJQn2YG
abIDTH8hMyCW7+rJTmxDFxOAtRElCTZlDkRUpXf/ivdkpUnwi3q9hJ+V2JCOLkK6M+2ddqSt5thm
nOkN8UCS2P3YQacPwCYLzxmXjW8cr+TJNqOZUKPGLrrLMF99Ke2kjliQ3wrFF4+aQ72enLQ2I12K
16JLwzMMGnc/sueAV5dcim2x64dolPCz3KCcKBL6elWhGZgq0B2bcR6/la42M16SIhUDj9o5ZFt1
jLkF9pFzl92kIrqG1OLBhvopQAnbJzZLxddFRmyg7Fvsegzma5AUOuq8nQRb3uiXN7sh5kcSgTMJ
VSCH4f8HQMA/tD0F2FXwUZw7duhc6QgR9UPyY76MDjL6TMRjKPSl3OZvcA9Aky/NQu+k3pELM1oZ
1PzuTM6c48S0WbgvrOS9WNp7XNTxIrjVQ7i2RgMf7YWgfVJTwcCkXGIqtWmmTICV73FEgry2K8em
PscAdFjIxFEV3O7Wwzr/burENV4i79ZpgOP3Eet7aQ6na8D1pvTYmuqHMDQ8/hKYKwKc+rWWJ7uX
d70XKopwtKU6uXWJbV+vVmWtGsDZa4N3HGdmCJB7aXORk8Xm5GxRsNs7CxFKeyV8D4NMefk9F893
rNSUZiVwJG6bLGWunTUDOL/LUOTPmd5S/g1dcZ+6x2CGoop379WL2r1VjsqaAPvtTO2m83iqfLGk
0+GhlTZoQVzFBrKJrUaCDxUGQXr2Su8WOIm4dAlybt2FERkoHJ3z6LExv/QjfCR8ARtCXtg+c0ER
8V4nJizcHkhQvqeRMJRElRHPHMNEypPinPPLSBuRd86tFcHMpzwoerQDkrYpMev8nbYN/UVUmwOv
skuFbPuwof5XZobgMQuxKDiUTOcIX1SzhCrJE+j5Pt/EY3HCbxatFY9J73+xcL7Y9thJt78DKIlW
FHeBA3sXzrkEaCe0CXYucHYmkfMwMP4dn+VylEtBiSSoZzaLhGVFFuhYa8j7a5/bB2iX4ClM3yWH
ChMa0DPbxB1SNV4Baus11K77fTeiXPgMabqshJrebqzmAgT2yGBFmNdIjIVAoqAchhRx2HDn68V5
VC5NtJWmdC7A6ApqZWNhia2lSDPuFgVJYHt8DjmpfjZ/XGD6uXrH/PnupIxHwASDRVkq+6Yr/wjB
SpcsWDBZ1ptMMp2QoPBKc87bg1GfCrcqi6jRj8uAMjXmS32HZ9h/ExLhZacatN8wZ/ngHZi+/Btu
byzppf470zYR6reLJ0cWTFFgMKKKRrneMEMj+bOAp7rl9lei36hTLJ0pPyAFBBKUh4UNS6F6QpeA
S2jv43enhSiAtHjD+qV2i/gdOGD1H4RofkRaY2HG4aNvObPFimAEFw30WOWO1eDhA+sFjbOE8vvr
Vp75Oicx4s/YNxwBECRO9W0gESxbQ1D2mYa1EvyTLpvNQ+12dEpMkKNcEFtdH7acV4Vi+I26IjWU
q9a3rhl5gdXt8u/Ykw4kXgy17BhhUJ6aO+2DLjYVFoguCz2UC9/Ld/Omf60jJ4pAOpWNRH0PKO5G
gGk6d+X25OsAH+66YJ3FPjvvijJmhnpRQRuQEUmS0P8MyMPhxuXsXjY+8GKeAuBqMRXs3GLiI9Ym
GPHQSbNQc7jvlqIJnkcIhTzuXbzA9R2q8VeJiwwODkA9xSIal/2fklYWuPWHQtVnmg164uOlWKxK
+U1z60WoK28uW83LfpDxyUtT4AO4IgkdylrFpD0CPQWGQVGqHJpugUB4TbUsQuagFQw9g/XLe/vl
s/7JyAYzJvuO0jjuaIzkxuyNT1wgxydb5XEJlHsZXI6jBfK09fAuNU+4CPo3eO6rfDjekw8XOAU3
E7jk3r3OZbmqujGrQLf792s+xPqTVISlXi9OlEHr70/hwsKSp34/2at811Cr0VhIANWm+AloU7TT
pkQILw80acwDH2nLlpg1q4jBM2wP8xri+P3LCyMsmwF7kfg4SjfIpqjym0++SeDR+5RUbD32qn7G
pw0M5Q1GnIdNCIAzv4/Sq2H0v/aM8a1lmRw9GlYOaZYXwX5AscoIGtCWTEVlL68RDUyE4hD9JHua
18Jf9zCJH+xnI91qCrNe3nNJET6qGJEw39uEWGY+TuXYMnl09n4COys+UzQzeDkxspyqDTKkPl5J
3tYafCEbaR4s//AbwaJDr9uGji484L0Neg8fDktm6Xt9LZNq5jfK9lmCk/3Wg++LOlgAt+HlDx1s
5nZ83U+BQzj/RNDLzYUUfzPaU3YzRYeOQ5FeqvBDE7+XbIr1t69uNYoKLb0ZFlZD6AmLUGHQhn4m
a4ubFPm2u80G0KwdijUYptRs8lnkPlCPRs4ayeE2onpI/AJTmW8fsmbrjzX8K+G/ZzV/pZxnsMRg
CTCGKoGxJvw+Ol2w+YEQlRd1yL/yLFh9u3b6AHncZIF/znAAhWV0qCBsA0gF+fHmMevrjS1k4qqt
p8ueSM2cM8i5qD3Y7kVp/TCy7PqlnCVNcYxpId2HTq2GLCgGSTZ6ZW1xdCYB/DgXrqKuxMfF0E9a
lzoWyaNiOLq6sckcc3+Na4aF8vn1A/aVtEz1XcaUuKmDlchnxUuuU/DpfifuhriD1hs20PiEQ61U
h06UtENsP1McTCdhIZ+0pn9/upQeRs9cOgsccG46qFzmesp0KicETW9LjXRM+VRQDpQFuSESa64u
3IfRpsogECjN1AI44X1RZ65GWo/yYwG9fZS5hnHTo6QOHmTdRLbrAVhUnCXNWylcwqt/GK0MfoWl
OT0pRvMp7BAqSTAxtfqLIBLQbcmysY+v0ghdBDtVVRv+hgkgUk6kntAzFskbEwVX2DOhji9NDCWe
rsWGNUA8b05zr2xNG0e5Y0c1pHD82HeegHuf/K/Lru/mHTS3KSG+MDEaBnHmufAUO6nHptKpahHw
TYkwMo6mUnImz54jetys/CASb3HomNpl2/NvV61vm4r+qfLK/koZJwFxUoAnGiDvh+1tzG4xkk20
//1KtBDY/KwaICo9svIp7wUmZNA/6I/RK+JHCpd39KaE1moMQH/Z34hgx9imJwSFsldWidJmUS6W
IqCeSL8amLRs78BJUmagsP6ewMI8vgzzTkpr6ZrF+dt3JwbUTWI7UnfGRWaCvhg+gQcOj1vJdCjz
7qs3w7nayUAbl0uYEtjztkAEm8DqzfGv0pc59yZCiE40W99FrsIXeWoK+WNeiU0O9knjIlUzoQhi
wBmOaI0EQJ2JcHWdeE2mjAF19DUxi5Wdk+R42Pm0KX/vrS8BycrF5L7GNmH9ZIz99JLXcXegcAa9
8Bp1rqYPoBKFHLmGLQIgw+9CCaYtPd47rPoabr4EH725TU4Juj7QU3M/pR8dxUTXS1DNAGjT1RTN
gDwv6ddLh/0eiSVKwCfUtZ8fFy/EuExFCzYGkkAZA18zdJmQ9oQqJmVk7TwveIp5l57wBjryIzA3
yxGHz9KRk59t7qMVtfkyUjEfILQNwXEcNc5oVLgB/wciLA/sX/IW+VBh1iLw+++zbgWGgh2CeyIG
+Ig0Kj6i5iBxHCr5Z/5A4YhZ4A7TrOVmju+ScMEiQ90ZUmEap5bTG5KrpA/LaBp/3nCxfUqLvWDo
Nghbgh07iOEFh+j54z//l1T/GjlgU+49//pbsLV5EkrkGuRQ7GYyt1n4vJZ/KocfRtO5DGBGMahe
J3l9XhZi9LsqfJ6JbDjSVNVoxY+plmmzkad0on07Qrjf9e+LxQ+WBwrp5hsPERtfkNCbjuHbPSdo
WgW9nEWGo5Oq+bEPWb+0+h44nRNP0l3v31iqxkHLk3rVeQwgSn1fOn1NfJNuxWjDkxppgAukLpzD
0hNarlOHnK6HgHBrbGGO9+toaEKNQxnUMiftzHPipP0hyXLa7nDY7A2EoXF2tqYaxec7zAOI0Oho
hvjZtjhV5plWKNtgRsFbUTnKZla5vgZglBnRK4Va9srp7/3ATnTRNsyWnp365i3Jk4KkJSNUqIUo
cG01KhjYm9RAWZGZZ3t66bPCZeMLTKLc9OkmumwpsH+FgqH4FzvbtxwZ3O1swyXyYgAjPRy1wRan
LE5elBmic2GjoGJfxRkA73DuFxKA5WLWaiFacAGCpUbc0b9/M/ybLIAJW/XkJB1yL5C29aqkGELo
FguEMeP44EbFcvlFFrowFeepoFTa/tAM9R0PrEBp2glA3ZnUZJAJJMlSHj8fh55U5LGQQbx1fvLS
tm7+sevwV/8eaSkJ3igwZ3v1YunWGu1RagERDtibYHfb7Gt1bE2Yh0jt687ATrvXy9Hifnv0StXV
gUje+mZ+nuV/KzpidBVbsqcXU/xQimpKa+YkoIUxiSTYGyToKcdozVD1KgYmYXBLhnDGDs7jd0VJ
Db3OBO0jhFn+mXDk3d7Zir4U46wqG5NqleRYcIwlqzoCnQdGIHwV35B1/KD+wP1pTrhhMFhm2Ajt
WUeQXsmkPBc8UaMosMMf+LJWKWVEWtzTw+EcfiHPF+vXwBmQcfH9KGHM2kinCcsmHzWgNUeo27K0
ATMPVzONV9pX1T7CFm/Sz2hwII8EzG4vgrSlMs9tGt4r9NnCI1ZxuNXW0J0t93Wp7pVbspRbZkT0
0hV64LveQtSQYk953NtJ31nRKzvi7gOzlTLvN+3ara9OsQBD0/0ugETNR/uAYaSa48fBUGyLLz6d
wsV9b1tylRMp914qgiVfTegbMtquUoVKpD0rkTJbnNL2maesN5Gqt3TPpXL8Vf1nYWE+vzzDzrlX
nmWZo+ICuKsjzDrkGKksweN1rgabhYOEMG5m81rjBOr3QuP3J+w4hCZbOhc088DzjoXXM/45narz
VFat+4v+06vvnVY8UJwTkQwvHUcx/9Ir6QwQ/DGZ+UmFqfp0LgLgkfpeHydblDuLxtPhFdi8ZpPT
Jn3NID+SeegRUL9Qhxko3hiJLEBCs14ReQhWI0+mwTRHkuMxyCh2vruJmaywiLMwxUHyoI7hhjGW
7akKg1jox/iwB3cVO0RGTX4cLvLqqM4F0znwu6rWsP8kIESjMyCJAmDUcAXZfw5uEsV/saB7W+VL
yPO1GoO8dzOVNRNQrw3zr7A66W8IL8LkAdiFk6xcwUSPDo0cGP1ZQvakmg+Hk4zcZS2zcZaQfVAZ
JFsMNnvphF3WR9iBGUG1xCdTb2kI8yxd2+P/gFNRsFKd0K1PdQYKJ6N/TAWB+guI14bROCNApwck
3dLib7+mjrLIR59+RtyTXlErTiJtCaL1bIwWJtI2DJNjSh0IDy1djkDW2tLTHCZQrDgzrhyQdyKA
37UjA8hMHiHPmmnxfcg6A2bFGLvlvZz22UhT1HHDCkFmyXS/CijijEL87QaUnQjfz1iUSXtf6tM+
/sc4oyzydfB/0IwSKD3c4sS8B4RHvBQSCMeavgVPM6VbgUOzU9qke0ljqZ+WGVuPv2q9CD4chBoc
KNEeOJH250cZuGwgaMQZUUwfS1I2F7njaxK1dcZixNKVBXHg1XYMf+dokyVYukm3rhgAadB3f30x
HBopyiGYWfEbIwOS89Kp/EETw+wLsUs4T0JH527D61hAFOtPwDrZT0P2TUDtRErXvB/cBEHMMGH2
YOoAfnMmJ6mmJguQLyO+PrdMvFiZNBMmR1lJ+NEUW7MTFpE6uCCHARs55w2gdt2AfhCZoOcXLwLx
/JFRRI+2zKdU67GMFqOnLYzXYQ3WiI5VUj3Kvygi0n0OZobRGW5DvrQfz460XLuDDCWGb9yZyDm5
vI1C28VWSTT+15G6SHvoygQAgJChqpVZ0gaf+JGITTiHwvvaRup+In0T9EXTnRFJU12XuHwyHE+b
ILZANbl8STc3UrYOPDNqxUB0t4neCdZ6ir4codG7ygVh/luYfBWlFVIL95JHpHcse9cGH8TQGJpU
Paf/c4lSpQYmWvdeTNGXUFE2FE1qagiGnSO+XCS3RsUwknvPdggVqMzQ47x4qpn7PfJcnGQikxVs
qBSRuQl1GmHeNGmK6k0EiNAS5Q/AVblgvq8sC6xzTK13UcVxHSAtXMIOfZisrswukXjWWX5h8y5r
HT9PwUHJia4WBzHTg953oF1G1i9+e0Dpr5B1u1S4Epfik+BIMDj20HSjdL0rTEnz6MxfhRlXncMP
eZtWytIu40J43g3ANaFmWmvkmigvwOaVlley/ouWnhFXB0UjRjGMmwQxWXZMPkSQdFzWYQqH71Uq
tIxFRwz401SnjM19nLcMP1lSQlPTr8i2jIPtIlTz3tYGy7GXAQu037RbaDUOSUfS/etqof8zsuQ6
8CefHOoOuv1ULXTVCbTgmm37pHxjdYmgBxx2WkTqiHX1I7gQGmeuVltqcJdeeXPZxIakgY3SKTT7
DN//BL9GxI7cxCi9yJcMrpu1AGJjo6fnFT9PmrBfOIHI0BbPQRwertMm7qw27T+nNNMOmXEE+ss6
E1Fjz/9Z4AeaDB6zPRCxF0uslv1xvSmm9nzKxn37+KgonE+IhMqkxJW1tiNCN48S3LIDVAHtyzFH
ETf25ui+CVkVyOOvn4AbouB6w7kV1ojSC7+dquEcDOzIs8VF5UBbP/RTU1uS2ROvETvT2AQLP3/L
y+jPBcKkS0CB6MiJv1DsIcQyz8y+ftWxc7UGXkqLSSTIKdjQrMZgda1r92qAFVtxa7noywuYXNkV
cXJMtAcMsvWLa75F4jstsow6PdzVFVuTKLPpM7/E0/ow1FhfyYOjk2YbL3LzQoaBBEffN5XvuAys
kmud5z0j/M8tVzkjhJv4zV1vWI5lQuSS098Zp8U5KwRlqN92qEEiu3aiDddJz4g+ynQcIn7kz4yE
RRImtEZAXlPy+02lAWVwj0+oNpiBAHQ9x4T7ywZKMeGi9BytbRz9XHP9X5cYS7UrR+419lFFaZBA
D+pmKFdDSPYGfGggsIksBaBwLN3PotNIWO6YrrS8/BQIPPAwtfirT9icoPqGWvCo+AffbGI3OtqJ
lXSWF7RrE/bhF8FnN1/OgjZtcRCcHnjy+8Bkgp2Pc0qpZgkUWmTQgh4Z4RAOgnugeZ58TYy+jmTM
gdVbvMWWoQFyrc4sCW6xR8EAm3OaMbjeHqTutMim+gcRgvbwaXPnlC+mWQVsUggLpCzjSPwl3VHT
SnIkI/ujSzcOwOYJUXRlV9juMD2EMupJV50jhbX9iDa74Wj1Us0k9kPRCYG94JwnjSc3DHEajaG8
QIktYfLmRsij8sPNE53MbbSwS62XoHEfvXb8HktjFzMTjutQsbhuBORHAg+bwSsC2pCqMhriYf09
pA6MMOnacCRvK708cgrDqf4RjEyfN8m+jIYxMV+aAOKEvltQdf/cwp6CrLFWBtEx0krpi4jqdgYQ
uJ9o+U/pUTVAJxpFPnDtMI72iNNbPI9dm25G2aZZQ7umCwUYT+QRokWi+T1E2fqs3znvjYoHdgI3
b2ckt6qCzjFUiCM9AJN8L6xLjnvgzKsDeQrDNXanyVFmTNe2yaievTqNMcZliLIulVbmXIZxG+r3
t0XponOY+LK0xxTQO3RB9p432UyQVfDDk80bn9TfGTnVuwcyJmA90oQkLapJ8/QrppBjUDYL4CD4
wjM9kAMoVH5bqF8BrpTdjJU7uCYnKwmOCdAi9sV5vgEcvldFqfQMMm5Q4oW30fSH+42ytYy/4GOH
IowLUaNHh9tL3r0K8SknThTQXe1qiCmsh5/c/IEziE4bduDTfnaKMXLmgC17Vx95aDaAmz5bpUTf
RouXDDKm8Ko+Zi2zspeXUQenu76gflUlye5KTq9NyfLRMEFwbxsrkjcZwLJXxfuVjXlbH2pfLeP0
3nY2aqqjAo3+mkUYLIJSSjERl02aRX/A8DODRg/9VmoUA6cDAPgrrHPoWC6cilK1MiFqldPNZBlZ
Kf2wqTZVlVIR1x/qoTHJvjCdlfg1T6qCCBR3l1JpDxz2j5qKdT1PGkDvwshUid8XvO61hYBcviIt
ZR3qHh5NTvY8og0PvIENP4LkvnBRh57wmFQ1jR0xCtHI8h/QrHV+uiN9Igrf0zlApJMTBaDBD2lc
HA6ii7SqIGcbNG0OjTZ6LUyxxhEM2jgN1c6VIS78tzAsmbUffp7eoepoQf+RSVP/RP2gOmjiszSv
jWLxdgj2FtJ5D3W5BxdimOk62sLwq5hj0SGnWD9qJRYaPa/1m6pI5knEone2D0ciJoYHZ2ydp20H
rzW8drTQGj0IfZaUGC2qkmNCK8SYnoVIarOWtNYVsqDpKtEDZTCBvF7bInf3Vczebmbewi2inNYA
Som2GE8LViyme8jEjijco/RTZNpyrD21BL9myf2dKIcqrAWRy5WO0ZTV5wZkEQAoUuiV2VWffIJc
l0R/si9z5IH8mmPyJQJf9/B+k5Nj6sVTp+pG9gdwrBMCbNFM67px6tgVHn1SkdL7a9Xa9a5VgEOP
NQYG1u9gXqTmFH2ItrtCwT3Dtk25avBSMn8SpG9D2yu57+VfyMi6WuJ1GGKl7w0MnOsAy55uWlJL
Sby6UUE8hb9TK+2tcm9Rbw2TBzph2M5yquCpTHx21rLGPKxBSCPO6UOkUdxbdZSbw5YLwBm0mNt0
kIVx77IR+ywGHERl7FB/hzoFe54BubJ7lJL6fZdoZldrKbW50lUADGNgTS4auiA4xOoICWh+s1+k
zrEnXIw2GPiCfA7xA8LWQ1zURkYtDITO0/Y8pZNZMubKKhCmEk8eCh4AauMKc9L2GbLb3jhentt0
e/lguxrjGT5dN9ddXEiBlO54WW/vyiufMNDcyyHzPgJOIoWsSyXG+A020CI9f/TJJ2AOUgUYw4UF
flkmvoYpw59hVe2EVGCl1r56riE4EKS0GD3PdxxUJPbFEi6WWUyx6SEPZC3lGHsYYXlZS0rtqMmZ
HDTWIZkiwaaZjLDANXb6lM0Vac2AOQMDfMjaiX1hhNDPef63HDUin6icu5t6uDZHQHB9AKejC1ff
t51t81n8Ipg4QhEnvfzA02vnGgrOlwYCc6UvqzxNZfm0Bu+AmSEQIR32BEHKX+huSOyBopq4yKSP
4d0sFtAJBjSs6qntXD4PyZVQrNR6Gb9/bfU7/HqXFbhfVDDNKA+eJyeajWxSnbPt3lUdyIvv2HNr
DNwXFF9Q16f7CZvFKtaqNSaDibHRW4KFA0CtRmwnAXkQKsVeE0ZLHd38T4Yh0gl9AiegBjAvgzim
T88X7dcHhtVHc4gLUmTn7LsXSAis8GO7pljMt/a6pukvnd2zToo8vDm1dIZNQOIKAYHWCgMa8M5E
DZg+oaAfi2SxG5XMwSZVN0tG3oNDmvWAXfMHIDJ1i0eq1tUUMbdVgDjruHSdAfvaSDKZ+t57yv45
rwPw0vo6AS42b8SYZswendmIHY3RC7c9q/k0bln6oshSqPODqQejFZkwYR3C2iF60jpea3CFc1Yj
Yu2SF4iQseuXq3e84KuX8MOBM1kRi3jhEmRAFJlFxJQpooQxPXucp8YL+t8ZEl0sGNOj2Ux+pBve
KPJBeEGPNVN+TJRsj4/nAwnP8O7wXsI2i+YELpi0fQhceTG8PBhWKCiIDM6pe+2VnLD9rm8kLSCA
GZ9fEbvORAZ3xsyegMXDK0eA7fq5PJD1wHqxUNvCy2ozOTnZg30f+hI7PSIsJ9Dt54UzA9upziEJ
ebcp5qJ5teugc46Z8R5WyTpMNdGis7S0DQYdGHf61Sbi5CIExvFug52bP3D2uYFk3FSyo2ehV2ZO
R7CyDbu581mVP/gqNu4OX9FH7Yiv4hnW+EB0doHbCKmGKTFCU/wLfoIHuiaogMpdRx39y92Xnm3M
oJioVdKJ1twQDqeJLI7+U33PyxzBOA6UIHrZ/2BS9io+DckTa10C/L9PolAYxnHANvKHOetcaAtq
pd9jayWMLVwP/ao4T3OGWT5Mnd2k19ztNlmRDYX41QZt3vD0lEIJ2UqTP59kcc+ZUWeVNIF0hLOr
MGdV8Z7u6BRoN1s1qp1PrSJYM1mJdZ26xb8tTghFqLu82mhwzhYL7N6StMgyBvGoCKMz1CgHF4Sy
9ngdNXfHqu8n9GeU63tJMW0d/QaiqjCdWTdc2q/cr9nwtWP3UmeNy6UzQN+RUqXo0JE+ivBzQcrn
croglB4qztIjgldqphlugb2qz9472B9t03jTogGzw9BK4mT9248WG9TdElbgPngCn7WR4/FBgGf9
lEvxPuIiJjFXj9pSCumfCylHRqVTl6WGjvRZu8pAi6DQ43eRnkEG+1QMXiKBje6xzltcFWO/GyEM
OFGGb05YwU6DUZd7B91IafPHnzd+ojI268nH9eDEO43WyDPHH3W6Ylbk+Co9NejmOmuKY2dAOw4T
MGjm9P+c7j2HvAiEXgZiQsTlHsGyv1i5QjZ+sp/On5aw+YgTtlyqA2da4QHJzRWQHvcSIHkVwEog
IDezNi25gcY8AIcuuG+M+slDoKVmcnIaNl/jXK3JUXD2P47eEg/rRwXlWWfvl5Y63hlKp5tSVWve
GyKfeXRKMe3FSCk6hwRnX+0cMOJbvNupkW65+PyPs51hMvTk4epkJy1P3OQJhZOjebZm0TZ48Y7J
7CTTQU/u3MoxmDwy63Lw+5qMBqBfI2cfIQalPYYa2kWZM3Apq2rIIAGA3qJIBbqZVUtwZ0kqyGaQ
K9AiL6Ip3PAkJ2af4SeHqYSarJ+EMDI32vYX1QmmYR3FGCoJA/Bl8itLI13whBvFP29G0KMnWiBq
KjE3rQOlfxkbXU38QQ6DdCor+ig5EdULQslVfz2KbV+QqwNPyF6WROKGLhuDtcI5nLlzcc4DkLd7
6ZBYkCv1tqDnIu2WjnNTjxYINK3HaXK2vizI+jWJTJLG1GnXmyrA04KtJSGNe9Ix8nUao/lTx/15
Pl7Of6yvHILTkxv6k3zX73XkOwhw9dJAY1WYGajSWshQLxYXQDwCQnq/ZHQA2sCPYxNbcDN71dwS
nRKdYMqxUiqxmZ9cpqcdEJ4IbNRhl79eAs2KDy10lj/hjGo7LzOp0qW7482NI415gNRBIOcR4aN8
xE0jLW4IXfOadlpIuE2j3LK8K5F4fQ30COqFBvrwP1V0ET4Ch8jwDQceEo6peqjfSNMs5kZ2Sjba
hvl8SyYVdKTx6qjKLo/rUNed06bWovZSEjRv7erfCQgD2n7mf0Rw2CqdYoDYZR8cbUTMiN5rIz3s
/Vre8mAvesCwX/eJIe3CR59zqjJw7jS7W8jWrek9/lstjhTmYuc+ZDAGu/1pvpYZAWDyhPF7wP2G
zMUD8UKZ+n/MVYCLi7wTlfw+P7Anqi5BLOanIgT+bBOabbHtHeNUsHzn+LL7RtDQuo8J3P5ee1P2
Y3emT700OhdNu/PQzsguAUiTB6+6t5w9M3qQTJSDlFP1zKrWTjvoY4RkPR9LOVG1rGyJzSMHUx3S
O7II1Foc5/cHnuufZiXTdQt23vwJ+N6ns//yViGFMFL3H5srwGz6f5SPaF9ncCLlnvBx7WLd2jpi
6abyu9z0VEkP6R/yElNzXdc1OgwCxhwfHv9eiP48arpcUCJ9+a+kUfjLds25Xr3mpsEGd3sr5NhE
jLYKGPHOwqfnFAr8E0VDQThNbDUbp8//x+JdDGtg3/W3bjd6lSlopXkEYl6W3N9OrolGiEM34ep0
oZt7cKAZ4mclcwehb9yGl8oO1YtRlKSLfaVOjhpocpBZe9jHIuWE62orQxMyIzRXQc6v6HRTCp9O
cTDXcpyuUe43guoTQuO4FMR6AlJHtnOg/39CT9Cn1FaZdsMCShKrKdvfsQPUPKjjZeLgH3lXbUUx
t5MQqT6ok3aH9yqt8VxdcwHPZtBbm1aO6hJfemcDKmpuCAeBdlmasi6R9LzNIGNgSUi5/wuMlPEK
agy6jULA9Roruike6BQ9N1JGwdEcGD9gSaFXrz2OYmf4o7soVbfMWb3W8EyXHv7ipZIQuqPb2KNJ
t/ZQ/fO9VaKqrB+S8gyVgq9Md5FfBurCalvfWFxTUvSV7wh60w+VX731N3TN+4g8AQf/s5ZauYMU
R5yui3QD4ikaI+6nwmkHrQU9+IDRb75KpUYDvmqTGFemB3DQzb8+xTXPG6Z0dEV0k1KweH2d2r9L
poJTumPRv6ExOgQAZ/NQduzKM5+sdbVb3zfKyeopEUYHaXDGqV18IWVbxc/VLCM5YwhbmETDCToD
eXgKAgdRT28fKQqWHEmVBpYevPYmdrbNZ36fBDo7W+zeSTvTVPr6lXK+z46Af7u4PwbBQzIsAcnd
iGIFU7o/6vM2vHV8bfIMp7fyCOse/7HoHcz/N8MYhMArxH/fXEscUtLpm87MPS3ZHyDydNbMMOLI
881yK5QDE/cuayjH8rOIn2ixCPAsXpulQZNxJ/U/BLO7tPE0AwdLHaLxEpGoaynE2EDeTdSTbxiq
9no6vIGrc0vuPv3r4FkAWsEyC8x4CB38SldGp/tc0Tl/Yo14Rjfqo35hjERlBSEx+0eoN64MDJeL
p5dmSq7yKKETYCaXRON4bM8jsDeTHshsNpeD1WrQjyBt4c6zcoHCp5HSRFhV/EzUCkzuCoiozgng
NlwvEgj4yh1zQ3u0jSK1kGF6JWyFCpQ9azSa6eQYvOnMn/P/W38u5CCe66PKTSHQe0ewVlOq4uvc
hbUkmgSxPbrEvV23XmcHEZ7z6oIZEsD2nTc8TKUFCMIn3vJqaaKnmpPeqTf/anSaaj30dQUQ3IB1
/Z3pG3pMU0qL/prbOyVEJI6GshU0IlS2/qOGI7Q1YeUJN9KUeQ+JgrumilXFgBZDV2TsqzVs7HTz
J9E0P4f6PnGx/fKWk0S+7WzHybrwdq5JE7CCwgpqW6/Uhi0v1KBeFKSm0watYYjSZFvTjU7aLiJJ
XzMCf0FDVc0oINOHSp1BN2l0xeWpBQxmdLgLVLTrjK87cujiWbW9xaaqvqSvR7xzN8YTBLWi+FY/
7pYkp7QYu1tuzLjqn4lQkktUBIBlZ1JMlt2WzlHzR3zA+P1igclxPUvQNkn6zshNdw//mqhMXGDF
LC/GvEglQINVeOu1VZSPe/paMr0qb+5DICIpXWS3/TACQHSnfqfY/4St5QrdDBfVxR8PJH6uHdK1
6oiy7Kq6sRTyvwNcpWrfCUrl81zMkh0yB3XmNqZLwgJFRAPy9QUilhHTlASoLHdl9x1Cxn2/IvWD
EqGF0EDn5azXAq4ISt18NkJ0scacemBzJoVxupDdXsmAiNotQ6v7b9M6LlSrOeZYY5CNMxNgqGec
K0FGLaBJosmu25FXlFJ9EpZpBCmydDqd9CF08QRvzxX/Ph+l4iDwmge6SJKKypTTRBkqf/xHs36m
d3ikYdeU6OKmSn0apDYt/AIJiEgCP/fNsH/XYP2us7HDx6IpeDDqlI8E2JnV1nJEjCeUPTXsxSjd
zObdU4qbRmhCnCm+n6Jw4iOLvBuriuMUL2MMjXRRbrDw0L2/VI5kM3wdJJSkZUSdaxyR0rNqIg/A
mXpMugmK3XRwG682qqx8gj84iXN2Pr8B0aSwTjVRqgfSEgWybQ0MjVjgaB2dpQeyYkSz7yTTLh2X
WmW5+H2CzQaPU9H0qWW12KVRFVXlYPHQyh6fg3hhY3xwbPq4sTTRT5Si36+BYgH36shFUDycFk4G
QWUHhOZaZqlYD/R4qL4E4u4wBLJsNM8VvTOScZb6TmezTcWBg1w91g0Vqq3eryCIjLRrfhIEX6bR
aFhiMBwyXcDH1Z7qNxJL7q6i2YxODq2QpPP1HTE29yvP9+aXXBg1vV+f/K/D7R89DtNtoow/2YbB
yYizZASOkfZn+aovMhM7KwNNctMABML67GBbvZM8d7Hlmfj75elkw0FZkp2f5xhnKAvPwEfvGb9p
QaO4zIEqRVApakuGGSD25YLuLHB1E8/KR4rd5k21DhmrutKTnldNeg5Y8vDd9NZrWfaS+j6yaHgd
901HHwkrYOS8B/k85jEyqo8mJagFi0F374KOwxnaLhQJUIP4APJqAkGF9Ijk9Ld0viZ2JaryrS2c
j/+Xtmn5m8NFM8rTqgm4fOAK2VG62cFfWqBm1OAsmw58O3LxqU1tFyG652Kp30fWlLGd4sEFnHXr
fXmh1Wc2aEEmm4jHXxFMcOU9Yhn+ApA0t5M2ILYCf4v16ACgvvLoS4CI45rafxaW5ZSXTr1zjyEr
lpgP9SI8tPfPB/diNL4dYC6BeCZzgj48rhx91hgrCrpPVAQB7MNBMYmZPL5TvIrNFunEBF3vxVUl
GUqy5SNex/bAIhL/AJFCzT1A8CJUwfxrTRLo6iEuIRGA9N6flY2IbL7/fXcMqE3oWPurAEn34WdI
mz5kEbT9OTH4m902vPGkurXeKZC7biGBFyr87/0R5vusi4onek859kLWTpYC+4ZhbGTYKhOZmY4v
EUqXKnn4hBWgVTp+o4nCb+tiEfZFUgy2E+z0QnrhYHAVRgAt536kq4rP6o4FvFtGQVx8BSsZiE/5
0djcqmF7lQQtTrRnRV8xlHdZ+FWkZypSc2G5Ol6O/aeffLbAU3u+kW/mnZFRh4IkiZt3B/EFKed6
yH02RqPrf9m36H+1abRANCt8qeu0CksFT/B1A5/OqVzREgY4Bcd6m2oLN1pjgc2Ldq9GSb8nZnSu
rqSp6R941rKDDAgX0RNwU0CjWQa/lXB4F9DlJqcREV2/LjdPhSaCrOzJTNph8XKpOrJZQilQaMh+
6y2n2uBNzp9d5m/1WkR+otOKYyWYB2VgE3GYv4l8njl8VmxHjUG+8XXkrkCPUVeDqc1uzUO5uVZa
SUMT71L7xDUwZIw1ERyxZdckj0FAFEOOSBXg+03eBFmxMSyT9fa26GYAhHpMBkXTBqh69pC3gzkV
7JaHFPQ9PQPjgBipOjPyyQf8hU88cCIt43lebrV39wBgRdoE03hnt4omtq5AHhQkijXB8D1PKL3V
zzZFbuWtop61jLLRrhY6jqj7Ym2q1D2QOpOAYKtg3e0/NDW83Q0/L8k2dh6UiHyYj7Au0tqiB2OT
nC6iWYmN9ZhS9mc5c72wcfM3jdfdlqOL+lZf+RPIy4nqtHNvc9xRXNfEm+t0wpyP7UcTyIjrnNwi
emox4d5bp3u5cLW1d9ijoleYoZr15eXNFNgWDVwqzzMKIcogfYd4PmbEtGil3WLs7hcx4KPZUilJ
kUZWaSJg7Ciysux/TclYz7QoKg0Za2ovuvVRN6mlabjCsBmmym8X4Ej48972uiMGPh5B5ffo9lPI
m9Fwa56mXOoPdKkkz/irwYNA0VnWWBSMLUAtim2K/SGZNRpHMBaJAT13Yta4bCvgjcn/TPQ8IRgy
MGtT1r5I1ysj6JRFeuYvS40COlKd+C1i8YwpP1n2bsR6DvClGrI5ItFv6I18Bp57f7PSNAOBHkBG
yJVSn0QII3iVRZuL9TydDTLqy/0u0KcqSnxy4RZxu6lus4gSokh8688OGbMaGV5WW4c+ImzyTYcw
rwSzkVU8Serwi59QcsiGDe3kqrdDsKzwyvG48aiPQL0/PsJn6uFj7VbONZKxQYar6FFPuRGXi/rW
L1HsB1O88gCNAeNBFm6NxTOMBJ3CEUVhKywhulSDQAd6aQ1iNrOfT1ZJ+EIQkppAIglIzXu09V0C
afwhGRpCxvkdou7IjtwhqS3554pltb4cvLuEnJkGAvX4kNv9zlTTFOZpKLrk+S+oTeHFINKF4Dj4
rGcJISGNMtSrS4WmSgbytw+KTCjY0ax14DgDWd1YbpeR6Ut90QPujflE8P4bCK8bKn8qz5lcYlAS
hsHPmfPqVO89D+VDT+/M0nNsp1L9lr4eOqFtwoAtZzxG6ZKYkfIJy3krbX2mHJVbNxSGdJYu/J8e
bkZRvekQIk24v1R+YaEYSpdWvyK+hdFnG2PIX3ic7918lD0QrlLXRU5iOxH7zm8XT67peQZT5jBT
x7T9DAFZWjaHmBV5X+IeiXFazq+aj9H0JwckkW53RigwWPFxrsinVYvOMzI/T4/Ri+G0uJ1xV6pf
sMYFLfqv5cL/9s2RQSjY4e8affEFSUrXR4tnF1pFQhLL+7pP1y6xwVD0MN4jIOST6Sv/i9XlbJA8
KTbB+2c3IFN9Uc3nZ+H2kMukQgk2syD6Nk0DgrWU738KOtiIQQQCOy6D2/IT6IeqF6hsFRWuwPnz
47EJlOHnyYw8q9XzVNuxKPB3jtlfnDaoYKFVVpb4j2Xs8xYysG6B3WfYQFQkeo0Vt8R+YdDiwjb4
b/XqKexiziNahe09YS/6EzleQw9HK6Ykx3LsWjD9zrzWgMMWmUzvMaTpII/djR0X5jspfum+K4KU
q2KACJ0H1Tu4s/rkef3ag/2UM1L5VkqTOorVzxgmIkd7LQC32yPaMoG/eRWiI2AEETsYhMN0v5Ic
8SdcV1YOAVrhUcS5bE54Pk+7DfF4CbgS6guedKxiPqOrwsuj+F7/qUwdvjHrkpZQvngy3+Q0a+xM
MR+wAKXnCadrDmS3c6M7WgzHrKSWfeK9IuYcs2NDvTEZGPuyu3vR2yjsDGriRpovU801pbfJTp5A
zN1c8Lc6eGcS1U2w5Qlm4fDKaHGkh78qD2VbEOD51H354KakKYWbmjloabvVNhjS6XC4B7lhTIX+
pD5fxZBOAiO9hLUVng+ReTm4eC/Dao15GOCK4rcFKEVv8r2Ahw8mYTUq/X2aRpEuZXMf/eIp52qS
FlY0jJ7+919i7hcdFe1SsRM/Qpu5RHZx4D9tlwPe01l+o0DoTu8gBQedCKx1j8FGBxtBJx63Av9N
nQftSIVuXCWLKVkpzX5Jba58tGzEnPUJUdNURxxF7ShP7eakny2l6zdNNMEbPffDgyPo+jtA8FRN
DqrQ4lnKk3BOMLNZ5l1XDxfLG2tBDogiJD4xILJCPU6beNq809qtZKe6b7dJDMu7WQz2qQ97Y8QW
tuXiAGW1AiEqZ731wNenesCFWxVN4JCErejbj4xP9ewsd6WSKs3Ulhd3nNJEgXKsIb9D9w6SlpPv
WKVKhr1/PKmkSXTdMUCL2ZN/yzF08lSVclcRqf6sMafZod9W+F2n9xN+X5CnKHy3VnPkQST2b15P
Gvg4ryB8Ae2ouGoZREdQMPAAoFZDsIoYGN1ub6hnr6Wni1d9vVCYTBMl5iWUo5XyqLQEg3mzjJsP
GGX7f3FLH/VbeD0xUt+uL9pakaPtP1J91RHJhdYGmbEIUjvATiyG/2IMLPvqWcaAwz6hJXJTA26Z
GZmh7/8lQqHBRWM+NRCj13uELwEEqSjKfFUP0QcxhKmNcdBay7l33/TSVz3SG7JxKU9V/mE86grY
TkPoS6+stbWVEFgDQOdMfwIXnjG7ZyAxNTwWHNwBgCoOWsdQ5BHPmLryB21gUtdAhImoqssMAW+y
V1sccnpcyZQVX0uOxz/8Gv5wEe8Zg5tra0C6ICAQgEejQHRCpyLQQbU9gS8eFUxNLW/f6I14jUtf
TjyUglKbDyu6mfiOaAFA/8ZmgmBlv68EpcjeXazLMoFhDsK3J8mpAXCuwdCQni0D0LRBgrSxq4l4
lzrlizf+z2XU0KnbZ/zTB6jOFXvfOr+r9B1S6Lk6xTI8VzZv60+C+786HRmkJp5rDTh2UbwDIo5T
BPMNGH8l1QS4Q5GAHnyMyFl2TSBVvkUlxp6bc2PQlOtSR8QwFdVA10PYk18iOfEpx9znMEhn65zr
tzcoW6AY9+u4PPY3/EPnuRjYZ/5VbpppKPrbgQleT/JyHDs+i3AlDIGWXvkKsnmPDJojd4A5//uY
6/lHptdWYxFMV0f+7aF2OG6t+qjsWqtWMBN5GvdXwbN/oPerAbM9TZdOwRaPIq+sJqBGViDByIwI
U+Ig4vVwFaSBcyXBpGv1EVNDHKOpbcBPtbbWw5F+t5JFoQBjTGamVEvvuVcYBXrdMlnEblieCgVS
g5yDhTtCll33Et8w24sN8QvQoRQbCtcVS/OW6h1ESGMPYpNblX5nS9NGmVNTtpNpPugBHTbwQFAn
hQRrdYq3YTZvAdJFy14DcK5MQtvPEQgDvzOVBuiuMg6kBROU0g2FUmlHrnQJIYd4cgSx2Us0jIW5
ksv4Wn64ldcVOSRCs6re/2BCdAzJZvWlBziOzKuDgPsn6NVS0DDgZYdNFc0WJg6LmoOC6z/x8x38
HFOyx6UzyHBzpe5QdhL9wigRKMnJ7SUFaIkhpM/MOderOwyj1VRl7SM0rHIghAbb1lQlcynFaZmu
hNwF2ia2i7NKVOJoxEnDJeadeu3YUms8WXsoMwYUJ7GaXutHmKFra2bW2cf5Pz8jFl2rvptcJ8vQ
23YGnuGu6nBg+J8ucRfQboTumVbzAVPywTVZLOgb8fGWyclgz06w/KrQ0aKZC2RrjBJNnedn1GWd
WYeqiNvr9PqovZrMPwE8slHl6A9UWmdpu8MQ6/dugW3T02SEzHgF8xUWjawJ3o/jCvz3DT789ExI
jkLjS7U5CPGsgJ7U+xLw+Y2rxNWO4rIarIyu9PbV/tcGiCxx5yzT2ZulftmiAkaA5DYgAmo0ZTOu
lJSsXBLFa5E/T/D+Oouh0TkFWDhAuhTTZ0GegS5JjsEz/GrK6Fwe3fhoP5pcFfVZtFjoJrik1l1J
mPo3GzF+2FIk0MczfT6dbGaa9L4n/Kw/AaLxDscC79EPg5F0IE8Df/6lo7+/JPWZswOzvLfpczi3
P3kRJxloiVmp5rjSBPyNWpNle7cVKAEsyqGZmTFB0ukWpRhqhLm9iZCSfojgYKnEfdweImwYgPjU
uQZSooibestsGBsp2kBMoIU78L3wYAO37wmbfg4SERFzgv+ybXUUBfXLJ3UnCkTi5RryC7JsG0sQ
9ZAeLCLIc9vkV0lf+AbpS35hFe54B9yqQipf1Pg1PYExHc8eBimbG31ZFiouTZYx0ujZUDY6/d/R
Dt4GATvozN9KVdPY5ORKufBc3jCeEZnk7U8ITRajJ/rNqXebowfd0vXaXAjOUmcg71LfF/UAhXfC
o90ZcbF79RJ+0dhofBgZC7E6PXnpzH6xjX20L6t9zAEu4ahCKp4d8hM3JkDrI78s7dZsLnp+1bQF
3Rsqa3aYl32A+rjHY816LXkQPUl2PHpr8uKPI8ncNciwk9bR4Ok4QSU05tceONJEtzclIB9+gSpE
qjLqd1dBnjSEbObj0YDty0iS4qbS/VF9fE+D1UEKzL80D0P8FmcuYCP0sbvPnkGgfFavfqeQarsS
oldDR2edcGBbNYeSZiZpLoU/514ZFloKe+Qbh6v3a1U3ZW4PsOMXNVDVVK80wHObyaDJ8NQvXxUx
UmH6fOoV3vMU2X8EZBQK0Uvhf3N2LIAQ/sgVbP0mQdJSTtTk67/AY30dqIbxQggHxLI8ZoQA0Ras
egKyQkIf+WXt0PlRUZQstf0j57GYuW3qD6cY4Bk7KXntosM1awz+pS5m4E4/rZdOt6r7nLV38/LN
xARyjZygWWBoxD/kbEcFJ0kH0dGhnE600P8mRmxx48GxShUG9KzbKL6MIaP0KgFVQlGfdTwCfF5d
9X9lmfDO+eG/4Gph4XIMmzqCe6SHxIh/3LkLdAgfWaR79UAZiQhjNdaO+0yZx0b06vYz7g6gJOwi
a5DcNUDhO+Dw+djr92m0EtK8Yfi34n2bkQJtbR5/EPj3q0VcaXsUOfkal62KNjOInYVlGhBr27mv
OrqzevF1N+4VyI3dDX2/vJ1lM7yhdZXJDkGTJ1T4kJDV/gd6tNwJWCxwDVViXr0xXHhSBjUc/o0I
HEeYwvJjE9Qk/xmObD2KGJXpXfbkXgtupBX97csfeB6NNCsSD+RtO3wbZSZv73HhjLxYh01ChI+f
5pQJFCXXrekPv5G2YN2H0zXY0eeHl3PdcWzgWJZRwhkrfdqWbz5NUH4H11+ssA5XDLRvg3eWXnyF
sHPIrMcjmJyea5Gy+RqEHazihufQJksNwwgwXrX0VdFp0EVrcgyBdQaSNT0UFVb852M8wKk1nbN3
P7h+h+bGNq7kwdsV7I/gSRalrnoWbdtM61uXwZdz3ke3WMbmaVT0l0xjYHOOuiidBzm6WRrjIkyi
al4fVXqt5JrCpOJZz1/PjaCR+lAPK9APdW/YRJ9GNwex/b6FTWCB4pvyCZNK5jarvHy/U1+5GInF
ruvwZwl+Bdlwl4eYaRDvgnyyCc2gpl9YZbTqov1nob15RpKKLVIvrkwWu2Cg1Rb12xgDcpe+vWph
lqxAqhI3/aA1w+F+HuuOKoSLrgguQn1QfzpiwAeb6tun2lYq/IW5kCZZaligcNW9PzmYqYWpuYgX
yIe1FqHEfYBwNLHNF4YpK4Daq3czabVATTgWMyzRIgJ1BWYAc47bOF8LD+afe1WHEW3XJ4ibNVij
yw+wKe29IvcYlXOrWhHXSFUWqEIN1oPdd5rtkefogy4dkgQt2vOi1XRDnTvGEe/328LKKsikwiN1
/0lP2iE5qbR9hwyaK2WI/o1KEQgtUVq3O2ojt8fSXcas9ap1OFGjDPel79zldurm5TRU2Ss+vMrv
dwYo5DPlSdmsCIiZrGeIO7HTzjVvK8KqMsG7U3igPWTj5HRwGAMPnQCFRl67O/xmhLl8TvJwDMEc
qJ2Fdxm1+LKJXhifGHIpJLjTJ9/cCL4EVnduvCQhODhZfPVFoQuOTE5Lc1jZ58L6S0+l8RNRdIVT
1Z4cutbZQPpEf7EWNolKOcgxTwnAvPUTZRz207DEPBSpPQse4n/nU+AemXzF8acqHP/o7d+nBYLw
a9InSlzOhuuPguhOEYhpvHzK+brZbyHJIb/zPu3lekMjiaSL7R1n/k97GuQJc+rPI2phMbJ3xo/c
us1Ks4+8LUBhp5+ha5Fdt9mOuQ1vUq82O+e92F3tV2chbkqOGmVoVq8Z5lPPqEeUVZTJYXrILuP+
hRTCbXSKBVgZInby9N7yOkAihX7AvzAMz2Q2qavJNLuhjGGfAS6j9xyz7JeFW3LydBBzOsIXe1Hi
o6h0DWeNjd+c0/J/d5rgawewafCtSIEyOvzwOOHIUC33ckR5Z5NfEr0QAILg2c73hCcc3b0QZTpK
K0RP5KO/Yx0HgeaaazKNlUdflNJdR52zk8gb0A7YnGhZldUxPEWHQ2topPow1smtZkXYHhB5rFCt
fkTbRdx7k7vb4cxWw+97scyBYL2pDr6saCgfjf51XdLv/+pwESfLbKWbJjrJx3dqblP15bjkeDZN
CJSkBW/AhbGJHJOwb4mDlvMNkNoRFJc6aBQpny4AkBNTNiYdDDXrsB87jTQdRkJKBwFHTv51eh0k
Jbog+VFaBu/nQha6U9QAun2lcjvnePdwMnKAQj4DpoiUPy0HJHRvZx1Wf2aWzubgiacdUzvtXXB9
vSpC7ZeHThg0dP0dQR9Jgo9bp+roy80zpGNcnUV4SpNBfQ6L+jTvXwdF9g0k67ZzstLAETida7L4
lIJ08jqinjhpsrUAGdTtupIlfJBiCXaVa4MqdY+VN+z2AAD9mgpajX+iFqgAJKEtJCEMTA0q0TBx
cX3sM/lNyLXZ+qhqe88MR7NUEb029UsOGimqC6xwRs6vbK3nvMG/HU23svfxGKaUUikXsE2wOFw9
PyZc/mpzUGmiXVyy2MV8ASO1YoJQBfpXyrFbXjJEyWUtXBObXjEP6MRLYmZ5UKcySYYKQW82gPTA
ZLkLjmyu0zX51qwsWOZGj/znm2qJwsINHyoY83JkrSIzodLpuqC6Nx27w7apIsOUty4DNiL+QbZO
eDYi1raTysuMuY6WBJlp97GeoKmJ5ra3OL2ImwEH7Ded2dlc2sh3ZxM8cp/xei/oZ65QY+rG3pW6
SVNwb7BykcbnRvsi2L+gk0gPWP5oDAyQ+yWT9cgMgFgHfBYq9b5ZDRDlM7WiuysivtdnMeIft72P
5LzhXm4fKwmJ0Rf64RShJ60odd5fB2oCNX+6gf07H5MT9s19Dxf+oIZ9oAslBmKH1A4esVGm1gM7
ng/4Le9rKfnhy0AAt9wM3jkSlVrxZWGn/jZuC1s18VUTOiEL/IaUvZCRM0do0MHZURlFO7qA8Ar6
FhlJhE70sRX5vIXujnk+adQQWKQ8GanUYH+MJJDIYfgd0McAXx/zTDSbfPQIadNUWBQvOiNKytUE
6UZSS2rcDj7tzkdeKCtkXln1DPdAD0DokEvWMuZte/cd9TO69U5G+zqMCoCsSkIrhHdC20clg52R
gX0tXKawEmzocOKWjVD1JgXd8CWjSoNLLIoire9U5PoIeiGawzGMXTapda30xE9iBL007sIUHFmB
lrDsZLeRuArJGZuaupZi63PJeTzi3MZDEgVyrhIyPjia724wA3f88BXPDhf51wtdfg0TCh/I4Ig9
LoQpRWI3LkoS1iH/39JV2H9+CBxhwg28KODDFPMiQUO7H1w70ouI1ovv4w12SJbzCg9o04ODiH+s
FQaMH/ezAhrrg/spDDS4C5dcp7qwvQMRCyVKmlL2LZdV6oVPU1hrPAPhroAj92E8Tl66ckePcH3c
TCFj5cn57V88AM3BVC1bqGzPgXN9/y7bh4OwwV6mE55Q95E6a3xakk9l7srp9s0vLHUqpMJWXe92
i4mkoHV/u5lrzxHTtfKC6J+NB12luPQCtrnHamDCbk6CwYug5AUXilONeOZ8+EY7wLEorf4TTNT4
UUOdSegNcLnqEwv355EUejdvvutu66lfNyUkmUQazDIqwj3KVuQB7GDq0+EnJ/bHg//vRHNVTdVO
D4nKcjbj6bZuj2TkLXZj+D07CSiiryo1COxMsja5OzK2OyMLV33OGKM8HLGg6WgYb2I0W6UYKikZ
pwSKhKg9AMYV3DU79DV3UIdKFW1W2/n5I0lD+o3VhdKKuYgDVnerhMEvrrA7FgPgjJzSLkIWny49
TtfAxX6RSwLZ0KzF+DwkkWoQJe5wFsiu3Qh9okfVVRNOg1Yq0oqcoQDniSXlpSHLCsuu+0IS/bSQ
1r/m2tM0DXrAfTtpoaJgWf7ll6gO3njnMuIYIGvplQOo1+MD7jjGjMiwqcPZXkVl3mfw/NmZAA4g
bkyJDOQE4gVT9LFcUOQmfFzwEynzXNxWZ9fHV2hZUpFPnUm0mdDJkgkSmjKj8YYG4tgDLZjW+gJR
Tx14Mnvva/9wE/JmviEw4ZiiYG5sTxL9ONfXjyXddyR416wNvEZuGdBb2lCowPUWITO+ppFUlFQI
JeztKWZzZOUzxqXhCEvfk7OeNf8xLoMOfJ9kFogv3ZdYI1gIBKkQ/+gzZhHwTWBo+orYWGHKJI77
sMrTrcYGkKk+3xiUsHGa/qdAvzq4v63J6673chzJUudhPIcnTmqdo/9WYCR3NkSlV9hTpasV59RJ
mckXpAbba5Gqg7OZs/upImBPMZE9DWuKqxa0d/KH+aZgBEsAvwZ/uYft0aWf8yGgySdfJxocPsy7
64ybLaO6Nl1OjOfr87txEDOPOXX/mij7sH4HLSD4U0lIMzR2E5kSVoZVqz91DF5GROBtWk6XFdCY
gPT34EV1E+/zPkDL9yab9snJFd9Y5DnEhdjZrm2Kq79k+wcT/8nBXL8wyIABmdh+27cdPAO6ofg6
Z1OtkVXlWQ7PgzI52/cewQblLozhus/bP5mS9pmtv4O6gFmZOtFTJR8nk2nAX11lwI41Usf0gQL0
RsBAb0YGr3NCXP8//lXMey9msT/WQgjbmpOkqC/BUTDT3nUfOseHsoJHp9jt0oVXPA9WHCYDS+zD
1IU7d/OItfAgIFeyRrdM0sPe5nfaEJ67EwMln/robcY4Of00hbzSUGzsbfg/+u/+RDkOt5P5xXoA
kc/ecIl5SNgFy2o0jeCU7O+nlhUkwBl8TRrHpX89mETqYVvKV0Q9ixEkfh0X4FQKInCk9ntbSs3e
oLqJjITWMuCu/22xejEvwlNL5UefeDKmLjBeIaNE68nvSf6NZYSdpS9JIXvEW9sNgXpI46iNMRjL
DAUcpqTpLqT/JFfHoO4378eWhxl9dhADRWJZulh5xdOIIHflOJulWvMmhqV2qbU/ihRxB2CauKTx
rV9/Q4UCN9hOSziEzI9mWbwU/8fiMyzVzmf00TGB+NvhIIrz7wfzBbvTJpP6Yeq6MW4keVaWrT5c
iSXK3oWPm/LGD45TR7Coy0DdT9KjxVcw+w3jB8YlcLsy0qNy0BOmdOsCDFKFB97SFO3YYcGnr+eG
u5ammedTPIowGjSLTh5YWarPOAIaLkxXsp/rTLLLdeCVkIzBYluIgNNEKtLk66ysXopipnnX0nkR
2gURv6oP8mypu3EkHK7vpQ6XmBK7It/GkQ9kSyqEQ3clPlllz9Urc7Rmlw1gWcQBIwfO0DegqG5P
jsFaTKV+L3zcsUOJMUeDRl5eE8J/jVLOwzWYa20fvTXDnQSBO+yAaYPUqMppvASYrNm01/qaajez
ujuDW34rf9bRIn5x9CeX/o19CujdvCXtWx8Ar9EY33ql0tCDFlnf/GxICoIp9S+n1AbWeXEd2EY2
/obPHTFdpCBTRYKw256mbQIoQAU/zgx4dv6YBZrCgX1alKWQRwXZ7odw+cv7eyzuJocU7hzFvU6o
HIu/M6hTJJN8LYTBZn0MrVjPmAJmo2jPBEAVDBkrwqrvOCJ3OtVDQFHhLGJULQ0+63U3NBA6FM4z
5UrI+cpR7TRrf39Ef5NajTuNlV7L4Kq2v5WgvCw+/pdlSe5hpQwzyI/Cmp3ROA59v2TQsIP8P3yi
4qH0hls12YGHP401OhfbM1KASv+9Ei1sj8FIg+alPfuQDckHqI62fH388HeLdB2wMvL62Gz9G3ap
M3GoiKYT/yy2RV9run1kt8RWnkZIyK88e4Yrb3/5OKT3ElnD10gqV805qEnEux31Jiz4Jo558cpa
Nya18LhiTH9EWWXLr5qLeHvUcyS9LlH96PGwbcCtAyhEfVvL0q98Q+QqFNoL3Rjvgo8+KUICpYHf
JG/b6gYK4IrlgyrqyEJ2huWdHzY17b2KMZgSURP8K0GVCxoFTWPBKWohNNVimn3N2CqYdWrxECoa
Jin+vQBWdJrF7oGytxXo2ROksxmYCv1ttjkYz9hVYrpbPFYc2GPpPl9K8lhCCM16w4XUBnL8p9F5
oNaHeWV3GWBq5kIDJFjjMhwtLrU1yDqeRhgB9fBljKWtGqBQ40h9ympZvyHha45QWN7WVeKLs5D+
YvsqOFiWRFwmMXkw/sjglM+/YMCXlz8SOSNDbti0FbEBMqSneMDzGiQtOyWkB2QmxeftQrPn/ftd
gbidcNjO7bTN/0WVnWsE2HHXaa7omr0UO1PvQ7ywtcFauGNAHHrwHNpbyAK2sHmD6BOPAlRawyp/
BPexdl0qdYKblg3eQTrygVAsfcNWGq3PzfgXY57I80tsT+0VIhhbHqvAxo3RF8pUIU86CypctdEe
mVAdapTuUc5mVa/GAD9XtY+WzF4ZnJIDZLV2aB+RCAbysqRIHw4q/dXOF4XhhO+c+3o54XXKWhQP
df4l4eSLsv+4XhnV7GJ5pX9udcmxnHIpjv8QBObYE5HuJ8aL6KfELv2ZsRXTF1vxxaFSlJb8u9CZ
OFwk5Lm6mEo5RQctF95x+8NsMGBmEB0lbMzn6CfsD9K2lIamPXU4rrhI3dyJ/diYXdArZkDB8sSo
H/oqR4o4nOR2NjGvHPrHVoVUy9a2iHmJM8AQqwb75e/kbY7f9E/6Z26XRT3AfGheWF8FgtE1WImo
Trw3b4U+gE+MIO5n+DGZdS2FEkkLs3tJVIyoNkdn/5pze9kpPXUJo2UFuYIvbXgMCcFM8fFBwOu3
U8dtLIiHPa1KLqvzunpmBE5SsEraFX/ncdhnrKEYD3rbwnaz8E5D/QNRD1cW1mIDj+nCZF/cS34l
8feLk44WC78KFKDG8IslS6KeyBE5/xB/LclpwOzCJZQESM0cb6u9nakhecy6fHVr9UJyDNp1A/Ip
44zMxEQTbZWqoKo/8azxcvDDSVzXin5VGSEgR/AKvfZywZY50z709ty6QWACu5uRlQjNeckp73A+
kInLchsoBvjpsICkiMFVrXXIPVxch9Rclv5FzcuLOrfka3f89fv5oiHg4tV1J0UFFNY2j9FxHTHg
2i7osIOzZlhPWAn7RLxRChLIN0sIgTIDeDuh5m4hDdzn1+u+tUabNi78iswsKlAxwU+r+jn/cIhn
o2at62K58eOHA3XAZ+egCGAKBd3B6fyGAbySzgaQJc2SRgvze3fP2W0pzECuslyLShySwwmVr9hI
fX+QG3JF5X2yhNDGU1M2u6YCrOv+3Ee18dc/jGdAkqiqsrNjDVuRNQo9aJWOXbZ7HDDrEHGS/1lx
t8LP5dBKQ7tiBjbZzJ4Qeguyg06RjZHYcbAbr7Z/6Ro1SCiYGZdVKHGOgUVOnjONbSDjt965oen/
Noa/WczFmBLHS+/bDtrwYqKdlfc89Nw1j0NI5LaLBI5e9vendC+cPBx7vcgvpCnNdECgL90vtStd
eA14mJhufl2ROhO6/mFbpo0NGr50cWz3VvBkDTkawNDub9pXk5nFX25ZPpCVVK9cC3RqfCl1CEZj
IyD5zPN29U+tiBWPISo5RAWqrUcYOy7wGxJyAHxFQ5AoUo5T2tq+GgW9IjNwVIjCiepUEvm3idv3
vfBPEKPfkLC+OVKWEeBe/SayHZaGlZjbDxsu8z5rF6a9dnYhd7zDgpW7mejcyT84HYra/YCo46c6
YqsToQuFFXlCjPj03kJ1mO/xLPfgY01kGB5Mpk/uTY7IsYJpEO6UYSk1pnWCn5RVlas0MLltF9Ny
7TMEMrUQPUCbDzipkzURCt6/WzL3DrdFvhNq4768rplWV8GyaCmKyhenILfFiV4KbzGnMrHgVDRU
69Pg5B+WgR01XsHCL21uiIOx2CBHJeMggSLx5IkdUMAOBFrYJYLq2daofP5/ejljrlxl14dM7ALU
gz3O2XiIlUsDx9BRLOSelNfCISFv2fQX8VT3Vftikdqu9ZuDqWpbrQovzlKBbDrl6ZN28opdzzKg
d33iEe86lyTJMo+049YtZZcFxxt+1r8j5oVc8MBX+oJC+aK4UkcTArwPs+S05TckldCDpJuQkoIp
f7Se3sL81s/exrFzYbchEBu6rL+lKnJ7eNDrFDFNPCYdX395SYTqKKUYL3X8IAM4a2zEU/Rxb7/W
i8uyB0baeECPuNEdl7VYynbqzXOnrwT54CHyoDk7b/BJMz6XsoheZnJGxoct0PmjB/Nk12QJWDJ1
zoqXv5GEgHXZsvJW8eqKvbmHqS2ewHYAZu4AMtLBsQF/oUQlXmru/2fpoOShbRkqlCF29cI02Y6g
vblN3c7DQfMkxqT4laNkIpBQjvJiXrR/VqFIlUM7vs17PNyEanLuDU0tFiDzmRG1Ec0H0ncKZva/
8j1pA+QxP+ocihb3yHnF+7lgvfeB1p2QD2KAZH8pTicL3PlSutpizhciCMDgVX7+zNMk4Cb3+aDc
fXsMYbUp8GNZi1dQoh578cISNkiFgDY9FRfqvk79kkXjvHOoO5F5ntIys14D2Ukudi0ssdZIE7sV
C1jLGOx1Q989McLBnPjjTjd8P07antakiqB4/t2FcZYDvT6rZxP1CR3sI4jqNEcIaPDVZojV2wWk
XWytPMmKjc7PU29Dwatsc31oatje0lWMwfBLuE5AaFz5nfCD0ZUbHrUKP/ImWZU4x7Y+ccWk2trs
QioYi4Ik0+91uhqiIBqwq+o+M65AvkncUu5ZGhPoEtcMHJCwcVgROdDfNGJNkl9Om5ARvx+SvWtB
tgE5m4bnITb5E7aLyolyhqFQBOVN9qlDUbO7y2vpJXMvDSRg6fhx5c9PUABjUIuwSsGKkh7jmvPG
Oah+2jYw4ufsFXWb7f7A5jQYpCJBEsPDmQe4LK4uYFy3lQLu3zlK5ce2cKpZ6fjlmh5quMgqyEe0
ACNHAREz9kyidoHPQgFzjkh0lrZkezhKIb8oIqVgUjEwjnrtZsVYAtukm8Kid7rBTq6lPZOXjh69
5fRgu6tbD/ohhgGhWmZj305QybuF53jlSUUf+iO144nTi1y4a6e/gRNCe9kpwWtZUM8AVc0SUuS+
fS8YFZVhKVasdlORL3FJcZQGWQ2e40Xe9iL5qxb33vnAdyttKpzJ6MK5ULt9WW//Sb1O57j6GYRi
ldFKqXmWg86IYpwGuS7xlWpfc/OFf6DrdVNDWghr1lBU5Q6PK9H3XTFUjroow+dI6lrfjDuxVcO4
cZZNh/vWvN+uRK2bLHIucM9gD9mHoIedxELv6tfo6US2m8rYc217S4w0jx2XN4y6ZBalN6biGYNQ
ER/mwvnsT61r9HhCN92D/oJ3OGLvbdoO8gI3cEY8DB1BZTjgykeuTpEJ/OIouEvGeJ5vgBXT0GSV
z5kCwpPl+qmFNIKMzwJSUFWqlJosadQEP6PZMByH4024r3QDD82DrFtJzE2G3+jK8xZdiKQ9YZTr
Nrt3d7olLIvF5cjFwIc3/qzFseONgwUiaFqAoML8WvIpqMhQwUY8x5PNdXWaEOPwMXrMRjfcLhQj
WS8GvbXOmbjTY4HLS7nMuxe9rZPrwc997e80dY9leEU5d1TQx43rATGWivq0tQkKsVkDhzLia7St
5LWvfKt27zqeV4OA2lQXiytyIGvzDp4Cpte/QUNA/mhphQy9WDp5F6lyFCvyj54w/eH/bAHDJo4F
DUeOo+EinXI4em1qPoDh9lWQ1xRwOMQfqH7RoiK1gtjw976O1cLojHI3SX/XjHNl3aRlXrTrWDyf
S48WRTbf9kmWwQNF0XRYEjfDbLhssCRRvkb0oMRsGh2QBpFyxG8AzQcrB9HTX9jlWrIZSCFTV/p5
d4BOcztVVzH01xnF5Diw5IQ4xjCXRSN1+csxSK2utUAW7XVuaPK+FQKYh359cSReT7zVt6diW7ds
ugljgvfTCpcHdtjG7H/MHtWaufDPaW7+1hdsUnGTu+AhTgKmuE7/IMwpNKsBURzr9Mp5VD5TeMms
EwPn4ZSk2i08SHq7J6KhzgsacYefsKnfkNh6cVbN6xwQC1y5jrzcA2yswjJAdTVZ0dhWgVDmJqUF
skPfOmXPnrm3ll84g7uKvnoGTmPpZ3Ty2Ml92cmCGeWWn4tUDlPNssy9McdxVvswfqYjoQ3k1j/5
jxiDbYppZOiunhW99N0izFBk2fIgAfFg9mYGh3wNo7ZsisPqolyUt8UHsbUebsOv6NwW0tXbf6L2
dRhEjSGel7kJUK66gr5e55fjxtzeNqL/BnO57oQ9ANlrYwfI3zQvheznAsS7ZCFYVXb7k9BXUSWR
8z3u8spytCbv+AIPdOk9L1nIUEjj5jqMjSzxFLUBdmhwAgxR7albFMJUvm8IxqCVTv5SOmUUATYd
a4v5VXm0W0FBIDaYkSYkB6RXcDMtpEFx09GiNKb/Adb+WbeAYZqT8sSS+IgufplxCkN2W/6s49fP
XIAjR2m1KNR9NFvBC9FEH8rq4obfAR/3+f1eVw2xoYo1u5A6eTNVRUi8gFcsBvzuYMVLc7b9S1U6
HkUQbSG2XmntSMM/34na+u40bk32ckRAtgVk1tX5sL3x7kSkyTeLbTVW8PL00BOJr0MtiliUdvtd
dnRuVUX6yIxhpP1Ri1+t8wrD+fqiAimxMB6gFzjJADnIxq+E3rtFN3xAvywXBqwnGjurMvKCjhYU
WWXMlE6PZAW9Alq794Zh69hFl+pzyux6b7/7Kr+liyezNViGCgPL+72OpnGy2Tpu4VlbYyp0r2Lk
7FJb+wzlmOaUEwZugVoRVEwfF/2CJrfCVIdyHwntZjHZC6w8RBTst5xhyJlGeq1Z6NvbN1Wnu0zV
i9O4KXshfl4aajeT+gpy9SnJv5P8cQ1SdXj0R3MSMriajEymoZxA+kSv1sWOIk/uxIwvOaiit1+Y
CrkCVcbdNRkVfOCk/VDMmNkTSvzXt6kUWLaS3J0Xr4TsD8ePL08wZDJyBT0vmsbVfOt/hpL3qbPC
0mm41t5vfoaenhqg7qH+apLPXACbBWMGG75MsC4gTJB7yNMxTyIms6NL6qn3xgjX6VEyIwpZcrbG
9UpfL+pJn8lQIjGpZ5a9KAEGmYjkPPSckeMgM4fcvL9PY3tc0ya7YzaHsC1FDVUj7hcDblSGz7Gf
4GNs9zrzL26phMlsuYeTiNvnBqXfUMIDzQXn0207ViEDfkxKCUfw8fA62Shh+OXs23vLsL9uM2y7
X4vS0V8QZRK8O974Km+/dSHSAuXaebMzOcj+GeTNzXdQIjYvEkZUVI+pp/vVOrrynKIl0cWZg0w+
D9X53qBvU1XrwKsHq4WslQRs1nqnuLjFI3DgiZPyzv0trod8Mh/BIayi/Gb18EMgVbq5TieKbeJD
WBkgy4DLgvXOYyevXIg3HkqMPDtN5h87FNCSnaOU9c/fCUb3qjWTNra+dnLMeFgNDBRtVQlHcI5B
IjKUVd4tBmaXlkuockLenvEgc28mgpPP6NzO041uPMYFIQwMsD/qqk9sr/3YeScXLQ/5QuFpq4a3
k8JFWJTNOlP8dtsx0+/rLCwKY4FJRAV1qf1rEBAFGgaDZxAYReBX9V08rUd+gMPFnxGj/id/HnbE
ai09ICCiUvxdSZ/FSH8c2rVRv8wjuitTGy98vs5YLL6d+tZEDcmVJ/aNNLmRjxXtN6VKPtrtu1mo
KSNcpryD3Pcjer0VDKT6AOhYp2EEXiLajg3hVwIyiKX4fXf/WQynfipIXk/BGW3icHpB8TQuajlP
VOkwknk5gMMxWkgioM1EmQ15h7RM9A70HNWvxJtuyc1DGuN+xCnE2wYwTF9wHhCzm8RDeH8Mmgs1
58RXa9rvg4ymK7kBTQ/QlTQOrflvJrf04eh+qmbKUI/nX3lJRvlW21++jGyGDLqHVddDv3qPbAMI
wRMHEBVSI+g1BBZkQfBnBoStlbNkJ+sRtjJj4ssZNDG78zcLKnOMPhmNDmYEo6pzLvcHS1jXbmAB
+4TBY6c5GGi3C9jaiDWrKf94nhYzwo6vy9JkJ6Y6EnVYvwguduMzKalBNO/5pyZWVx7LmoAFw2vO
r0EMyplhT5zRziDCC6IBdhRVEekK3jzxJElbQ5c2leKslYg5opsXIuoMyiogGd/RepG1X7AGP8cj
raTuQ+M0m9dih0fzQLJ+yqRw1s/jz6v3lMcbghrJSBTAHm/vZZ6TJkUlT2wvfJ93VzYCjum64mRQ
rU+fqQOSJAB1rjzVjQKYM/MATUwQHi9lpsx85sa1MkW7PL+j1F1vSbM6v7N7IT7JUKLf2HxFjQhs
S+b7LwT/DxaQLbXJ6zBZ8I+aVUuYkfNyuHjjQzvtZKb3wWWn9DvN+nyJUnqK9oBfyyzmJnq/C5uc
ebrFchD+CFIdY2zw4+lKm4adCUi3RoqC4V92s+XmDf+T0iRaMPW+OIIynH2KbABMeiqFBMcX+17O
LOijMt0LIXM81LDKtpk9TI+/b61n6sc+3Zi4DOTQ+8wGNJw7UN8+II5d0H3bS679f4O3Xj5M97Wq
E8dDx0CMWy8mtB4GAgdFBVyENaCseTRPbKUbCSl2Xk842xltoJHJo7ak3wmpcNsy8/SJAlqB/bLw
brP+RQKvK8NHHZa/kj2KP/Eiskw95NC+1xVxWYFYYjc+2ifcngn+NRgbthsVXT33i6ncR6tD3BHV
jweNzZcil2C3TiS2HtsDcx0lnY1orodvlBUIPCMy88M9Q7bUKIt6DgMvPHzCiTToxibLo/SUWC94
pcJixFV0aBKva4F8SlH5x9zr9rb0v/iLNfB9k4LnbRAXu5IPULpZiMLwz5X6D32kexgB+3Hm7OkN
xIUzKPp63bp0Cr6/80LsaN4+EYcWGOw3moG5IWc0bkV/rDDsqO5AxRJGX9CbQGfDqPn2oI10foaO
HV25Lv1osszxZab7S3OS8PpCC71wrJGlt9XeUhTbO5R1OOxXLysQbLAuQOyDiPlVA2zbhQ5Nkz+x
przJHmHaz3CdnJsHD3FC7SFrbV5uNd/SOH/WZCo02otz2a+nZMIoCSDqtyfgfiebHlZsfYu9mflQ
z3S8e4Qg6WGOGQwAubCIKxxAA8izgztA8+wgcfM2LYjmdvy0c1GKQoB8AQJJ81OBqAHaXIpY5g4/
Js65TmCG0z8CiXzuqdf3J+5AJx5GxtjixgiorvSgDh88ap/vl1fd4uCvkIrAvYdxXFElRDT07WKI
TOaReTh117XaHRMx5dHC9sCkfG7BGk1sZ0ZT8IQ0FPNvpZ1XMX237/vHbyNyuPGvgFwCrzS3YsuW
rd0DuVNHNGnDi38Kdl7YAbRcRYgocCnwHJuTw78ti9f4iDuBx81LqRoY68VXE4vSlBH8YhfxWcBY
Sxbh+pVXypC0o1lqDhR7pC/7rsKyhaOT7rNvtx3nCba2u7yylDuU+UMj76eXqA64lFQi8jDGqsZc
JuEOoXB0tmw4ouDgCnpbBI9LzEvueTZAFdYbxuJbrZrlMCIwrU7w29d48nu1UxH5/LojL7Fsigfu
WMTpztRegN07XbQAhf7ODDZTdaF8P+Ue0XR4utdU6i5KL5+0BWbSVN04IA41lfnoZTaqu+7nmaPG
Eg/aNls58eAMV+F1Ni/RiW4kXlkLRA9MWZqdk0qAsciTpIDu3yi8F2C1ct/pp//GKMHM25PXsqYv
OzU9evV4xwo4qnr9bsvrhpHdMTuNUUMEZIGNPyhmM0pj/QMxzf/8qLBdnwDfvPRIige6w1euTReM
urJIbZuUSK9SUAYOD7HCDA3QBIUXpTNcr+/SB2wzwDUIDfMCotI89RdfEPILIaLVh5qwUDv9U76u
eGtcok6ZmcnVJI6u8Dv1ROSSMXJ0KnGmniR87ifhEuDEj7VRmZXsHE1MYIaPqPWgUzjHtZGbdikC
siiB0OejNLhUvffVXIFfyflyghHAFpj3AUt/1yVb58wYmytAzfw2Mh0BZADhLc8OrqJN9zKzFrf2
xqy/1NiwRYXpekuld6jryZ/20NDsMfJNMlhMjQGx/gtpJ3J7JgnR7rwehtaUjoWwZva0L6MchO/L
tR3iCZMX/PMX+TGh2weQ9u8VOk4ROoywMLP6liM/zLt7+zPAYDRdK3CSh8H7/bgLVNKwJowZ+XgN
N+LzPN38tDc+AhVxOk4jQLebBg/lR2yKB3bEWb2dOO3x3o9GIfRdyPdLKqZ06xOPbjWvQxDmTfjR
k3pWS2u4i6/PThk54bG05qTVbel6bJ85N3N8byq6nsxyjCmMIVjUsRKQXeOSIT987gOZlSjQPasu
pRFrBxvyBRaNPtmWE0YTkHB/UtDLdKKsYsAKsvccwOGVIhX5bWL4TYhSaZqNGZXM063yVkHdDbes
af1Chhm9V3DHC78r4BHh90fZ0utw2V8hC5qq3HvK9o4y105TsSXLuE+yBPT3jqluruAlwusvbL8Q
HIg+APvsTuUpENCVW2JpU0zgtWOkYY8A8ofkgkx0VQSOEtXiO4S4ZSrc8BSDMVVKqe4YhSa+NjXY
o3oLE/hurAWwOQ6MmpyfRj2jGL3V6qglj3erwX334XByDmRx9aWW3aJWN8OnBMqE7N7sWu1QCpDZ
rvEnsmo6Hq4P6cUg/VY5hjYJAbOys+83q97OkOJFsOZ7ken9F4h4LTOwt4a9jNZcEeyxt+VWoMzQ
PzK04FDViWWiLD5jWcVruGBLaDpqKASLEFPtuTctmxt+z3Wg3WnKFsCa3WnKedjKevxNJjnmJ+oz
VW0Q0UtCn8pQyZWWGWBrvpJ+WoRi5+F0QLxKrvWn3R8r7RgDB+a0gmf1i0h1gE3Z6LJeYsZrZN/4
yh+sBZAQtHztLjJxWSXWGoSpgrg9mWnmdZIj0ovykw/+scvkfqRUHafeUZsJhienHkbg2RQ1dSaI
cYeOqS12rlH6APkIl4C4CWcXA4NV8vlUJU2CUBJIJYPGIjb8Buas9FQhNMCKKF5ipclYbvCw1ONp
U/zhLrs8UDheW2dMACv+nrc3n4VdYAx2W/43TT3EjBeq7+aOvRWx82lm5p7oTzygKLIyczcNyRng
CrSJZ13fYq/iL7DDQSoJvqklpe20JyA0Efs0cgt0L22IGG2A70rH27tgXAWG5Kl0sWlEOqWcn8qW
Uuk1evKKM/B8SYns1kSBHkh7/Osu2NuO6EFIkpaNhWa0m/zDWBdN9uR19m6hygJukUf5VEGuKbsg
FNeJEScber8OCb9c2iyam26G+K/fU9YSrZnaKON6quo9o6JSHWoQPnILn2ip6IVB0w4d6CGJGBPz
aXV7hNnS6DtFI1cd6jUYDmIll/nPyOazvCb8dU5IUQgq+PZFL5aW4ecNwzHEdnsyrqRswYJROjFW
x6nkPfGItgd3OezrJWW+Ft6DZYB2RsrsQ/SUxLdtCvAvGrY73MuObb9K275h2H2YUWKxO5URPhzV
pWIP26oh7yw+ubn9rGZk58tgrcsg7xTnGB+imc8AmfMT0bPNp0xc8uiVGFlQpxFf4z5I2SbFEUYW
pKECKGJ0PxhmNDPHyph0uOZ0YlEDQYGKlQBzGrXLrAS78St1XNC7L784+Ne5jVYZCZBw4o4i8zW9
EtuBvsP6i+1JEvYQ50i4VeMFCWhVrHdZoC/VQwR4ZfTlH6iWBQmB2odtPt0O8JnlPIFk4voxGifj
Js2+/dS9V04AlippwSudUQPJhE8b9t49NlTo51IQvruO4hO2sCECbFa4OEWP6PQZfnhya68wS24M
ITqJeQC02vwYEgaeJo2eABDXOfPXJf921uOyzy0Ps8AWgv0ZQGsU3Iae2HM8QFerZy6pN3QUALmg
Oh5kZe/84/8+Cdrdsen49iq7Fd31CwrYNJBrS6TUoExid6+yDBGo2NMuhbqlEWa38qYXEhSv6fOC
it8BmiM1WTW6GZYU9ImGsAWbPSfwhhS6apqWxnGillgDRhEZK4Foh0j+FpBqhMzZVRtU209o+yIE
SHJZ3lscejl9R3fEqLC0VwtHrU+jD4JQfXalbfY4cCPlC/GGjHCGmqHactj5pemFSy5QJsr1cGdk
OGagJb3bc+zKPndyew1SJWvaxH9lkQ7fTEcDAR/FwPlgJCnU8WUpe8jOZ7qvPJDkJwR4Z9RE3tU0
rLLLI1mX8trrS13+woX3GTgwc6owsEZiyXhVQ35+XDbpLPY2aSf0PBinfR+JfzXN9Ab7CIyYF/Qh
U9nVZeyDJLUApVdfgg8xuqv/rHnd5wJlLNSDxyI3ixexedKB2XtfXTe09qBVSxPLXd3YlBSgK/ui
XZLaoDIn6H4gVry/L+bxOz5UpflLZkzT5DrQKlF0ERf3CxJ28EFNfQakrQwlfXO3Z5Up+VF95tZv
ppQPDsNQAM0DvQ4kl2wFGNXjRl5vrbrdmXyndDeIi+mwShBtrY4/uQ9OmNlbbiRI0go+heizw0U9
dcZPk1nQIB4cfYXu36VqfQPDHpTpvfpfWl2qyFPYo3vrwdqEntdkkuYqGoVhvQSnV/fEf4wKIs4f
yIB7iEAuGYAmtIbrjH4kOPTQ0u7g3RKu9HTh+2KhDS7Pfd1y31qBruO5Rtuht1YZd2/87bHtabTS
SW0XM/VBhcHolZ9qiiWziX/x7HCyXsFJWCL9ZQj7oDJiLfvFddfHl6RG2EwtODs50VZ4VwAwc7BS
7uZ62YlIxb92cYYKvJusLAlvXknZdjp1Nonduohe2JsDiuqYqssVNJ8GuiL1kGHSAh+Cmp8AX2gA
AMtUZs7dxJ9c7IyVvqWG8G4++NvnIACuKUGAhwpsV3XTBZdiP4yMIvbcUKGiEC7ITrAUhyckOjVj
IbPJSU40RnZ7iTgih4RMwYJtLqQc2Qg2W2TQkKCLDcQHIfZ48nMce/WhzR8RVe2nUDKQsUKGBVsu
PD10S9liGogTXkFP0rxezWLdT+8WJPOEKZaeMKMeO+/BmdXDrC8Xvu1ISI5WlYzEpZv3N6FUUDdN
jBD7vZxEtXqAyXCUd17A8oaGu79Ge0VUqESEYGfOS17oS9WyDpyufVK0jfylD+xJO1xt7VVSmljn
1dwrN0nVldg31aQ8sxfowWgNdxBEah3frOPCKW3QUmifOeDJk/63GHzEureIAgjpOUppbiwR/1r0
PQz2SkZI7oExjBhP4d/gFbWi7hr3tVpOOKv/lSCWttIvBdqXHCRDpODQUDuE3CFZIE8zvbHIDpa5
JnE1ka4kPQqJcWH3KJjBzS1vA2n751qD7KsExQJVI7ngrbDOYekKUNkUxtb4Pzi5i0ulUSFHG1KQ
FnTnx7dxO3t001CnkMHPjiQe24OZCg7wdpVfXgqLF1flMBtKUMAASrdpNhU7G7gq40XvacQlfv9c
y37BURFmwDybhdqB1zdPGBN4S0ER9hRmPq7StYJwkHL17Yg5Z2XTUVa9kGyksHEPY3h2ILcbPX3/
WwD69OaPvpXG4KDYFBbUY2Gvg4vi5zn6AwQs4rRqzOYB8WfdAJceidIrHnYELd8JkugTII5NNu2s
BHw403Y2T17mxI0R9V2XSav1OsH2O9j83Kj8WEj50DAwIp+dtRJWa5P1iU+oCT9Iaf3Jnaz6Q626
R2vJVdkqJXCtVL0eHbNBVWtTbsvQaSa9cFxh8wBU/7L/dgzosXUnVqxj7ApYMVBkkGdKhpf3uZw2
M53N0lGVdrUkl9jtkIVMLYQjbluAd2osuzK0h6FBUkgWnIOJ99z8Qnw21XkX0x6vUDxJm0CY9NB7
wuZeYX9YvwkNeQE+wzTD0BeQ6vrx5NQxKqm4N1ji/WGQEfzD2x3y91/Ekz627O773Lr56QiCgccP
RLQAYmEEnhOEGBJm0LWRITPsrpuLL6at/7D83xmd6IaQjCInz4t+6sQtLpC3pB3N+vY5bIyOqGvi
XzM/6iV2a1zxNxftHArzj9zHHeIlDED32zdQhGVZWYP4PjonK83e/iVFvTALtayGRAs0i9xckpcA
YixOHeVb/BoWs3mfdeE9nE4q4tYddmvUwjgwb433VExbcjOQzbMOye1v8tTOhsVNoIRepl6z/x7i
tPkmBcYjHvVbSSYgZPzsfWf9H7026iWuK8x/bbLPf8ECWVS2naOKffyptYKjkUQXOnEAfE7WTM0Z
kpu5SK6bTm9WTRO+a1+Y3burLJec6D9V1ne9dg1qWLFcPccPxFZ9od3pS/ro8GVSzwHyyR2hSMoI
HYA3ZPABuMtvQ60leIu/rB75fAA7r+b1TLNvJ/odNacfAjhXwZgnWW/Kg5IllYVAKp8B2kZh2Ri1
V9a90qf+O0HYjQ01wRdwBAwKrMTTmRahu1GToagmk+6Rka+zYohJn4ayZE5+glVIrtpCwOa3eMpS
pTA9+JJVJPnlbw5XF07e6Jik9Y0raz9eVFYVeUWqTXiJ+Qopa0/Ybeh1X3yBBMklvGK7EXoAtHCM
orniH2rwVaoqeKQvguWUvVTbMK/uAjKaJ5x+MTlXCIBALjYW5QvTMciOUu6cpnaa1kT6YB8bopJo
P3IBOElEgCOYVpLMPe5yxh+3mQVRk5maT0mIIE7Ft0FNBct1fyHINXCBVVzAEuWLTCFuKketDVan
Y18egDdUovmwh6nb4AQTBvKX2qvYGvfQU5Rm8QLvzp+40mMI48DankGWqHaSzbDGpgAWE7GkAXpJ
z0xDQIhRvb7rsmXjfWepTmlXAU74DqeWXWd9hl3vrRmtHWN7kXRFNUll/HnGID2vDg5t+O18gE0J
6iBU0YCOvalD4HHn8u1E2bmK7z7i/Qp3Iy1yLQy++2dgFmS/Ly1wj4TJzGkyAO2QLqNv1mnXbV5d
DmffhZz4HogUTna8U2p48r76EdoQkkRS9Fz7cCXEx9cyoBLW/l9Jot+1xbaJ7cDlRgKfTKvWX11n
HaLadlXCv4auccYNAPsncHp82w0RrQaKRbzeTaVp8VGSwb3b6A/j1W8pJCVbtuA8H9AHZLG1AKm8
U3av5NTp5apsq0pS/v2A3gi0CeuPxuweHVLQevh3RVQpZ6Ok7bXGgGb7PT9NNi9sVyfRdheoiUWG
hLPxTWFWgrXWoJAkBfe+YHxW6qU/caDc4qNPWzuRNuXTNDRWqExkvL9w7l5o3bULAknm860irKhx
sgdWxDYtSfFi2s1oyjDx5Q0Cf8+LcE/Z480YzS/a7U9gKS5HrZ97Tus/R6QSAldFTAEuM0cY2GUw
H1+NyYJkuIc9bmv+mLFqvIHrj40PJY/ug4tcXyaGzOn57ExwjqhPDltiZ0OrnZxsTz2w5+qAXcV4
MLlsPoOtQs8sxx8q+KDDIyf4B53ymuRL4EhHjSjn3ssMkXR+3vjJrI3lYVwBSQrV9CSnRbZeFoZK
zqexYICSAuO9Q+/Af90wAcaLAD08V5oFdFJoJL2DKDAaDi6EPptcGIVhmBgV0bDjbLpiFsuH9NPV
ru82+CNxUzYdDqF/zjmemY2sRbXnWzMlANoRgw4cdaPzAE82fUjSFaVNjZ8d8bZ8POVuRxAs9sqM
pJwHuHG/FwyflocTrH+nG+i/XLorV2UhUAN/8snxp53m3CqahxtLYth24PP4LxgHM5E8xTG756li
uWQ6UE+4KTqIEtPSK/xfwbg1280vRglq9vU2mFy3Dr8e0KxpD4YapG4CKuhuRDlj/wUHZ3wUSL9s
hoM5YEpTXv3MDBpI6071H47gw4PaRcsdXqnhc9n5NOskVsqXfDDMnyblegs8f/8mNDjBHcluQbwC
IDAFPyaBL5vjza5IkOPZXD/gCl9M0iK+MFCWPd2p1k87dADknAHeV6WylnX+OTK6GGPtzW01D8st
JkkImYrsBk6SnJOFap23kCZD8Oq3RnbyoR4RNuRQXVU/YpWcPn8kwfrNJEqvZudIJAN9jhbmvdDv
QLNKht3/4cP+jBcCK0FE6h93Qk3puIULuKyiPw2v7PNx//RQf6xKu6FWG4yWsUYCJzsFMvEwMZNa
3HlNdt5E0gpZyGvbw3E1FeR9SkBp9Ey/jhDvbBosExDYyMsNBvSsyB1Vit9Wwd3Pt/K0/pyKKyKG
UBUjBR1YIWudria2WVizuFLkswn69/S1qjE/vWp/B2yxmNo6GcjzDRBcPS63tlzGfdLuM6yObP9r
SNIFP4ikGXLMxTPaPkOQpyytGudQo+sRzKMiX11mss2IDEjoPmSToVy8obutj6an6BXDm/N67GCx
Faf7GCSr41+bKSYWYFJ08QW/bNFQ6lBnjeYkhauKoNAUsigyNY8Lw5CfuSVdYNAzt3D1L90zMR79
9CjhW0yLwLKzgjISvlcg1Lx+2n0N9ApwSdlvIG9WvWmCdi8x6vm8irM4voUhbTiRTY1lI89u5dky
GcF1xYXSdtSYGStceoXPE2BSQ9rzI5KIg6FBI0CTrZ31RcK0DmGzQbvLbay6fmdywjbCR5h34IN3
CwZU/0u3hnaWjvqzOQwSZWUmypyHwp0joNNn2S8Mmirzy3NTmRZMQ08VsD09y0omHhsA7s/fmpjU
Uv0UysRfc8ERbImaZ6Sr9OCDXBwx7qqru+DxjU6IaTwqAlXD/Kbfb5clajH32h67vxu1Zj9tbBWw
ju+OPQG6VGxWDReg+ZBgVzxLxqs/+Pyy7HHwXH/I6DL3W6W1M/JmL6NZSP/9MG4Nc8cllyVgIRVO
0qtQmf9KPlbMyqMtgf5GKEhPTR+b4fdcvLx6VRDwv1qyZNduRdNXDuCIx9X2W1t2NcLqw2C6uDuJ
O8rjyKDTGORqDOeJaQFnQXwvumeQ6RK0vy5Aej02V5HfGAxc749z1QdQ9dvMUiPvKA+lsURRodlI
LY9C1sIgt2xdlJent3CZYDzZBP2fb9Ue93LT2OTGsdOtTSBgxfZh+o/iCwFe4qpyXoQvoHHCxP47
hK0GzTyBIXdDPD7DSDtrQhdcVbMni2u7Jqo9e8Sj6sv3RERJn0zVR+EC5oOFtkvFX6VFrb6yRxmK
lgO+tC99QKmq/3kcIkp/26fNxnBfa+ku9DZUQ3PKpmjXM2jbNEgC4AaYCZ8DMW03jJJfBQD0pR0T
JmQfHhXTqlBZIUm5QFIGTSkBhthDwYnlBYo8AyJms1pLPa4YU2vmj0+UzcUlfiWfJrqTEW+ACYYm
7wioEYIxoOZbJSCAP7yFrwPLUv8AiZz5lFiKpGjz3EayeE9VHJv+u+4TrinCMJTIospsZk36dROW
gTHtHXUb6nxZOBk0uhdnr6+eeYMHVKM7bakpO/+t+Xltwuqw7CL12xrLImNwSWEi52WM39xHr9SE
rFgHCEjrryAdqXTffSLqlL2jpFBAx58H52xiv34UFjdb40QtPZYwCAdCHgtTMZODr4rfxo9CYsBM
/6le7wBBVVP/53843G4uqJ3PyGZ5arMZIoV9WDk7ErraqW2NuLXFsiDmi/Ls8xPR+x9vxI5ZkycK
Or4rtO+JLhhedDHzLl/Zt0VnE5YnIgjB8KtuOZIQQTwhKwqyeqxP4E5+vVhLlCR5K8cs74LCGMlX
yDeG7qzFd00OvzYVGQm3F6q4tIsp9DuvwdU5rGm5dHpJokIAKQYGONvZvXJBHctcq+Mzbqm2vOdg
Yi1lER+HzyFMaMkw5YK4ClBrHwGVOm1T9k31i19l22cEaeCw7O2crWU7+vzFr7+mV85EG57Z9fUa
5k9PKtIdlbDRhyvZHL57A8lIat0RNTHOCspfBhhTNlpGItb25WYiwG8cNPdeweXMqIcfpl+gYbcR
JPrP9gAMvTZfB+WK715LUJfqBQcvS3EPL6McxucbxZjmXGDG46TJIXvL/i5NaxLTCL1ao3xDHdws
xWkLYggrZYdlowm4Nuh7corDZTZ5GI1fQ0iNzF2LcaGVNLwTG7xT0JLySMcFvQcSbvo2bDoHlOEC
Il+wS1itL7Wgux0/zVIhCT+LqvDKspjWAiazz/XATncnF62e4Xfu9YfvFLlM8SZaE9vCC/NTkm0/
T7oAeRJvuc8NH9qUMU1HM6K8mUQB2ONVEcCKxUIYh9pCeetjn11LZRxEONRCmHOznjsMxL81709N
g2Vc1XY5jk/t8SlzDxl6ZQ5JwZLTX6PSSGzVcaHDw+APtqucBHN4B/krwm7nqdIr3BjOP9O8fmdW
e84iOWYtJnXaedq6B7lED9rcxyIzR23GTz8lLGRxOQyNXHU9u6NV/uVMHtDF2FswzNZ4f6y34kfM
SKN5VTLOnHVNxtDZKzWp2lR7iMYg0c0vxEPoOahN1f+HHbdYKm70eNLQhqGdlNOyNPbREkp9D2qO
kFZgB0woh7m8syF64oXRTU+5BfBJ16qXT8Y/LwJ8grqkKoQJXrmmGNW2AVaI7CVipHur2fXelQsV
Q+7MUcL0RGTa+fFH1LOlmU0wegVso2H2MMzF5jnR0viOGfEjL3UM5T1EKX3o74+P/T92Q1ReLmjU
2ozZ+GzlAAy900Ul4VCZg1Mac4Ly9qVVFpqkERLlo2elu/5ammQjJYxw4p4+4dxf3Zx2vIY8wJqO
afKqdpO7WdDdWWHlstsxEa8f1LvVGmC5CDjezKyy5jIYciL21vFm4atefJBjNmyiojak6M6U0JsQ
xuWJLNud3JO727ObnmHcgd1qSRaMDuVx7y3NcISF47fHTDNG25q9gaaM5nVkwj1iMH0LHBoj9Lot
ZL9KqDhKe2XNck6NiMb2yuZTCkC1GMgETZJoIvIF+9Eg4yUMKAhV4VRk5qgD2hdqUoUllxhYMTcK
w8MaG+0dB3zGJ9waZLF+fFVcT7Erq8pr6UmEOoD4nu0Smaq1RPQ0sq97WKnSVmOGiNG1jr11pcS5
fUYhPBagUJCjMihg8os2c2dsO02H2AET8JOSM4stC0HYaaVY70xSDrIKKyPzqVT0y9BDQ0znf4iA
BnFoIBAIt/5NHktgdvHW3qcipkzQvEQe3bZHNkKsgMeHbZNgvCP5+4lgj/ctoCdE2mPhVZzi6ojC
h1Qb2uimPubtjwcduF0EviSk5vD4M8G5/5q6dbYFbx61WlIvKJOP3nsoxvYVlzcCcokRi2XrtSU1
NRIJh+ZSMCVJiLbivkQHpY/RuQmITLxxWk9mecomzyCM8L9SAPuw4fkNq/XcjLw1muoDhd/UtA29
VijHa/yJyriXulbQLM9Y1VwzQBVQBkGZpQA9srDB4Hul9nxZp+2Ja10Pu6U7vS1nA+MYiXZIFu4/
kM/Dp+pz24O22nTAWdLqUJbh0nGOAlS7icTgOEneJHSfnsFWqBjWf2ml4pvacXRPS/jlV+XHU9Dr
ba0qx4vJv/i55wQ6iRZutnbRxSW/1FRQYjGU1B/8EMh/WSyVCA13+Uf1ChuFmOzSWflO4GMtAMtP
qVgb2OET9OVYnQqGDkuj+uoqO7jr5/xYzrGFff4uj/MeibaYX/tjyZtsF9/SVeoJKii0J4MRDTgy
C7rAYUIg20Q3iBkQvHGkQJ8RWm382diJQfydExvEYo2AW9KI4/5vrSk4tkZAgon9IhimP163Sfh+
60NIi/G2cxkndzGeSQqf3s4ttkul3CATTexiooOwvRQKnudSqbNBIvCK9BNcKLCJ9h0etgX6/50u
JGhYfrKmyN4vM4YY5BzoKKlO1soUFi/YtxddA5J7FYBUxYGpiHJSW678qwKAKFXUIdOm1J8DuSkA
HWj968Ek8yYTLX8+qS1WEnk7FYvcsYaoh0C93ChJwofBtDJnKgScwBnSnc0ootShQbqtCJdA3Z3j
2OpKc5w0TQm7cI2lPF1p3B2eFDjZGdrNZrlb2DiOD1QHxghB5CRgXbMIfoyBZHqzW7boeL8ZNuHc
F9NYvw/9zMIij2/CvvJlLafW25eUonp6KDCgM7TWtvmehz7furxlNYehXe7mbFZdaN5iQaaLEBy/
5JQpn/q1TsP35g+uQGMnfwWBAlcqMR1ny0WH44ZAT2230WCiJXpV5ZiVNItT8o53oxRAtK41GsVE
fKuJFb4IK/Ze1TVKLsAMBlEDKLy15hi8//F35MMFY6s1bdaxEJBp+/PrPiRWBOEXIk3gLLxvAe4f
Jt1xiJNS2sGSr7PYDHMGBVbPK2UHWxkwKdeEfdwo+LCK3GwEmZiQ5Rn5eOy0EfFWG+w/bdW2zx7y
H2LbMibGbCt5CQqlbbzatB0EBBgc4Jq3bNlKl9/rFnSBxReYbmXjZPBtNIUGF53G4XXe6rMz7mu8
dATtF4nGruAhXUQPYk697FsLmHBuFR5B6wsDLOXk4lzVc2GB1KRNaRMjaFk/jFQWWm8d0+bV5SkO
e3ECyZscpSvp/Sz0G11QVBka5NThWzlUoIRVpE91XwSTenlNwMnhnMnZyTHNd+F95p0PrmR1AUIL
/Yh+3En0VqsOtjJ+PHKyu1jTz6YK3Q/9U6Gg4C/oSaNdqTVDmWSR9GqwIW7ZRZtvPjo0oD/BSQBQ
cz4YQUyjHkeMcyOsRVgKq68P444bGo9atirdgS9BHZ2qD+Vt/K0Bnz+W+bvFaOor0hPhR+n/CdMG
nJ07doWaAoypB1BG0btgCj7lzCYI8EflBCQpfniB5JmKzkp3FmTDxPFtk2fa+m7HhMmp0iEMo4t/
0Nl8D9DUtP3GkEOgRHMfSya2HM7j0oWPgMES/cM3ora9hw0fxYYH9vIYtHJgfluPwbEYSyawvIay
7KkMwDm3q2eVS8o9OJlopG3z542BZM99cId8EzAAvNrSMSm4EgEsJW/cAA0+AUWrklMlgHMbvnj/
tvNiUw5/VfSviuKmkXweVwSjk8Ya9x8/Gn1zeknBHCg65yvlTOFxtchBB0lPc9v7/7nIKmDOM1v1
eI8Fovg10U9MK8q4mww5d5KGxR8nXotaGzgyz4UHKC3vwO81ilcplSSuNt16XJIG1tKcJVVPL1IJ
Ipi6CkqWDb2iTc/WzLJv88zf8aM5Pq+vXP4FvKrvJmKPk8lG8YW2Byk0GicZ5H4VD8rlSyufzgcw
+BOSzYsPkrm5m0GnZuSz6QPuowO8yCCI/Qko9GXSGxBm3EtLEp9/x8ARkEZRhzTyzqdTDWiH8uR0
V/ZftuZ0yuh/ub5AqsXmmzj5l3avsx8yZpXYTJ92VTMGDdm+CIveBGJu+FBj+lmR3BQwzwVDK8s9
bJ43uknNvWUPL8Ojbc6kS0EWfcm7dJ7fXEj0ggLsbKLudZwQ64HnxZQWCmUhCelIZ0M77JaYBOKe
l5S8Xsq5HLlSUhaVmgVi84dKxG4VGrBWyJV8tcSG97xDFYHptELrapugoMi3IZb0Vp8Djju2UT5x
bajvZwmw5aup/az5Na0m2YeUqz7SPKW7H+hDRE+B7OPpzr2RvjXU+i1//QTjQ+69fch/6FwGE6Ax
EDlFHx5e320RFVhhztPrcBjkN6Nfuvdr/0FOoJIk1E6S4MA0TGf8K/dWR39hI0Z4JxrbfWZAikDE
y8CRKjSzRz+MGlyxrGzWgU84x2ZvURdpyajWDH1QK1tDtLxonczqjNsG1VQBaNltsiDKI9DylLrj
BUyHe56J2+AnLIUF6JKtMb+Q/hkUvbBV+YzSbBv9Eq+5hEoYB+iqmmwf+oUDM9m9ala4ef+ZjvTL
ej8OSrgwM+HjXYq/uYilCszrKeFEfYxXqSZ9uHjYA2KsQo1zzEoSCrxhuH7hK92mDOmKebnO9LiS
NmKqfojXoYwuC27i5OOWUnFvRIcF0jFR6j71dyqyjdQ9g8xQUNVfeCmtWMcHj8uZLOYmGvJAc7VG
mu4PocEXltz3+55BLopsnv7cINorhmvb9BNd890rqcl+D4Rx/7hLoN+dsFrG3nM1FEyWYeF7yS8O
TmfzC1jjGjCdtNGaDbkOGuHltg7nYnQNPnNxQClUFjnLRXrops9JWuMKkbapl7r3LcLr7aEidt/G
BmvQH+1ilESjZp5tRA0udBKfEp15eSU+T81RbqQLLGPK79lK3V2ZwoKuwzLN3lON6PVpgV1sG6Zp
A57jH9QyD7nyHuhdhpkwHN1bUMbRn7aHvridEAoTV9flp0clBuhOGA+WKMaz7VGcE6HSHrjHS5Ie
oymcqhNQ42yrD4Hot/z8IOpq6uw+gb8/Gbx9u71xYBYWeyF81Owne3ZrcjtvQWya5a4K7lN7CkEt
cDDihtyAWMVjYhSSZgBGNpf7/h1FcVRLrxkFZKutcxlvot16RORnQNlGkuDx1ALyqd7BTty0JvNP
A+pi8MrkWGgxCltE609x4P03tmM1trDLFzDCivp9sh9XxCqjnEHwB3yt8xje6fY0+vc3x0EqO4Qj
HFJCRNqt02hbudXWT0iQpD+R/l3UN3rGv6lvAwKmXTUx+WK/x7nNBqy6/jGfTll2I+MALET8LN7f
WEGrKg/pJiTsfBQNqsPki3aAxEUM5TYR9RxB5tenXg1y6Krkj5xlHL0hJRQlyF7XAhxtvKg3S5/R
94R//WQdvFton8ogvDeK+u9Q5rW24C0TnIBbITWes7mGNaFLl5Hn0/TiIZ3ZiW7FMDAZp/z/OO1F
lxcCuttFD0qYBBLAh6pezU+4A7ebe9IKiZ0DOlFBVH+H15fpPlsh8qC+6CAosfct7oaJ0UkDWqpF
8Qt3JU56/wbfDEAYZKoZhvaN+WLQCdaHEvSk9EMXj7SCFnImpOAGBavaZzDPvRPK7vUhprJuHNp9
RAyN7nfObbBIA9K+UsYWFkH/BdSKO0MOrdfZgZG8eoALwEtxs3Z7DJg9PPe2XLRR+gVVV+NRm97L
4eUYI3djv1Qf/4RNFV4tWqPaO5j3JSznKFfY8FUfaOepAuNjDUBXkOEdspu0Wkmg8C+PKQI7mogN
maUy1evxaHFynElPFPfjdOjq65KTVczCr9Hr9EWAnE5xA3tJ9urumCBgQQOlzKt2hdgHpgbAIBAO
nBXo+MK6EtFA1lCro3y0x1jy4HFCNN7fDUK+Xv4NRh4Tl2ZoTkoqHvk8hCBiySwyO+W+sNvFq+Iu
+z4ZWk6xApJoOhN7hNdKWWOP07i29+lvGerZ2libW/yNc/xdksTgvlYq/Pbay2gYpUUgxrUbjHDh
fYG/sf7IUO6xyXxPL+B2ucGHKuMn3dJ2nwWdibkcMTjbh9Db1MCrYNr0pbOZmH0ejSuAe4PMTqJR
chCXy0pKkyb0Y4NCZPquMeiJTzSpwPO9bjKJezgbEQtRxqn0D5nzRNsd9hvkII9KdUNeawJ+CpJU
HRR+mSEurHQqMtb+HhNN/coK/2+Q+izcXAd7QGb67xX0KR4ftiEhKdZSbbWE8YRDkXIdz3GYZram
WLPkg+1bJpTJGrV+L2qpAOLKo3sPyXi7CWNv1YPvIblgkZF8kbBYctiUf5xmq+1/52Id5QJ0oi7j
ozM2vVPSpR4swCZI1wmEeqIKbNE/x35lCB2cYYDynqI4pdZE5/8LFaGE8zn3xDCr6usAC+vt8yp4
KHRGLNdvm+m80LmbebIgjbMPbRzOy/Gmxuh7DIB4sWj7BG0YBX8fjF2YqIEXtYS5YwkxI/5ogKI+
Q9YnDiD3LU+HnTsLJPWPwLXyFZOR0fRP+HZCM3FVQzVoTwOA6r7fqXltLahh6SsTB+sU/lLM2JFA
0KqZUZcm09NVYqN148r6oxIfRPZVOPttGeLGBACpqm0OaKDmao9/ISTd9q7ZQWY5fLwueBp0O32y
OQVUF7mxB/y2pp6gPoew2/D4Lg3muLgze7k4WPBWw3brI933mD4Ica6g0QDgvkc37HwTw2RiVjyF
o8NPfrjvc3gPWVqcm4M8dze181W1As0Ryvb84nB08brWjxzezlR9+uiRsIi1XuNSCVy9V3I9a9ZA
X+YPVitAKhLN7Ytsi4yozH7fjyZNn0qKx5hmlGdeX/yXyMhGgjtgxqSRTQ1EkZIKl1ChIz+Y4jsj
TdUTCjyFJcui+m30HIQRu/nh6rqh9Jop3JuvbelZcf1LAyU1CwBsmivtqxWJGZmwHX0rGmv9gizS
gwqP0mZzI7ygKB7Sd3GMfYUTwmNy+yxdF+b7N3HS7b4YwRGED1AqvgY9PB+RnME4PMoFvzpH5Uy9
55ePs/HW+oAfPVrkoi/lZNetRuSyoHz68mxrN8b6saAcHTCxlL0ibu+lV101cYE9bZbA6md3mHRF
8oTxTxB9dIHGcQ+Z2dktWNOrqXWXdqzuYaKMAQPeMkf2fcbMjZ96AKd8J5Lnqn3ZJvqN7SBspVeo
wsHyPq6myp6KvP+p65Np50N+FFuCXenlmx2XduPqIFjRkS32b150E+wv6yd12V2qaOaJB811TX00
Qa4GNo1mXsnqOaIvBtKRTGLXJ5tetBhrxxPAnSS3fncrzYiPjdWkRRT9d9o2OEsm0awacAkZ7uE7
9caal8jLgr1lgLp9quYbVb0Ej6fDiYtTnfUd+uPmAOiQoUN/52pD+arpDKbc9VLVVW+S3f8hgojt
LcE1DmpKbW5H8Yyxro36RhXr2SQ6iPCHLlfuEbsvz1AjER+M1yfaSyXJW00eUS+cMsC3GbGqV7If
AFF88lisLQCoZ4KJjaktzbRsZwJZTwKcBaohGrPhgMYIXEqgRA1+vHScdbk+OuImwwk106L+4bWs
59g+pnaqVo+k1Js1qAn7gBTv/URwyQyyoHu4Oky0WjT1YaBkFKlyhzaZihLD0pSy1UD/8hXOE8aQ
bmofWR0k2Evhh7rSctAcwU3wPuHKpIXQLFqxPOT/5bMQRgNArObphsDc7pjyEx7W0oyNM2jNyZZD
YzLIelXiHcuxtGFlvNH1FqlWBrPT8DZGWjsCqFEdC1hUfW5SIj0Xp4wfPtKbMr1D75fdd4dIepHV
YmqPsujaLuEGKJTwtd/mh7F5RqdusS9bi0E7ViFcFRexjDQNMkiGZc1PVLZYShgxs0WdY2O964br
td0m6VuqxUCShfWc1pcw9VujUfugIcbtSXtKsLbYBY4NoEr5D0Hb9EVdWadUkds0GTIfS59dOJUu
iddArEcjBgHXGoENGDiHcUjoR0UmDTat/4QaJJ/un12s37/+17gp30QVZFeg8dU5SazCcQdte6Qe
/CdjOVThzu5WpPjzqyyLXHDpeKil6twHX1ctehCM1MTv1c81g9dbp5bSUGQuyqtRtSBYJZGeZa41
tLXDN4oC71BCn8DlKdApig49A0VG+HVDAwYTB5rZjILZKBHGDDnG8PYbD3SXR6+g3nVKUOxeAwcH
OQbpCEfP526WAhVuHiL10S7KIahk1fRRxMoVzLIzEnm3b9FWKQhNspQy7QK5KFjXN6isGGlZcCxk
elp6h7yU50ct1irI+7cUgAxvV8cUKSzJK3OvCBADG7/ghJqTEDMhRsakFDaDJ+ybK3IvpeaVLgup
yUDnMhheX7IZcv7tuvB7uCNe4cXO/v3Pgt403DUyw0HpQ/BsNxoTJQBDFg8esFCgKpSkE5Lhi66y
wFsKZaLhPcBmgZOJlGTX4D4cPjc6qV2hMZ9YO+YB9N1CfGx5Ain0zLt9NQk9irs9OPATITM3R254
1hWdMxlK2O8fdcY66/SftO+K+Q/CJoiH6fx1mM5QDqenLboT6WXkmn6IL3kJGlObgGPx+qjiiXby
pzMJvkpp+y+yO5S4+ZfDlNxaHw0X+Q7vy5weNO4QZeKEHWJMq1KdjKexcYW99DD+E+PMmlyYE97z
tqmQOMacXhphLcUowAHLXbjXrfnSbOOBmI4ciDHC9RTKF6Rrd2r2W3A8zja1vTeXXSYYohfMyTcS
dNOktEQLYQ8u5PpkXbmWiNhTN/GkR3zg1BQvvM2VxDhZ69DvJGkb9u1kWh5wEG8hoURpwvEMeoIf
b8VxbVm8inVOKYJu0qwI+zbhRHVir2qmTJpZvQu4wCOQGA7lcIq3kjOVwFwc1YctRTQLeHT9mc1p
5xPCNy81j004M2AW1LAHekOgOuEipUU4iGxMQ1exgifn6hF+qn5o59pcllQCqrf73UF+QiX2mUtM
0pl2csSwXqFRcA3Sgz+4Xku8XAUQ5vrHImLRbaTAILagI06k+GAi+VlCynoheFzJPkBwhQflobiG
L1QXRBfmPCmz61um/1kyPv21xAfODFjprOPMUvBr+4Rz31jMYoGAD8z4S5bu6MQzO0bLSZR8Nzb5
xyNUlHlLFUvfIti5Ip1uDJHjF8WXIb2XGFDFmirthCgkYBWUgssJUoMfIXWez9WhSmKSiCeMf4EI
aXMc0Y/GhamrTDhqh+db+oRiakd4gGPg7IkvBs8N5tv+NeToVK4yNc57Ivf9JPhCvUiTRHwPGkBg
hHq7CVNnGpder2/qxSp4/RPYgXxWzE3UKH6A+dQ1FGLMeZjHuIUF7+GGgt/NptYZIeEY3YnRKU/2
Eq1DgrUDa5pPlO1/XwcDXs/U6yNN2dsf6BaO0JnJRVVn2auk8XoQX31kGf9AatbvuhM87XlZDANk
i6WX3545HgQnEOhHobH2j1h7Y4P0Pr3ZV2VX4hEJV3dPNrAsbhyRpBpqaZKM1PnSJ2/02F/zs+1r
1BZhLrJO2lWJ5kZQXFCZzjyMXBgYVtYE9mh0awUiwLwPVTP/NxLFNPIjiVL4QNwqy8vAn004yTsM
bIRGzlIHW+v1NkSFkbyK8D5ahCAgGQyf1j0HZFI35nIhbSILL6oVNAjmCis83VaexwNEB8Qb/VCi
PQ5EN2Iegn+NrpBtePaFMCp5eV84BFCHvcezFAZQcYfWZdjtAz7ceWNx8Gb72/meIVzET5STRnaH
BS0OUeFabDFLTrwrW6RlZylA/1AqWBe3k0WCLRyTl4xJPClWhny0ozJet3hIrqF/xFqVTRrM+jV+
p4r+luJTE8I5o8AxJrAmKSUY4bsfVebR0zQJ6Re8wUosKTdbeGxui98flStB4p5kXfJMS/kMo4+t
/1gHzsHuVk2Ml9Qp+laIhJFUO1qJAOKxiIl2tuPyMRrMI9YVrDB91liErOVWqE9ooEJZQxCHFktm
yYZdnM7eQA2JhpSP69aHL1HCOszEdtwxGCLyAz+wnpyqB1ZGzbeoqUG2dczbQYJL7SxxYUj9OjQn
QA7TyGoAKVk9ruye31tVZmSxQ/El9ouMGWGLhy+x47dKAJbjzEvMtzzWRz9frE6WChUnnfforN+l
lPV1aLtmGgwZeXt07u+Ek2CuPevtpfCcmbmtXzKMq0V8fwpVmXwJxbYo/d2oDWOM4NKwZ/6KiOGY
Wg10QxIjcSZWm0vxHN+A6tuk6/L3LiSnCjm8M0HaecF6KagqbJ0rcEreg1yXDCgkYAD319BbxLTq
T2CqGDYoToxKH+3KaITJKWFm3SDNBIU3nulRujf5PCSCIC3P4+I75mLVAbN8po7VwyWof/siB2Lb
yN7OJo6z7EnXNws0T+GPm/hAXIzK1s3Ss8GL6FujkSJROQ0oMCWPdGbdcs4mhE+DbNDAbhQE5E0A
GMG3i2Dtw5waP4IgIIgnHSoP6TKnOsmHEzRiTM+wjdOhumiWAcpWO6Xrh1PxtmCTnYtg2wyx+c26
PRKEiHztR0/mLTo4NhVp7d48EgG+cReb75evApqq2NYsNHn0Bc8fH9VsRLenNP0KYBIOGlhzv4oE
sVOBDZ5+GpwuZMfQYVsYg4sClOa3lQILfiCCuyvoy/9Fn7rbjF7s3XcxN0adKkMUc6yKJQQwQ52l
ZSqHKMQ2gxQJaAamMC8RpR8easj2j+/xVkvpZWhpTlQOQBwKTpg4VqLPnoTNZyWfqsNt1nCMQ9tr
p4aqgf9VxtqDWf14YnZJUhVdqgaMtGl91igncPXGvwmWdObKecZA0nxhy0Mv6FHGLOvj949omF8R
Wrl3BSvgJZl+ZJ8bNQSbW05OLY3rn8ZTslVFXFbOdOvK+Y82wv3Ad9D3z+qxaSrqh5XhWbVSFf8b
wTQZEFmwoREabY53OGHYDBbyjO6QFH3W3+RvHDhzEfbTsh4yH6JXAD9501kzfnoibNgKmkdup1S1
rLMnwNce/vxHhCrEdHoFRd2F8jh57EsSPm+0TwortUbIN4kqq7CVauZvVf2VuSaB8pgALpCjqJBC
/o8JQ0/t6EzgYiMWotLgl8Rky8JzPpibqq+a3S7jrUhyH8BWNjlG8TozIx9rytXz78fBQ2JwMmg+
Gw/VK6qLRF5vQo8Lzcip9DHaeXmy4U00+IX84WP/e6Ib9u06qpjd9lXKg+rcGI6x9nvfsiH3bUqL
Wcv9EP2AFtVYYzYi5d+K7vYj3qLhVB+HbfAWh2OW8+Fwn99DT6JFfrbj8oZc1GmKk6fTGVebcqwe
7LMI7MLlEBs7r7GSiZdpO8hiEJIRf+A8WmcgopLbmzQ6UVnlHI3ejMpIR3uIh8SmQZYdNIaFvAoO
L9S2n2gUs0tXT9Ls+6zLA6hWbuLBQUpeE/7cbg0ZTosNaiX8U6tKJEg/gE5fOKa63hhAzaqtyYgv
13BIME8t6bpCAG9uGL2zMjor2Fg7AYzAs6q9ksRNoj9Wkwsi0ZdsqS/uUDX2zSSyOcS82WCxxbvm
K++rpAVtZ/uqPF5YMQCKuMGDFUNf63FcXLDzuRJV2qZptC2Q3uVpPONDMAdYDPVhr3lNM1Pt3xoh
RqKWWgFdEd+jdHMc/q5XI3hr3fpRwomE5ndEood1y150LamZCNQnFHaIWP1gLuFYEWQaCslm8dWj
iOh6B71fa3eC+weXdCU/fFo379s/kglg5GrlOWYPe0L0KRol2Y+mlp/P4zbJSBRC5bTrpG+Qpl/g
Bg+lStrj2nJg7Ze2E8gDmQ70aqYAh9hnViv+ZRHTOR8h5BR8bmd1X6iDLphfg49ag/1H2VM8hcPx
Ps0ZHh24dXIFGy6rg3my+M5YFnol28vM/+uSnNjIXoZm7XQTrG+6hV8Mp9N2P8czXpcKJcDvvEGp
oHXhF1YLEgIoRGtqVSE1IeproYvN2fbjvIX+SgEpuddik+WyGbO7e7Vo1odRTh3eKd17solLgeDH
DQ5XubCrBt436X4np14vXnOjp62OvU2w9Ge4secgFiIFrLsiBasW1A8sb9A4aL34K3mo/HliokAQ
5++wg23HIx6W2zwdONTKb0ovMj7qZuAUXCWnlBH/IrCinL+9u/D5He/hpsQjLyNY+8QSnehE5vyO
HMrTlmcoFdG7bPV08bEFyxGOJIg3SjLNYNZeYDRcv7IbeeVZOKHmfFuIt6fEfyKc6qDALYontUG5
X0G7TjdyphziIaCO7XGAkIIrhsO/M2A9KZQ88HDsgH6XEkfnkrvdbyeUK0JD8VNbCTXS5h8wzCQJ
XpqxwpbLk8dSTzD3ohkogpsPyCwgrQocPn7G7lAUWwWgzsA6jBnVMaw1r5cTVmqwYZiT1jV3KDmx
N4ylJEVYBUzQVfGINA9smhbgb1HxHp701HbaOl8IGKHeF35q6z3IZqHCP8+PU79qsFydm6HFnpOw
DmRp0THRSCGZAwTkCXN6usTk0BXCsFmJcYEswaz6eSHhbsz/Bgmy2kUmN1IF6ZVv7QI1kj1vTvT5
JOVFB2beUzuRtmphywIKu4xyrqJG5tvR3uKeRhOhTYGJBmZrIGXX6dlBbK0Tq27NfKtUWNpuUMrl
5y3HiGk4vUE8R2qXBZI+NGV9FNxuLiX/p/GZ4qtTCn7ElajuIaL17AqmigqyZr/+dPLGK8G6ujDD
3dDYz4f0Ftg6KxrS6U+Jp9H1DRHo6nINL7J0CNJqXDt8d7rQR8Vq79QbC9GkNcJEszpDjtcWNzw2
Pen8MU2I6GgpPKtfjPKF3Q+oWex3CM920EOMwfkey49gbK37oZpgfmF3xH3lQCVYEEg9iuLGlksS
FE2dQYGj+aQPfGhi0zdwPn0jZM/nygBW4rVdmV6ERxPddjjG1sCfmo7w6iP9n1iDscc2IlDsuIQq
7Glh441nnLKCB77cShmRmA5du255U1HaokjTOSYKRiMX9tAxyifkSXKGJ7FMCGhj7FHRvRFGn6Q/
HiydxxJEfyFTW8beY82lkcPHfLMVVnfOpXGy/kQFMfpmc79qbvPNlLzodifgOPlzjkIwREPRBl36
G7vr2iW1TOUIKuIPgG0Fm/9IHkuGA4oOOooR11aQRn993ocbm9QaexiYY7okJOEKiQAN30mkASaI
I/nMYFDObUbtpdEqa0v/FTB3ExW7IEeauZ5VTuxXTjVvRQImTPr9s8R9FmQhxIBveHHJP6/qP86E
sOBijeEMGgB8mjucg6fxbnyxucCRT7ZR72WjPFumbzJlHngmP9+/RzBojqDWhMQje3ngpGPmhInO
NIVEb69TsHFPJdle+tGuYi0QroSBSChm3Ji+d9fRK7AJ92EMOKTu2B++ZK7eUngjquF5jz/oABYm
E1oq0dzlmWX+nFKmUH77NjPHkAfFkJIfhd29D43FyPxKbUaayPtfCpDYklJgGnqEyDIsgqhxrg4S
hDjYGLOnkYV0AvLO5Ks52nZASDSzKT+yOLs6vaTADrIIEQCbR6wzGpotq3TMIoY0MT/3bUoo+X2x
rtx1VZzu1hJhkQx47dXbNYvNEn8t1uP3cI1ERmaNmhY5Z3UOsYGsdnPHqff8A/CHAaprC3TuHbPc
eiSerheBuDhup91MYdNz/8+Vz4uct+MYYVBv+kcGA0hVu8P3EIvHc+RQZK/0U1lozbP8QNETolBc
GnbU7U7qCMpHuGuyZ9dgvBFIHB4igjI+i9sRVWchmasrjH5kBzRryN7zNAyzS7IqlhCtyQG53pr2
wfjxHNjxVeVsXvkVZspoyw50GPfDQNpH16JuDlrwBLgPL0Tlw5r9ipPU381sQTpL7FVqts3qS6XB
cWaEgbNr/3zYzUk8ZM4e6wpnVVbbdseJmjeqjOjDxz+1VYBUF7j0KT0YVZY7q8giOKXlWsT10rvX
RHeER2fsLXF5Gbr1ZqkcyZ6PozWC6BJKgD5vvg9iB46qskIuAqVBCJgLvKvvIe3shW3Qt3Pf9hxy
r943MH0B1y/XuyxVuiynaDMGwSAZ330l6F+waFig8rvacbggczBEISfU2FM7tjrHFmNomDg2DkbP
r9cyaS/R1UVYPsy68nIRqbKs98H2/9N9+sw+EQJvpPsET08+5Byxs3Rk66ZyfKD+20pY/NzJJ9e6
TLd+NeWpOhMeohVXJsXFEvPDmYBkX3Ksa6wONl8SYh2KvPotu5JYYM+2xuc3kRPg/Lkkid3ANGtC
Q2sapf4VkClf+vx+bLpEEvJgHGVhrHuT64tD5mn/ZoTP44ROxO68a7sh74MsS0+kNaDmkm3N59uo
IljaeHcpFyxNcPhWBQCAXP42VCb0z4L5yDraNP+UAmCyfIQtWu/eCKfnsbAh1id+8ZFdQXsBmoJ0
pqD/RaT3enzhDsUGGL2/Ogg4fyJmTzrEypRfg7cp+OzPnUEgKYdd3upWEi/5H4fEAmYAHJ5hnRS8
bDpK8OGlF7/JFeo4oOlrLp2+qmZI9yEtbYzazDWQiS8/cSKlxhJ6BHTclCsIn2B111ynu6BowfgV
AxFKyb5s3wizyb7stiDcigikeT8wE9wNFdQMMAfxcYFacAIbh2XS6VT5F7EosKo5idd+wEegmuWk
Gxd7M29OWdFvjpGjrTkpA2ItnPQjlU29dvkC5IeABvDLbe3095Oju5NCKoJISPPj+FMbBASCVvtm
Aer45YpUsnysSBjdU9/RWdC51GpLe55ByTNUogfgCP3arl97P9fg8CG+ETcydHmt+wMFskxH3m1n
RsxIBo1CPWNy/XLcoQxjPhGUpxilvRJeBOLvCep09j+fwuoCBNsxGXkAp4X7SeJFKHlfCzQYY3X0
PfcJ9uq78dwYPbCRMjyGpod1+g28ImNQS6cqkCwpt5Vef83k20TsMGDXPUNdAHVxcKzUDEt39H6f
7GGXPldnOe4mlWwMEFqKLO0Ygd6PVGwkJCjdvDyxaz9OyD3c20fTNPdW/nqy6fO0frxBmai7ygm3
xEgQbqEzNoLdbRkc7qhNjObt01vJkeFCiZar80tg1uvCtdX7me9nxcixnz3Hb3AHMu3cUBvN/AZ3
20Iq28Djcg/PHxufMyJsITXOerTNuWYNjqmkkGiaBSGvJ/kZSfF/yg9ypAqON7y4jU7siz8w4JbM
yHwSqREp+R1J/qvEc1rEWUI8dOWgygZ9/vgaNBMgvOMXtELHZ2eBzQPQtam/hyZ23lSndWJOxF9E
fwglxVCiIshkQGEkmw2lRp4n2blPZi/YEDD3e2PGRKlT1otormIPYrZxYZ/yqA6nzMqWqN0JgwhV
cd2CHhMqz2Nj4j8FeVxP8ynt477IXX7NVs78zRigXIlhSEPfBTgnSDvQCmyJ7WKOzuV+DNDE0cJS
NrnoNIrLC+WCH9VQQ6rDBB2tY41iETCsy1Qme8DtdcarzK+PCF3qSF2QhqI2+unF1G6F/7f+E+jy
FuuOqtL1oAcPqaYLji9jNK0efYx2/u337cqP0Nt2IYoQset6zv5TnuZeLByKuIBU2MrsYpFPEoRf
YjFUUab3Sah/e4Dv0NxlWFIz3c6dgnp7LEJduyAuXUixbG7oKRpS8cWFfUWzA5bRBXYyVU8eFUZn
GFm8aQE5YofnPV4bcqMNkYUs4gDHonjDZbKf+86rlCcaSFt4uUg1LHgeM4mu5owiFz9zEOpsvnQt
zDkcSRvn3ioVOYyHvxgoetl0e3Em2cb2ZIkJVffSpVvttV2Qy8a0+x/XCwSIV6zzChRWsPi1TNje
AQzeeoqd4/i15ttRMwqTrhYaBKStAzwdkAE99/UwG9zdHQilPoOfbPaHgESoS8SNQC0U3Sin9PSG
BZt+0WSpxUQ7RAW8URKqgUpsxo9t42/ZGXMBrMndQ9sjWpWYS+Tsanv7R2K7jGqqlD1OJGZwRklB
qZ+R6F3KUzaNYeIXe8YTDPm/l1Y0597tf8F5+WihkdWT+gn5pm454LPr9KAF/E72f80T9xS33Apc
KQL8lsjJdjC7jFmeERbDM1G/prYUsimqb7JaouiF+ZBryMwZgEcVTkvJsUFXQ1tviRo+PZbXirjU
GoEDZYXcO8KnRnqCLbB0CIqOJuv3EkF4eyAA3vHmukNlqtGu39LMx1N5Jesh4kmDQtTx2t/8R+lT
La9g6XHQ3Xt0rjiG3jH0BvMo6DwlJlaT76MSnaDoW1PQj+QDQmQz4V+hGOXarzNDpI/UVHHThXgA
Ox1OBSd1tcWQbcFj+mFapY9+wFrQGYWfgIEKbxkEJc6LSGwSjKp3MHGmKzmbDUVrV06I33+ju2NM
GQ61XL6wfAujymV0+DWLI6DSMUaTuQtVQxLAbv4Yi1rkaJocqrhJ630ENRYdNUNBh7jsaf6TFN1v
GoUiITd2pfGnOC9BwhEegoIUy2dg1YAwfLs3Gc7YpG53Nz72H9mTtjlvHQIeFYhirSsRHR7b99J6
+Uf73sei1gq9pI+zJGBM+KfpOYiVouj0u1uzbw6rjZDUllDWIk6OAekky8vxErqIWE4F9Nc68lXq
HogOBkYQDiRTVIZzfQKEiMIGnm4C0IGkMgwr/08kOxQJzXnwW0/Fn6LibyQooGwDk9R+AEok6LFv
j57o6AypZ+INp2jdAVN7IaEEVX2Iif8uin1xz6jgCbr5Ay/8F0HbezjxaN/lk/PtIcFxnXJ2oOWI
+DgAMf8cthyY/X6c/7h/aj6dm8DSDIbtvtlyLuQ9hbtyKTp3bSk27aZfnyhG4bsyJsfhCiIlYkLi
MqQ+A8cRYM9ITJdlQ60R5LX6F7IZ21lHuonRbb3VN8jwvQ3GmtLBEn+cerKyvjDqzdL/Uph1b1V3
J/jq0p9Z7QEo6F8V+RX/GhFl0RlwkZGSQ/CuD9W/+dVFR9m9P5Qc3Ku7qZss86k9wGQ92MWgWkZk
FAmARgdVz64RWLQ/XhSwOkh59USeWdgr4B2OMOhkabohbqS9qaMNGtoqnLdMAWwg00683Q8PkeMp
WMeaiSDup1NbyZ0Gl6x/CqHvf5vaS+qJETq9VDeI6X4nOYYskZXXy78Fe3rLFPlEb0xriieWgWEW
PR2F0U8iAHkoP/o5Hpq1RqB/PtuBDI7iEytlIaFdYS748M6jBA4nYt7w7zTxnRirjd85W5afsPi4
rbj4GWVg5ry1apGoGAZ6nCOwHcBPPj41YDJkwMfP4124dUVQ/6Ot3QF9q8VaElT6hx1CeJE3v6Kw
2D8DY8IzCD/fbHTOB28jRLRx8kWQwyoaMoEFNS36wKa1jhkC2zsZKQ+KSBGKyL6YZfyQiPvpVB8c
54UQ7uuHuPNNcvROBx0pR8WCPW3dChzifZTrfjkdIKzfBD3R6wXa4YFPSkGYnZhEYawCWDWc7rDS
Wcu+iK8iooA7rfJEnfGKb3/W934FhsGWcwZKqUL5rnr5WpiMQ7oFosEIK8VLWbuEyIVW5eXwUK61
fEHAvDzS8eIsTdFGfAw54jMoopeY8IVLGi2YnBaldcBI3zODnUXHHF/tmPq3Pmg6zjuCUB7Wun7B
n9uVEV5pIAM3H7gW6iOUVLL+snjBVDPdmZQH9RiJE+wSR8Y7ZzrCsHhg2TX3Y33wi4dvlZfbodPX
tg7v3lHowUTLKK/pnYYlq9LKFRkTrIVQw4mMpvzGJ2o8EokMVWZEQHdbVllv5HPQYGcfG2P+NSLu
Ir/shNYDsoCM3uFmO9zHglhqkuIzHg0GNuzklj9xdYu3KpbJVrkuiaysdanyaLGRXXkO+eKobe8+
5k+hBls23jVl19300kUpFz1/k9TnkQ0y9M14xLM/fYNmqbt9BtraGln+kEFATJfCLKIrRbZAwint
JRfqPHkprdGa1wXeJsGYWbmToAjQAM8dDG2LiKrI+ekfKgYv1pMr84giO1cA5aeQSfO5AYr0evY6
G/JbfFaGbYKA17EJ7RZBnecyEZPy1nPKe4v81vvXTLZf+LIuMhCvYdlBl43bOrUUK4LZgwNU78dz
/SSQNfGWJvM8xBCPVcbI7DRPxPkffERtJioMCGCuXieHRFcs8EW4Xsz7u8SjOuGqpk5B3/uOEVxC
mZUFU2EHhOxik3ABUFvQmDnvljGGVBDJoCHl8GsfI8kKlFp65GnHFkC1CXTKOI9UPYqABaF8QgPo
wzDvfCtM9WwPtCwK6qAb1P42T9wEv7TPOcZd3xNtpAYLwrNVf3+ywr0TEnltKVnh037wgQOzM39a
ww6JBtdhQoSkcHv8qti7GW1GuzN8AZsZse5BatiRydueRZBx0kWFar06dJaDqJXNfi79CddnXoUo
geBaLRT+tC4K43wa4RD8K/aIv1QpiLNKfslxkXXRH4YXBEie3h4t3lvzoCWySKQBHckI6UjkaM5i
LkIlhyR8r3znf0GigOcmuordSejZfzd4tLjMumC+mAZnvichXSvq4uK/FtN8iVzG/EJwbp7HqZyu
0PA6ErgzDafyKfuvEQqisXXCEnzwX09Lpj1mUX9OSuaI1T3s99mGxjrcNGfrexkCDin8mWux1iyZ
bHqMMAiCvIsR5TlyXASkCDVG1G3ElfaGwoiA/eyH78IHKfjZKA+nxZX1tDQr5BjFMpcQVOVm5iV9
dGQ9/Xl3i68+ZgCYh6D4Qm6Ix02fqdpTsM5KfBRVAgFRHAZ+JhqhxBk/sqCC4HUr3Rf7TvzrMmrc
93OUF9gnZIUGbKL9aZUv1dognHyodS7ass9PR5DZgR1sJ2ex9ydv6YFUi++q7GxNODgm+thjFnX6
VoUNE7ClfRdl/cAa3FATXteD+rub5YlBDoydm5z/qg0DN1sG6ghySNuXScxDQ03IAO0qA3m+hK/D
PqMBSgxN8u8/LBFoCaqUbi7NewZsQRiQ9RItYPbP6T3ybjksorBBAOug+xLaD0Vc1KT+t8ftyAhe
rI2GIr/kmwzWmIXwPuLzqOzjRKPGMyQwfbtY+4o4w1AGV/hppt+MIskvTgVvj4SzH5Lk/zhWOCW2
nmno8g9f/Qbde2hTwNlV8D/7OfPcfA1HJ59qD/Rcfxv9ow70mMWOsOeFJxpe39mGxcf6iCNlUuno
za1OtVy93JwYy8bcRFJJT3OZzEFu4YsAmdKr+mDD8qLrB7X0xEQKm7GNKJcIp7PBfUa9L3hBSLdY
gGn43KAKocNP97INC6Jx18o4abHYFmSwW7l0d3dRpXrHVObMWH3bRsDZTONaCd6sQiFTScePXD9d
pQp5imCO76bQsHidYvsL0rWtdcBEeeaT/xE+W2541qowNWDkPm6eNjVmldesa39PJuRAYroN70M9
Oa0dN5cy1llcf/xQgm803eDZRl2DAAzPxkMcr4mpOASKEmLDXNP2wHLuFnz6g1c3hCip1Ke6TkDI
Aoc5VvEv7sZmpiA3mTi2K8510gLWP8ylO7ftbCO9ao1qnDZdFAdWq6PsmvWgf43oapVZD9GT/MUR
/En1lFeWNSufpfIH9VuKMhVVpdLyaxUsk/kJ63EEhASf+FBWL+5qL+EcPkCU8BAozHhwvvy+EfzE
0XSkipSZmz13tY/DvhI6a1K16DPtGWoDLstkRSjjCrgJlRZGBcuLdPRgespo3GDeYvK9czW+h9oZ
gvmEZC5bmAiUoFsXhEbUszZp/Qn8K0gw1XtKsk3gLFq/YTqb5maAwoLPhKCyj/nkdKtDGAaOJCVn
raNLEpu9bThDbJ6nQJzjCk7LqrlsrVj1Oq4ZlRZUEmAavgRQvlbRLmOdoMQ89liUyYyk1gbrebLf
h6M27WyWz8AeGg9exw/HkoVUf+ODyNaY8aOD3zG4S+VY7zO6PN2jkIrx9lsAxKFUJLBmbVZGD5r5
vGZ6hHuuhLJ2yqB6kCzjMSIrMXEAC98eLdjNFRJphucRIcME7HBBncXW8GGbpcRmPVI1Pi8sCBfN
bTrzyhIw/hNP1Z6wU3qSQVyuWwxwo2yQ5P+4zM/GyTXdOyhY/gLVKMNU+OQlsnPI8xrXeepN++qP
A7YlT2TaqM1GzaFeSWhnaFlBMDoL/Ji1/zAKA9y9tGa29vUK7JJVB5CsE6YcOw4/Bd91px2XZ7D8
8lFuh4sMj6PosgFvnAphPAZl5hLznlXkZuGIO65G3INm8hABs1RwhBt8PEKf43CAQGhzd2+MMwPX
PP6l80AQF3ax84aoYvLwu5G9S549sBlkYYlYwO0yAdoYEzTRr4/ZOfH/GO8E8rxRe7SzDuSeetAG
aBaE7LV4ih70wrkdqJsNRQH6J1U0UCDacmEHpUPAA3z9lNovWINoKUtMEex2mVd802NROg0aOz2/
ZBCg/5Xk4p2CEaoTBBdKZc7byMlYXjQ9nGC05v+cw5zNGCDWYjebejx3fn6mODf9nz7DvSXUpjV2
s9lrcQoX0VilkngKdpHV7uN+rHK6TfcdIBmKMlvl7irkRAtrhlwOHeJKO7If0psZEqee2i/6xq7e
8lzkta+HNk1Yp0Tpf/WBfwAH5s5ScQ/vkKrhX5mx/zCuQbXDxrpF/uxsyEaWOPtUAzNonx/NOxpp
nyyi2ncp1uSV2eIsioO9ZbxMx7f+5xjRip0Zf/b4XUwEqnL1jq0lVAloksn+iDB1Zk6Rj1KUcSek
doFDN8loP+LzDkbErhc2mmH4JwC3Rk1IPDqq8TWHbaX5voHdzFMiW8g592QtFiOLdoCITZQgYXvw
EIhwMP1U+wIW5xc6pbWmGLe7mtyQovUWrKdchCXaLN1yW4AP0mW59O/pyoedPBfJgoD+SlYFUvS4
5U6q/3qGr0jpfxqMp1PgekdFbJ5ty3x/LPg6WAjTrcsl6bmZSZc1Im4UOGxIlgItcYFm9LGW039Z
/EDkHaRlMQbmvpDmYzuNqC13aLITyj+/88zdMpRzTvewzkVYndPgOeK7XS1fPstAeipteR3wBuX1
f9aanvT2KM9HXLPr4d5FJttBvjp4JGh6Oc+aTBabMaMFu+TijBSjj1BoKFwtNiSrC0pF+xjrwUxC
jiyxJCuk/3hZYjDv9aFH/A4ZwGble5TriSRvDJuBbdYjSM7JmE9ff2QoWxlozR95fG5e+ROfZFnb
Ms3SfOLn1gLa1H+kFu47XS6EGylWen5WTHwWrzk3mxpXx9jjY2zp+tuC9CswY8420jtk5nQfRwHS
j8pLo/gkQfoyx/+JNV11nXR/CasK3LUB2LKZAL37RPc0xTIkfQ7/wS69uqu9lTa4lrCS6AACqn5g
tF0rtWahRdC7yDxUiweG+J7dgmlvkHMYz6Z3pqV7B8LbSjrF1/TMnLw1EVK1yN0wwRaVKt9MeQ/J
X9QCngF+i1jQYTbzC4+n/aSFD4ZtTM5yE3pAthrOBmLrEAZ49ghM8x8Dht2adf6+jf8Tkf6WuuIh
jzsSsC1U2oFY88CLYbK1MvJfqBKYvXrSqx0gSyXp2mpJmztnZ/VZKJrJqpSyoyWNPAgYxzznQ/q4
uMSMXtBFm4SpvqFJx4iKyRsE+HEMfnAYe/qcza7CyRC9+516ZMpL6NEZcVOHmwbjXzTc3rswgV5N
XxW4NdH8iHqeTBYc12C0RIpDsb3ggTXF5wYneNAO/IATozY0FW+yOfArXhR0pcHb/SrSKcYkt76v
uu+JdnLSUa+6wGwv2EIbjyRiXdDEoxfh6bd9PTghljiaQjmCpbkoz7pbosZyO8LUkXAb/Gy37Vgg
CUUPwMZGKgC2Al+BbfYw5f2jYGk/oczx7Cyh53dLNRkP4vqp6J9SfZFM95yJR365GbOxjs7D/Np0
SXB0SlrLImNlXp/lU0ecmAv3bwBN9wCYECp4ZXVdzo9IiVulKvvZ2s8UvaKT3JGOST5zokQi7jCy
CrKVkKznxh8LazzWA7s9jx7orYgQCx99mimfuN6UjWRBOodbnQdsnTRTFgq5TuBgj0vpwlKdiw8c
mi9C3avhsPUGH0Jb/8kYopgLlaP2D+xfZ0OT+H1kTM7pzdeM9pOr9RZ59y8szWzO4siUxu56I/pW
tgoh2nbpSqcxyqxBJlUwERQgsJaOrqUyJBmlIBMTfUSU4h5aZdiC31+8//BKpCcztK7MiGVLPThf
/JKTdFjLB6KaWq50P8QyN1lZHGqT4yB41djUHinr0fHCSogL+IimwzmHPrZmpSIGALMry4AVR9Rd
d1B6W1IaYGmdl0N4wftpBLr4T3QCaX2B9q/TsjJFQVo53UmtdFeXYk9mhkf72Djh6zbDzPTYCIPN
4N0mhz/WKwH02bfXuoxfjt83xU0ociFUBUDFD5gWkAZtfCZja/fsiS52yfiMqf/wokEmwD+NB+K5
kfp4usWyvdbXaCcq4mhvsy05Y//I80I/pQbyohZPL89zWeGc/zGH0mIMlk9+IwpmXy1Ucjcg9EbG
Bh2motijM59gYa46yRJFxn9EbU6VygHS/F8FzdIuCCdK97Qfyk9to52sX8jF27ADRW/7mfAukpv/
qBwIIV4qXzCP4pLjRPpC10lMtT0rWKFTEIX9dzxGfplLGSHlGaFj5lrgm8OKmGBJ53I4iELRMFTP
NtSZqeva48e0n67KysjCeejqMkP7Mry4LgKq7P96OlCaN3+BUln24LPULn9y3Lt7kSSXEwVNWEs+
txEp2PzeIiyiM2kdao9701kj/EryMxnrdoK5M2Foxa2/7cMoG50uF2lZ2AX+zjVCXZl6gOXs5W33
kNb1U9TmfQvjUs7LZEpWk7tPbW/5fix+pz/1P9S94UmwAf/XZ9pmqUx5f+1djW/jJ3/xKzz2Migz
MrYHX4KwuYwYReWTGaL1wWqIGB/0lE8nekJ5gfAUkRaXJ6cCAt5xFPvQMvdr3fDu6OF9b/DM1qvL
l7Y5s5kZxoEBCDloSL/n0OZG+m5ZtcuipFZr/IoJMMTnfWpYc3DAyYqbT0iOcdw0+aazeQUKUWiL
B4bABMO6U3tJP0fhLO89nA6szddmrh0i15mQVh5KirkpA0CwFU1h/o0LwDg3WNNYhc0XltPFvtfe
nhLs8p+dwvLIt6v056tlfIP3qDFPhYpvA+gCLDkfCBpgz5d/4Cs5oBbGehmAdn8KDsPzVzIA535f
4HqXOLDAmBi145e1lZcZMkjJHPzFI4pPg8RDAGlqLMImmjQgeI4uS4LVLLOM1BhroJ9K86xfXK24
2UBQryJjc/wH/d1QhLYM1vbY9BGUKNo5oH/c6ESnoJI80KA+AUgdOvLkHzy+76S72vga7XO/ZpCz
AhErAedlfQx7amlUsJR2QAGXPtEHgJK7y6LwnQFfMLOarZxJOW8IUmci8Q5QoWhBvCKyvy8+Mu60
yVqnxx2lp7No6XSUDmlf8JNUvbbtv9iHwGjKkB2LPe7YHWTGORK1nCVGDQHbwjCypq47lFIeYM1+
pKuigX6Cv0e2x7qZkcCXAZ4EIpzIVWcVRQ1Hs2qGpbdjxHCuriHInuH9Kqf4FruHPKuAdNdkkCCL
Lij86pIHF39oncmG3SoC2LJ9yLoXY/U5fSiq1mYKULHkfXsRAJ/6SbZIgLsz2QnnEHQEdYCohp1/
zEKi3Gidhrcy+BVazwFOLvFmAgb+qiMo/j4hp6q67V3CwbLyCOYxUlNzzVPUxZbO1/wQwq2n7Pjx
ki8M48V4InNmuvgJcQFHLJy+2QDiA1NHSaeOT3JfHmpU8DP7ewXZzAcXbM+/QWofc7HL7WLeiPA+
/OsFh/5PhGmvKHNgpXR4P5R9m14MI4kldq03dDic38HcxQmS0I/kCdfKoePo/1JFh0XMUHgKcQtl
cO7eSuqiOHgZtXqeeWfY5H883zYvNDXIKEDZqvwJOpjnMlhtd9nlj6NX5FLWqn/+rLRt0qwh97hp
dz7Fds4ebgFi8Q/UsXV010Iog2FJcQryJgGxCAzkFZo4EwDXyL4Ww7NNh7Qp8HqcbXkAGp0OencZ
5pVqmZdljFAPXfXrRkBUY/m2lW0rzdq8NKJvtXIi6LB6Erq/rSfc5Qz+GyOGxfdJcnevTYUIGizw
67/EfLBIgTBRDs+NKG5z+F94s01BbWwTh3n+0otJMt7TGIVcYqrjeCzjfOdXaYlbei5HlKbiND4P
2GCO1IXYkrFfFWJbNoXwhB5arUcfehGOeliSUE5qDuiT4bwa/Ky2hdYiV+Pbhr+ghGmBmxsdHAVC
W8CkVpPMDpTYAbdH8d2w85eXYe1BipBqKssxXsK5e8syN3m4AnOb+YEF0LNgCk5lOgZEKbmoNZLK
8gWZtaMoyYvwO9vPGHxlE8dJ8kjLCxDLOxkFeTeurKx7WVxbku8AOJwduoEwVa6wsHfVnAKOAXWu
ZiPUUw2WqvQdTybMGOBS3k1AnMynI+ct4bMehWGiYfWWJEwNQSesuwEOm0/ZRbnVURbUzOyWYnSo
Ex5DftbLLkrWGuPkGuzd74gv84xkBNkGlsaX4YlrCzAQe5TV8cVIajDUazSL2lrE8oksJivw/Gm4
3raetHSkGGuuaJTz/gZqM7bViZ8BT8YXLbbI2noEivxVJ0kVpCx857dg7OCKw8qg8xt/Cn0cbehA
wAufENlxb7D2TK01NdfxIjKVoaPzcThkWgQ22iBpoZJ2SaDaUdgjY2fLB1vu+s7p2SjRf1wikREG
kZ4TVmV298r7XtI0Uo0ug1V4FAG6/bpP7O6wve2EuRIy4oONVHbjIvi04A5xVYOCiBTZiKIgZ3Dv
U8ogKd46y6ntbScR4WDT16vl8GHTezZtYXuGcAWZmaGCzxbeeZCXcbjumV6k6u7Tdq7GCe05jRH4
F7fVWOevJpF3OCVzkjwUPMSxSeg55LgHvGItfUHbj4SO9N8bTNdDCHVbkQnSPdQxciYPBygukIDJ
PuObmc+ZHBVKcas7c6txr3b5HM8qIc2D3lOm5vkka0efvEwkpYBvd3b+NqYFMpgubTNW6ILG1/E4
iRwRDdUSoC+3hLBERH81qTeREnDpnWwyT+IR+cTE4j7y9im0BstuT1N95AvxDDDffnVchzNhbh5r
vIjR3yIgmBwHzH2/Na1WjTmkLsOMk26KtO33eJJqF935eLBHvHWc0rvHlOgkKHV7hNjlOAiFrYuN
FdIxBkem2RtBCVca7kG7DCZOdDtWr/ja89Q/ZZCFqgGKA+nEhdIU6bvn31ePhFyuM2glAcxzjOlE
fonOuDHwpaQMX0PTyNvCJhz+zHLR+KPT/WW2ZQvZDQ6NdMouvH2q8ef7V+BpolXKay+7CWPUvBh5
rFRvy31XlpM9boKf2Dneuolc1A1PsTf5P61kJyvszya3MXkZbq+4f813Z8B1EW3F2ryQGSaEjBAl
hM39jGlOfwmfoZx4YM1LjFzuwlmn7r1xa1qUh2noI4yvgobtOZVRq5DDcKhWAIF9zN/pnAqoZ6m0
cWRi+y0k1b2aHPMx9W0khrvjZwlqaU0N0d+7PQu6avJWUpEPQrVOLL5UzsOtVMnBIb1m76Bf3IPV
+8SasX5flFYHqmKNFamVWwnQFNFBTpKnqO81VtMFm9XAvvbdmZeQUCkbKy5wPutGSb7zf0XeP7kZ
MA2D+52yOSIPcUcjbdFfGItxTyQpAa/nvX4+sU1ARuvCyuPaHX0K3egx9PMXCZ4AkP3xH9pNd5+x
eH7VNTbMbb4oux9kP4kYRm3DVa96/G7+P57j3vM5qsXt4A+z1h/jnSkZ/ZCzXH7cglZUV4iIOw3K
EY8b5Ep+DGPZN1hIXt/LoaUwapKnwvI8rvGXO1R3w8LzcaFDkxMgJlprocI7+XjRBeTL4qdsYv/9
4FoE1SUyBTrOG5g84q31TVMSDsacClVzInZt6BPCuToGxtTf20MyxHez2Z4F7JV1bi/C4rpkblcA
vIU6DmOTagqTJvoEXXlOUYw41fzK0tnln0YXa7Mx+gWZ/ei4nsSesWauZv+fVnZdy8w2+cHzhOTk
ITx87gItLc46YuaP9P7LybQcjw+vKbb8NGkTPBbp9b40vGUPR/wu2fdc4aQCwkCl2t0cfzhvTnES
Ezy0cFvBZBW29vS5css2ga85svV0mELZcZRAvKAPRQfwBDxxTf3K7dgIB70sIvBSGFaZKWsWBawE
UXXpYxLmM1h6ZW324RhimSX8uxhB4pS2ID9P8Zvi6agh6wUuFxZuuTpVg2AkJS0IYLLQNL10q8ZA
7u57CZGs46xPy8rzPG04E4555l87o5VSRRc58uoCRjAMvAQ+DeUVM7SZTFV2zpjzUlmYOpDBpBFN
YUt4eogHdorTC9Z3tRsk0mwdHpZWBetbd1+OZEiggr9jcElH6rEBqOIeX/mvm96HB5g6KLWgClos
LIm/HEHFxmrNvQwo6tYX7n6hFLH7FKcf3ST11F3AERvUijHWpDdNrcDpQeg15ldUIQWiEBEwNV/h
uEK5Ejd+f0+m4Fob9mscGxH1a65E1QkC90mYRVkxlk8oOqzlBCw337iWUwnKZGTyEqsF3hq905IO
A1FNISoLkp4Ts4BOUmZEmmi0Ss2n1rnEsy4x2BzMfdveIjf30Xr0c5KCwdF6wTA1LUWLGakaHnF5
ODic1ze702ZpAdJ99qx7Gyj0vSD+9rZLsV0CZuGQAQYAQyxqS3Y/qsORb+A/yq3fFztqYhF/9fVD
j7YCfVZA2aX84hyHQY2u0uLUJcnRZgzHRvjAid/QtpDgOdtB8BHIATIgXEmXNMjfCugUtCpNp27i
zWVPAnn2ntZFXhntP1UnkXIYlcEFwpYAxFpF2gYsOBrInpUX+sjCaYJHX9OeJ8uqgK0KUDJEgWsK
dogYOuLJTqAybwuCz8I4dMcETu9QV6E6MZiqOakvp9gAR/glttdIkGGWtFCK6l5TYtU20aMm2v5Q
9vfZSTd1CDuCUU0shpCYc8S3IiemD7h93f1hEv38jRmvYf+9nJGYaUjQQzPGrO/IUzsWRtziLv4m
FylDWQGJGZ6bPoC05h0pFHvn+mxLXVO14Da8dwtbSVBlGlICSDdlLbmtY0/uKGcuXLx37PeUy+7F
RCZcVCIv0i6/2A4HoEYDRAOT+FojbwP2yQIrpN2ciWTQq0Mgam+SWtT+gw7RIUbRTeXuHOKu1cNz
WRsCt/+S9msUsRFRRnBNHBHMaNPr7fOIv4LKCMQq1SwTD4234bSVeNq8MlQ4BAOkPOecAAtstIRN
HAhvS0jYt6BGY59Q6E4qz5Kvvu6Oo9GI959Z9DFbC10jCpcW/xgoXxQBZ1uqWRgY3ItgRX7cHMwn
BprUOeDScmAyx6kbTHrE7pkN+/2T7jY/+1CJC1i9ADbi+LbKCkV5aSakRBU3i3R/BAZeSCtLGP4X
KeWyxqa+jz5X3jfJI+uKUK3MuxiEM7q3cWugL1hzAa5z2bWjDdqL4LIrycrXPvgCUWk6ccNm/P7N
yVhvfON+cwf2UuOYD7NyiclEM33gfEyUkCz4qQvz8SOFhY7cNEgxuxqCqkreRQ5J/XNuSu7dV9Yg
q1HGXPbyr2VPG3SPti237oU6sp/mBFI32qqR8Sr3pqyln48RbhzG3bQ2l/kUbYsuvC5V90k+Mn1T
ugskh4kAJg3kgvcNW65FleqOJVH+aywVMocTh6T4iBz3cSNMSwkz7/x1tsXmCuo36nTAsQW24kle
1qnI/aWMrsqKL2Td4SrwCnBy8W+jUyg6cqB9LMZrmW4j9ye6tlDGJO0IHGPXyKY7Hg1PSxL6KwWh
TUNwOZHjXTPT1lGEB/7AUDCVcFXhbM7kmGRjYaGQr9i7V8Yzc7vhuuZT+VdhWLAQFau0Nj4ihWqs
obQCx+1h3q4d17GFonAkxGZfNFXPvkzLNGXxRqwL8aywD7vpbBcVitZBDnj6LdzGJ8BrcOWSFSl/
7srTP9jbS1VtlmjjSBX5WL+X3qyH+J+MVE4KLiX3pZoJt9UL+g2OBNLt8BolObyq/xbzyqyQHelu
6ratXuc+6nS/whYkqdrbI08wK9FtEs9etnauE5iKRLI7jzIIhu0ApskEMkoT16/bjeVjArd6erjp
6J4Pblb+2DvmHQLUlrVulMvP+BzyQb9IPFBZen7L0A2KGpAz9TmncdtjmRCsskaNMTlmr958MpWf
2VpYoP7RtrZ3Olo75wTR2sI0hTN6H+vvlIQeBk7R48oT95H7BLiBNeBB4tO0pwQzYJhQdRLkLVUM
DePESyVEfhrTDaN327YgRWSfkqyoWAAWRZ+HmWP143tpqtUO+5dat8jDXi52dpczNOXPGNvKpLyN
CTRrshv1YnndV4cXKFchZj4rtzu+ARqme2cASk06jU5+f9ViiHXz1bSJxSKhT2IDSw1ay6dlt7S/
5KdzxccCfUMCPRACh1keDukOlOK/hiPFxrt72K7+7ccV8yWEtYaXMJnoVo9jUMEb6nHU2QiL/KGf
L5KZqUqAma/8W4LCGbyETsdRwsTQdQ5TfD9xPPztnQOx2v7DOpzL/rpHkEKT+OTwqUPcw47S/7HY
/DzPVohSJKAOVg/vCQVh7AEQG+vn4gAYEAPlaUHXlgQd9M27VHOpILNwNMqdhyk/1DWyMk9JnnES
VaCT4FjfoHarzqFGc505rbIDZd09YEUZVX/kajNvktsQ5Uq/pDZuDFvztMgJ/2isN4Mo1kPvXv6z
KeExdGpObvlmi0YYPMQYscRHsZwill8b880Be2KzZIg5cyNTqQBEqXQzQjZqbXnIGoRJezIv0oGm
COxYwxJaBRlkL/NWlM724w4T/FGA6ZI4MIfOBHoO/ewizdGPA79HNZZeBF/j7Jqaob6kUnQ1GPok
1dB+L7RmDZGrDniQ8ZrwthfE3kMvgvQr4KsdLYVO6Q3XABxWivLRI72WCM7QCCA8CyywY3KneJ0W
TxmgVYFe0WdE8n2riv82fIenNQEMHnnyNgqnpkJs0eCRZMSYsnBlR4/Ss6ARHCFvRoMFBE7AdDy4
Yl1UCotFWqpDm5/vj/ofZkPix+GbHmLG1WfAuhkcQex4krsRIcFc6mFo2+2zC7YD3KjEELFrkysx
eazDsYDRKwXKoW8bxl9L+ahHc9raHnRocpt3ItpojAdk/Spf5znsqL7tvEyHcV0hhG3+oE5UxINU
pfzGAn8rnKvdA4jQoQTlDPHRDKn6iY2dtHeDQODXZm4rXcauAiQILEG0XuiH9tV6KMpHAjUDEmsl
Oe5s+Wbxdlx9R8cNF5gUm42luE4XGcD6fPZZwypN/Qq/QVFWl/BmxovruklbHcgV/may6BsPwIP+
uusgcY/hfuefasH0yvzlufo6/wVSw8YKwaELGVyqRNA+PMckfryqdbqthKUN/8y80RlM/FVvJnZq
akijLRvLyxthHPsp8qi9C/sCl5oe4uuxM+GTF+0gDZQlMES/8GFCU14eq7WaEVD6rGO4AQG6nYBv
2Z2xdqyG4r7i1AJ1za/xsMhT8kDCOaXWLC9CKBcCFjyjfpsvp8vczC7jYM17qo00Mq+Y2yo9/J3u
nN+cwj3bApsb0dkK/XuHFztDUn+DZLMp4AVXfwBCysiO0q4Z3LYpkcvL/TSxd5be9YMWx9QIj0hB
uJjq8d8YMUKSt88v85oaYVJiqiKNlQ8fyGe+01a1m2iDCj0xithZ9cPvIjXnbFToqVWhgTOwOmco
dxZcniP8K0ZBB72Urs1H9wFzGEEO6om76V+71IrHPGUB++raHa93L0I2Zas2dua4FGY027stzI9Q
5YYSdbXJzzbmVu9N0z3S30MzmdxkNGzQS05cG3RtNboGLYaDHFt8vGNAkUrQTBfjPUybGXizyN0C
bgwMbFggtERhiIs/Us75boa6xsBvmFknU7YRyywQjIDHVjDwsRfdGC0Zo3LU0UTUaXF4rNDdPoh6
L/Kw2QT6IAX8hxu+H7zkEeq9Jv1o1DnZyyoyVhZfjBNGowpexBuS08vXwZ7VfzJki7npvNoXAzyg
WWjtf2FfkAqpfqtpVoq/Kta/3bIyc8onksOhoykjsr67eKF3S3/xBjadqlxQhrKx3rWORRLaBUu2
8HddSsSN6fUS6oClfbDAnMAVemndPvkEF9pRHd3KsRdLIU3ufdkipNV3yMe9r9vSFdhFLv52zcqW
XPNlwKpOiXukcco37kZ0zwCdNquinfafGTI3nYRHU12g3Q6mCTEWp1SMpUhDWEXrt3ISQyIN8deR
fLvRAumcuCa797qjVbOHi/0NJpGEFgDocqQhhD3lfBfo9NaE4BxePFKEuxJR/GKnboL7I6acOKaM
+2MbH8O1Yqwx+o/U16OTrmTPvfY5/rPL9Ri/LzqZwgnLVTAlfx+3Nrw+n2050iOADLWYwZ44U3Va
/65+p1gafuraZwYa/0os/VavmpdL2nUf8uNMjCymPGv2ASn3G1Jt6DE9uvfln4SawfPFntUPrBcD
QKIJRHZGNPj8d26mQ27E/p2PpNp2h0+9wMzdhnNn0eZs0iJtj4gPIVO9MDWJChLHFNMjaAarM/ZX
joFdKW4WY1G5jQa/gSk6vZHmRXG1SuMGINpPb8dw+c4kCoTA99rDNyR6zRldkYgkVCoQFlh1Tjqx
Spt6kRKVpQjGrVT9Vui+HDZzjE7gxddLQwiT7iaA1tDh25H1FDEtoPlMj/5dFwAUsl3CfRy8Lj8C
6NFDnrvrEeLUnPERTQo1yliSpEB4gYgH34XX7r3/I67o3HzGLHPnMJlpchSzoRa6B8W9tdKrRYOV
nOEepgr6u9rv1CCID7YOs6M8ET6d0dWE/1PH9HmdiFmKRbNPJohjsk4mzQE9Mtkq1H7GH91Ysk8l
e00VUiioEUxlxV3ppzKHmFlEFd/mvy2folUxBrGpeDt7XI9bf31pZmg6eNYFr0VYaFiO5RtGeDQY
Ndl7TaqbwxugO9TPDrikE/XC/KcNxeuXtg3yi7QMjIMish3yzFZ1UGyHR7NdSse1oGAH3GhvZivF
us39+bWpYSM6jeFeTw23JTDYCMDXKBEYyidu2jq+d5lM4aMlrHdbnb0SnkqSyGtw+XZ9stKGMUNb
uXfJ3J3loRmMSEizmjhjHkzg81yAJM3zwL4kDU2tK3ZrED+Ec2joAhRDFkeHWpLesHTl27CLsqc+
rK0ohHGcmtef/dhA2WdbHoq7CR60FL5Kz8qZHuC3A/c783XrXmTs9grz9f/rm2ZduN6DSlHcQQx1
xF0mjxVcqZ3JyzNdhdgDwj9i/+GfZMiWXF4Pgrn/ukZng50WnyOr94v0qSReFct9oZjcagr1HOXW
Lf6AcHEN1Le+oSGc+RrTaJRVald1biGwS5j18qcM8xz6uhhXe6Dx5L5rcbcmt8keLeO84mY20VZx
lSGJPGRuT/SrMG8ueRIbIS+2I2dAmO1yvCsSS4E7w1Am5RHC620UhsFRqJr/ObDEabg4e1iKMYDn
qy/j92JpxxzptOVLCSLlXgbC8cEVkZVh4XObgW/xJnjZ3HZeHRwHjAEySw4jFPTC/rmaibxMajeI
z3V9Gi5R71p58iC2TBc4Ri4mSGBL3BxP0A42JZhP3pyuiYlzqXBHNF1ac6Ew90v+bNrQsGDTTNYf
43IIM0uih9hXETZyr5KewtDTeYwJ7ZXZEFWLjoxT/Titot/IEQfQ7Fop8RLobMrLLyXZ8nYvyYjv
HIeSjWCNwAen7Exikh9Ixs1Du2V/AV6+oI+5dhmCJCrLUI1zGNHCQIJ18b0C3P9UNzqx4goDtkPD
fyvE6jJ76ZwyLglOalgrcno4g8+4s47z6vRr41oVwC3hjiSIpD2U7UXD5cBbvbXgYSNzpuqP5QD2
eOpnUq2t4mxsPnbtnQnD1PkJMkpRII5mHEysRggXvmw6ap+NTyn0V0RHYlUeMtCd7aHyigKqW8pg
uCxEhUyh84DaOaS+oPrzyhML6KvrwUp3Cy03xq0DYUAnIBWNtM/he+5+odgPiKEUvzoiUtxItbKC
FGfpNVSKWpWp2wGgFJVAqApVglrCTwIc7kELZg2fThb1AUY+T60MqYq1WdiQZ/liVCwcCZQzlU5Y
sRUsB4OrZPTrcH+yDUSSqGtWmmyj/yo3bzYlHNr3WUiO9WolVcscBWpurk6EsWhE40NLyOhP6+aJ
qWfgwR5XNDov/qkINrf3BCb9B10P/xSlWhAQiWl0FkvHMWAEdhfp+10YJOUtafsK3Tf62SyZYw2I
/6MH/wcgyRwPpv0MkruVrUu0LSOhleEtC1yYzFCkQN4VoM8wSO/WFp9G4e4c8hYoedCXo5Y6SR5a
E/QWqTsFPC1n6CTBjFuRn7QM0QzKvhJi6JtX7IQvSKOLYxoyBg9qUGbq0nYHv6lsi2CKLjv6ug8q
/ZSwBH5atFbtk3gxEtbtqtcXyZpOo6giq8syXwfBd4y+cIJ9XABvWIWUtvUDzY+JxJYXbcA448ys
Uc9S9/39uAsxDXFoCpSSkndUA5VewWYlJllcao8AU/OBj0oKFpb60RFX9wPJ5PEnetNqtwxtkUMT
ydeXO7aaCUEI8jLBc8XouFN33FPfi4CEnjSv04lhd09RHGj0mGE5t1UNmhzarCJ25RBoVzMbBt/O
ZyE2610WIf1qQc+BbpVygC0wVj8ev0IPOfPk827dtX3/bkmiongtqrSrikMcUy2Y62/7oQ2IrzVl
Q520Fw3EyrvXcdt1t0oKmLSHH5FYJ9W9Pv/iU+SvatZA9Zj5/vizXYxIm4pkMxNLg5/qQqBjoTaT
G6siauR0T7yLUHAZK6dPrf6aLRB2GBCjQYQUNneeepRDTbaoX3tAtBCAp1f9TMNsWjfba8fiDWIh
MRA7u5rp5/eGzMWF4mY5nHSv8iKsqaUFOYyfoI3ELrx+btKT9Hf3jq3OkiTWomriGS3i4htt4JnW
2Cuz8o6lk9oe+gy3kNVxKmji/O1Qy8ZqAG5J6o7E5bcq3Xmr56FgmTv23vQFsRktEGETtjvNAjRU
08a7Etq8MYjKwMN/AvyTKQ3SsZBAAHCE7427f/l3q5jOt76P9b9Rl1D4gkB7pUk4VCuI2B6oHOZa
0YFiDCNsaRuf8Mlq6wpAomWfCjhoAv0XD/G3mowZCJhk4zeiQc2xdudoi2013LjZSWIPSEhu815y
RdzdCpQxqCVxuVyIEW8fAUbECa39y+DURVnOQKKbL3B8Wvtpm0+JiGCsNX38+XO5BVGNjlBlj1Qb
uujwJcjlynoaim7n0T2tfhfB97viiZEskqx85T59M8VbYuqoVIA+hRnfXlvJtE04/UclntWMKxNF
TePKlTYsctFxZHsoMYO6jInJcOxblS1Y97kSK/qc3O4JqNSlLQZpaIqsg62ewXV+psDaPRbQGV+K
dBqPiMgmDhRfe+CJFA4hsySwHKnv2gfZ2/1SClK6ceEhYz1gjojh2pYBHo/yB2rM2YkjZQ4DRJbR
Dh/Ny7iIrcY7i8MasDI/VPj1lvcbx/YwYw8MpR+w/84DtWqpzEj7hWvDEybQucD8WmeuS872X9ty
IUV/7PZsZUlQbUqANSZADjDJWGu1dXaVmlWZLw4VDnUhox+I06oKQVvG0TvSjMGjLPImnloMoNPo
GbM6hQbHCoJZ/91XiOkysvikA4WzVx8QM/zPu/hShPVZC1YJTpN7xOYIdSIROoIiZLorye9vRD5e
4sgEJ6OxlnUDKidF9hMILRwTaj95IU65V2IRCLByALuYGqR95TSbeyscRrIdnC+Nn6Sg0Wx5rq5h
GcHbG4Yq8xmjfJ2KngLCVsHpyPe7xB1UogpEdtQrmR4G0GBxu0V0uMa6KIpCtDnASxqiq/rgdqJX
rmcjkDmSG69wSvpP6vEbcUaWTIkF6Em/0/p5H3Ze57/fOud5cCSfMkmpQCu6pLIsg0+ky5n7XP1F
kn20xKFbGN31Zyai5/2p+I/IVoiRbyCPSezmhwMi9F2xh+zSEQevAaSRMkkyj3aRzqJ1b9JJa4lp
KXbY9sMPWLhuqZfELjIRlceKp9MOoCf1eF1bezxId7UikJNulFi0cKRmQ/wZKuiMaGI1TMjS+Esd
NcO6+DbQMrTbcDGHHqkLQApNtHEYSgPlZCCKyqhWjPi4SQv+lapyzaSe8UxvYCgDKQDkJGGBnCLk
4YSIraZXJLLQMLSHTvMLuCKez5bZNVTy5thIcJn+HAf8hJ0Cpqh3RzSfi17vAw/W4KqybdRaEppS
kjxH2CdyvTDCJPSVDF2lHVEqV3uNvkpfdg/THQKoRKpaji7PJvud8/Vl1fg8mr8fY77Mjlezz9J2
qWzxTuH/HekpJU1TZ+4txTXjXgMRlzeHptCe0VZEMlG5xDZKq6lqLnmCsvaQMpq3Z81MeNhtam05
WWg9tPwkTKzmWHbttY9CmLk4dMKCenZ/skVwwhDpKRWQywYOQnCg5hhmwYAxaGXrwUVCbmT5oWpy
PXT1tBz+yyvwmDFTmASEkqU+dISxFH0FxMsRl8VimsZ78BpyuBohA/oXHCoKA9ggCrYlX01ACSoi
mY9xdhUddm2ZMCc8sAyvPbl6JwEGWT61UYvILRaAYyt0cejGu33ETOnERGJpb/+GIc508Xt24cn+
i//x9f2Pajd8UL5LF0rGTDjZryyvIuJg2o1v4SgChMMKulRO5tioazLw5o8b1XhkPopKMuT1p8jB
D+U7S31RBqdsBztq8TQVhCPKzu2319cZAaacVu6Wj59J6hgOM1BTBUGPZ75PkpFHyca71nIr+bnh
KTQkOeNYZbrZjs1yExw9PsB0DaBLTjAHPXZXu8/YxZeSr2Zdsh2O1itnQjauQdnq4ZvdyVFzv5m5
JbwBvxqDBF11aIuBAlE2W6itXdGS6ToadybM8Y66iKuXBcbzI2guAIg67tNyZVMx9po4M54Qywym
JoRl7t/ICkQOSM5DczVeIjLL/61OtEbM+E47w6trvjKrDdaqvdq6oLP0g1zQgQ0BArxjAeMy0E8w
l3M2zM3rFsmp2ozGWm5paMmxjF4AMgPSpdc5x+fBAe0dqtO24BVze8ZhCFlM6vviruPM05s5viHR
ul96OpblJpyHixq2BZri0gX4Bs2QtFVRyZrqCsqsjbfxYu+Kc1/04AGsyjhxMjuL1ysPQTxtpOf/
eXHb/ioi6wM5AqaR8EFhz7bN5xx1/kut/4XG6ihaM4OD/8DQagngypD7FzzpXfnXqw7Xrz5UdeEw
zvWk6j9Gv2K1Ydek3ioRbboO3RVQxrF4EMDfUXU6MdobPzK6yXfh0SLRYf4/4sMw/1HxHGXsXWjT
LWGLuC5K39LNw1/riqIU3TegBoTWzRq1DtDggXEEQpRKhoTaG0voleYaQmQPXmoX8a2LHjQGwIg2
1fkqLEVpbxxeq+jHcmzcTvgUNxLOgSbCh7cxf42PkxCA2Lj5jQlyrIRePU9skuUu52DaJhtivUkr
0io37oZ4Y8enZJiGHjIMo1fQ883/GnuC4b4rooTOUAkNxJgjrtMVVmXycesQOZgy68MIyMlYdnOz
qxfi14i40sAJMwHmfHQ0udMjrFpsbKS+F1QlV4tzqlyoqMKVJ7VkKhVlKiNBKBg8Fx1EkuEdS+zF
kbZnXSa6UFSi80IzjJqC2YDdm+e2qAXZ8O0suyun0kER9uD+vhE/SDWF1PitLV2IE0c+X9nt63VC
46iMk2PLJS+07y8SIueSrvqDBCi6Bo9fr2A8uhlOFDGj1PKsYyAxxPK9nREMDbpNm56j6itlZLtd
f5XCWzjxsgbZUDu3irgsOWBYOVSPWFZMMnIqm/Gb8MOr5Rigw2aruH7OI5YmqMGy02ZjVBPDT0Zj
9Xr0P14BBOxrFNOY6SM8jDtY0DMjUSL0atKv9lp7rJaymMFFAspeWoTy1+ClGZEU/OOL/FJyiatl
HXJdAQto3ozv83I0tMGzg/ffHHGEAz5fFtluuyAhrsvzK/ObhHtIffRkXVEIpuKhhKTHdCm2eAUf
DrFj09/uQAJ8utVGJ+wKwfYJaEspBpTirtBA6HZKVMElABC76URlwUsIB8hPXObilYdw/q2/RbbM
er0uWQsaXN0SAcRXOxdEkw6NQeNmiakRgsYK9wxrH7RpMrt2n5xN/3pcoyHI1qt6sjHt6wzqnrq6
Snq1lkWVwB6Gy1MfkVEw6pT5OMvASor4uMJ6BWEmPLBkw5bD4DC4BNj7WaZQgBYFjlhWA7SNEtHS
KP5IQuPaHJpA5RM+y7avQIJGAIAOGwZWin8JYa6gdRIKM2bieWUgUlQQDnBPHyqNRGPARFCm3bmZ
GFgzX3bv1i7pg8IYMIFqQxb+wh7N7K7oqTgeFkk8Fc9f8ho+g7eYm5dEcmHW13YQ+Hym0IgDFBE8
R8F9zS+5AMeKF/eUKI70z54prU4uD1op4e9eAKT2wORFJkRWyQgIMADcGHBO3UhRY8m6cE4ouj2L
eGMuMG9aXNXcyeQ13O4jnig0tIF1rz/HUfZ3uZZAwFg+c1+AYEWHTWaHr+WDykiMn9pntGx/8pTW
/wS2iThpZ1JkCV5OR5QTs7fK3RRjZ7OS2ODXKJNlmd9ZoI8y4HDAGzzIUM04WwDUoldCZzfzwfK1
tHA4fRWG5Hq3Cyd5qB40up8gjL5CMG43aT5X8g59hveidqFItcoacScyOWdq2FBLjaOseHXrjDbF
MACJzm9HgAsy/TpXi3rzBoXzJ5QBDd7jpNnSbHf1D8nFleZoHYtQp107ZRx9y1FJoohyX0Kv872p
L2gGFxaNc8q5BPPC3mgrWIKlGH8am0UDbR6bgs8UgL3NwIneRKiDC9x84XHhzHo3/mWgFGRT6Uwg
WpRCasALrGcrJsxjBKIHBPmpmJqTwfmTeO6XOoN0R5b+tWKvTG1HYKKckrtSG9DARPRn1M+eOyXf
ziYXXFj55VpRJcWrTuqluzmjHdHg7AxQMGi38MYzpQ6QCW/W2G/s7A+N+GsWfq8CQmk70nCI1rit
NhKTgYCspa6l6/+n1ZaRPcpSAC4NrnSFMvM/yCBgrT/w0+4D+UaNtAwqo7Bi+C6lZJstNShtMx1f
qdbe5jPvIH+sz+bqUFPNfIpM1kJfQ7GfscgKCNhat9HF5dvNrCUQhkTZ9ZWXhjA2c3PDxA7+d8Eu
5fYuvb8az6gA768IhKmUKvketNYuF0dNmOeVicKQ73TD4eYlkprFVqrj4VYOoaiDPMZYcxDHAWVj
ay1Gp8xsGWk+ujFYrIjSL59GGjA5EO/0tedZU+DzWBSKSfTGOjkTyGg2Gg+TWGELd8+ddncVXC50
qSwOaIsHoctZSYvXxhGAA9B6ti6DW9/dwueC08rBIuhG02Ua85WgcYnO5bfMmdHg7EQ7nQx6+bdG
7VfsTS4KVgmIs2Bg9QNs3yc8GErJ4XpXHOvm/ZVLjNoQyu6e2/U1PDmilpkgjbrsRokDgBuyK82s
jU5GXRtyfpmlo77ad4UUGbIrLLqbueVZknkJOamxWi1xcMaNc6UdXrQgkOv6P+aYC5spdacnJ41K
UHgL6dJYohvkhJcvCHmhnROI75xeQuaVntUTbDm8y5UtRofHGgLsmbPXtTf3SQv8jnGG0k4x17vu
RKkWZRGh+0Q9h3S9Df4HxndNnCVYJodCc/tRe+vqtIcgqVXnCsaVyvqoClTCpCYXZ/tJuzewgAAc
NyubKp1o9QaOi0eNNwK/kf6lITHFGB31KlR7R1I/erwwu7mMQj0Qk+mMQvx+rJCHfSaLtVU41yqp
gtn5Dmp/MfsTKqqE76dJbtO2G/nAhYtXVRt1/06+7VpS9OjH87vxU0sq/dG8sPCLzGZffRQD6GYn
8p2nnqhDJSsO5fu9vuGevwSCqSw6rAMZcOfX6jmLRq7RJW3QCC7RRqC7sCQSII8pQXlNqdI8IwTe
MTdnEB6ZnOndfL3ktWoTxiBHiBD2FRG58rfXsUwMEpqf8FCruKBoW5rJR4AfBnO5PxUTWmfiwFsR
Dan95tsVZ1U8UFqiOvESyhS9xGMJ+sQqADj6ziISgez3yOxKhEF3ztP0WcOrMg7FhkKwi0QuQYHE
VNcU/aWRe9x/KbKtm8MUdwmdRzhQ1NsiVfH/D7ftVNCBBRdWrNsY8LLNM9Bi8DU54tGlS2FpvtFp
09uaeKBmZ8SRTYhzVLDxu8y+PcYz6cm9syLG9y1xbhe9h8dqXdxh2/SLkrtVz/DOux8cnsBuvzqf
ocI3jPR7RRcr5t5P0cKMGzh0fd8zH1OIovJn9EqSWY8kD/2Fd7QJPf+biikJ/rqfI3ZIJ03fOAOT
CjVmC5hOMMKhMsbQqdW/b+D+tcqEDjaOZIQBm6NmIZL2OZfFVt9fm0/kiIm4d0oGjZRGmoEe5xP9
7KmlZhbLU3mJuwS+lz2c4nypyFFsuMGloqCdpjRG+LJDsPnAt0anT0/sGu2mu/RNki+jCSrsv+nN
UrXXeffoqflcoQ/iUZS+xGGak1hAJ218Jvzso8w2CiXFpIFiYCcil215mEQFIcX2Jx2l4ERKmiS/
MtflDCGg3riZFOhA+gZmZdeRZmbjfOLrRh4SVBtt67LSvKT29eV7qVI2EMzBabYzT17a4dvzh7ZM
C9CaNzi91ceKEPVIr0pdHWPYxCfylXqcDjAulKuwQzhHBTfAljwcK4AIige89KxqnVOkv0RusGKK
Dke5EHAtU3bfqRNPnnq2GLcoriB31Ha1frSWqkwOF9O0qsEJJIO8SZ7jKFZLfw//9oqunK3e6j8B
4dY/Y6BEUmH0BVLSE2b0YK2Wv7tXs68zfJdWaCwJ5oxvgs92ocgonR2Z6ZBYpTYFDE2UIblQgiwJ
LJIreqAxwd5BQvt6qG4lqgMjkhJNB2jTKUG6WiZ4mIwsHjcw1ZA6TdApNcGGQ7TODOxXTEC0qNZO
EqHhWpayEqob+shfAinO8xkObV6I5qs8ns0oTE+2YepvUCq0wfHE70vRayJXZwEOlqfvezn+5Yra
/DblDx/6Ua9u3xpBOpKZ+v/pfusv1Bvd1/oS5UxuEv2TI9xGjSW2WgCDbXNGmd1tFDBHbLBPFM2U
5+B22PNnyJD7DgqTrmT+H/Uld60Uz9IXIeNgPjhxpV6LyQID1FCpuY71ez87pbVo9ROHZLQYvlkF
gZKuUBdaQFvWm86XPwsqxHgi3TCC4quX0OGXOKmPEFaofQMCkUSsEWJn5cSPHMA9kdDhtp70Dycx
X4cVmaqlGX0dTjbA3KAf2Vx3P+Qxi/0yhe5XC4mm04Puqb+Pa1Rw4Ltli1LIl1t22aWo07momXIN
JP5QdXiy1oA1lGA0jakVqcAPUUhqkE889mgR3BZl2qUTU0tJU7xen6kAf/ujEyJaSTZmGcAYuzoL
1x9zGfFS/AEIR6oI3fAr/ymaUS73iVa4twGASurtSy6Hrgii4YV/f18gQfn798OVHQi8RbeSyBK+
m57vg+0a103URW8rDajYkbdLnApU43a+6JPlGwbqobyuKER9BF6dpkGqVdAh2cx/GThyPKNod/3C
thbvvm90alx2+zmIxjBTSkc0cikE6nZVRcE1BXwTfqsJ77ho4uh4CCz9oPkbhcV50GgHevCMAHlR
urq1/hx/Z6lJs5mxnsR6SBgGZFP+IKASBcZorJvKaR+uej8CE9jHYiX3MJlbjrJLgwhf41s/IoI0
rgHEVkixeK+oSEvUrVKM8TOif4uo2Vl7wZ0fSiHvZNF2u05ym6tZ/ZtclCVTW+2tqrkR6hL4HckS
kyG9SAe3zGROmMNsCzywxFepocSWyPdapa6g07S/ce6J20CKDuM1zjIbCPRb2ZmU/L8Rklp4g5Zp
sVbNDR7bvMUt6JDxCI/uE/ld8TZqfjwF6gI8ZSXNNOgkSB4LD5BSeb+1Q2w3J3PFKccl+1XmzkFR
dds0tXiAP6wkWdlSCDm0+gVuraJMy7MQWC+NxRvTN7VogiFUFVMFBBXPdUWOhAKx0Yo6e/pTISNp
GmITPvh6YTurPREcBX4ECfgC5J/2UKSxE17W7BwOlsE05Y6kM4bEZnJKmdqZURVySqTWyyc5EE4G
sEXUC9rpk1YllJfgPo/g/xFkPJ4TK9gbKypG8cBBwO38nU+Gs9511v3JL1Vq0H8IiqdYKXnQOzm+
S3yiVIkEbiH/qVsvTwCelk8D/ANdLEvLWut2Gt/KKQrvfdAJIyQxEN22lE/Cx8nf9zTGOOT/O2R2
HjMfmAG3+mjkbWO2L2oVVcb+CK7SKrb3Bxc/9bnxOZVqStpUC26IGut+d6X3XNqAvnZ1DzPsNeey
iZXZ2e8ztgym3XKIj7DHA/HCkcwVr9emxcAWu6+kgylKJIm2nW3uX59LSD8EuW9wC/3W4Yw1F0Of
DXfAts4NNQXbAYfiEjRk4VVGyAch4RQZ65NdORacCiP9AC1rXIBihtoJc3K5HG75Egp6MOm7MDw4
n7i+dDu56wT2KHhjvHO56m7203AiC/CVcHCKLDnFxuKPmGk5HS9VZO89pm+ximvkuB24FP13mlNI
iQv3FUmT63jNN00IG151mB1SyD4rZS9Y7SeSYUve4u2mVp/XPyEcgB5pmF/zl3FQJS7U5CwhRq2s
BEBiyRsf7d2Xo4QlxaJbh5uMxpCiTFPCCmli9U9xWaY5VDVLeEKz/uB4nTm9hY2lROCr54tgEKZ4
vAdIWVXjiWAYIdkIr4p5IE1ee+yEGqHg0bOtrmS2g6Bs6mIxR97ceKO1A+dzTHYWec0Srh1Pnvii
LzSywVZ4lmVl4Lnq5yF1h+vxeSGdKn04TLWNMmlsOMZa46s4lItvO6VZDPOlg9Ofq6Eioc4UUpV8
sectzlpu5mcrGV/Y+I26a0SDjJ5MqQ3ktnuG99dKgN/oB92TcHcDn/HeYb2FJTveR1yfkNk0Zo6g
dVH5M2jEIVbzCtGaSkFK+2HyFTEXBxsuN+EB3qk3Fub0FeulNkbIlTRWiyLXWwmYPl1PCOWdvIjP
8LOoAuCtpGZAzcmQdlUIPBVGIJBM/7rcEJvupxM8JoerTijbCsKVnE5rWB4PXYRm1fuby1m47wNl
El9hLvHgAIuOKl94erOl0b7GqgGMC5YUPOEMUQxwLORBeqWb4qls+8Kg61jX5UzRsRYUVU2IsZlX
byOMzQLYw+XRgTEPxo69gDNVkU0s7ZbtFFxB/bsrSLj0HjGaUruOtZogFI5axWazLf2S/7HFyGmG
e5eOpsPYqoK0/0ie0my4+uIN7Q1vyhlu8Yju49Q8rl5LgEjI+cIJtSXOexrL/W1RhpEtAwCdgpTE
JJhVQFFSzT+VBuiVODs9ew0CmPN2VI0/HiGmOcB0cprDa9CPtSTh8vzsMKBR0vvA0t9w+vgoVvMD
5e/4tCOUSy94fmvzcIxkTvEHQkcgiBiOPIebreyXWpgEVEqr3Nvy06yk9RnOVMa1/CtJ+4W7s+uQ
HpCa6j703gP2m777ZAsRFkYHDnqayRor/ohpFUfjp6ANHuOs+XjlBphOruCfnfU6OLIx2J0Qecbw
trWO2ks0gUWKOyjIK7bdT6Iq/+Bo+BqhklVW1vkMkk6aRXPTkTNuwHLWSnj9ix+uvbgPotNl3MMO
yN/fUSJJnhvk1IYyJIduvJizgxl6PFTFWKOzQDCO062uZy9MbjExcfWVEBzoFTn8iKjPm4XBq5TI
+sNIDVGxdwqZ/b/5SUC6cEoRZnvNvVd6H6HOC1W80hpM+Vk1tFZzqDMOJo3NBwdefOPM5yaNQqQk
5giDhGo8eu6+iZY0BaNcoah3na69lw/qX7KPYbrx3FD54X3ZN+4FTtlS5LcIQ96vpPpy17pLkI7i
8Y2D2bKLSGqOBl3jRaNS4Z8c6IgHe8OZK+tCQoJG3C/hf89/4bmsjP2wLRopdlVTan722Afzl1wP
lKud/gvvEmp9kcXNmj95zVx1SA9mG2VDtZybmg4ZFMGBBt0V7bIUeCtGPOx1lSZuZHisOMExIwLt
YlRh2GW923lkf6v9WuJfVe2cuVyizel9trRxkj9RqwOe7YYZoE9AsgjSQx6vuA22BW72O0aBuies
lSrxS+ybMIospF+ENsRgV8fMEV4gwU7JbqYe1/YNa8ZwvUB3RBSGW5fTD1DLFXIJb2ulKAP5E8w/
9uXihDgUcYEFvAnONJn8pRP27mwCTx1cn+hcveT34ireFTVHW0oeVr7qUdcBkn3cxqBrqvlrYOvB
+t15XeRROyGwNOgRgutXCJWm/wjwD9HhxpEQ5VuHUw7yges09lXj2MMN0jTqV21PUoKY3IHlV5sh
IlMyWVyxisKK+YE0n4ukxum1LeqRiwED/8NGopTWJUBBtSLRRra8lwG+zdBPChKkHwru+Ja+Ubgr
ve5hjCTanqFSVl32MAYrGlzGLjR8AJ50YB9aTXoUTchE8Fs4acwwykkOlkxlBLlH20PGWRykDvwm
hsQZI3OWPRC8wayjd3KAkIqC2sGHoDpfpZSz+8JO1VeYM6e5ouCXoMyfmrQ7jS+Rv5S03AhYvJ9H
B5sUHr4YlnZPVQ4cavZHZt5/RUeoiDZkbqj20wsA01oAmMvDKI8lBS/+R3+VeqaZSgun5xYyuCve
YOjYRq9KxTgibFZyKaryAU067dezv5SBfrW78EQbr0GnhambUXbrfU6D0cfDhsdeTBDL/ujzjost
OoatVFlGux+Gj8a0Ykk1NBJMyLYl/0Xy/oDmRatodFAcYZteTTaqMP0deDBGBUVgZuRAE/RzePWu
hUIif8kCk0HxZuHvO9u7FhIp6gk6+6+yV1NRWpyldmati2dfH0jZJaoUx7vltQCF/+/PQYDf1dNU
S/ML2SMF1Ufga29ORf8XKljeEbH2WkA2qJMd6X+kyhZJlNDNMYfAMiev4zDsKPqaieoenyXA7x4E
wEDfObopN0m9qjyk0muAPcyyS/gDUkEfe2cYXjrrD4wCEyoWYrN85Nl5Mgkqe1tA7mID1S02a1Xq
8atCLYShWIs0TjquZ3NoF1ZTyFah2QAUI2ICttABTsMjGiDfNe0/CX2KSiTixtT9y9hWyG/+ZyQo
YzsJKh7eJgpWl0fKxqKpC8N7rCYZ7/x7EUXXYE6hxip6YiE8993J565GFz1rfSj/fFsk6H1Asg/8
alL9W0BtJypphXrV/KTl+KPCZE+JHIwM66Og7SS+mb1XmrbXKlBYOBSkh7r2DiAgoAYzI58ECyg0
AW2e2dbyOEDzqabLG/RV0/+cW6nvH5HXdc9SqvPhanAPn/00WHvfFJTyhnUAG63NV1w1/xXJmCUK
PE+7jhf3yU0Cqw5taf9iBFpzSMrVlHe2F+9lhEyvFSUUalTFPEZSCPJZprYajJNlYrJ+o1OBnpd4
2gwR9Nl+P1JvthIE1ny8BL3hRa6H1K3hTgUkzWBPXw731gPidzpljtvGW3ouH+FtmcQoamEnQ/Od
fwqKxqiHVG7RAswkRnw9jj57Iaamfm89Je1g0HI+ewQB9lm/cT33i2uNQ/aPPXum6ix2LgRbkYIJ
dgmkw5s/4+Ymoxd9tuAGWCAdgtxjjwt0DL9S6RPFi9G3ML7UywYIRc7YcozVlznY+rrgy8oOPy4g
liqZzIE9+7wXcuGEVLphWboDva2sa44TDw28Z1tqTWb/qZhHMallD0oC9dIl+8e5fkU/5Pd8IQ4b
lA7nHMXPX0XcUGDQXdAuuRF6IBoMiKQoBz8WsbPRsS6rE6Z8BHAqXuuXDRDMBt1F2FB5quch7sCv
UIznuIGrGPnQxgrSXNm7HP1NLQvAWITukKfOk1/UuJl4T2PvTE+KMMUKc+45Sv2VCeU6zPvghHka
grwWS9Pxexe0zntb1hFmMMyb+nJO59bQkAhVx6N6qtlzfNLty1A67zLcgxWgbkMPUV59XoQmpRtv
ezGoP7/RzO1CgmmwpekDiAisXdJaEfJomCbkDv7SA2MXLQwaCCgsPw7q6VntNyOz7HEN+EjLrtk7
L55E7QmN5yWSikb2YK1qhLYJnQ9Bbn6kvTBDvyJVUMJShK7WvlTTSZd6p2Hc3aYg6dztF4VpB+7h
XLPSbxDYNXVkYM6YavaEr9L9L3Ft+XjZjZEzW1YnmRuEBotFikjrIQpYjDbNQdr3bWBIupY9+4uo
VSHo1V5vN7BjATsCJYbpsz5cUa81lErTPXRvnt8d825pD8SWnF8dOUgwttS54u6AWWFBjzRP7UGm
u+ZIBqtz3ZT6IsR8DJDXQRfZ/DHkWJ1ZqkWu2frTrnGUF0VYEO50QtBkJDMuyNscKiJHxZneK55S
sEc/okMonTigIjS6LTBik78diK5mPeefPc5elte7bimiC8Ct3zwSKikNoCrwGedkPYf3vCdjBRn6
tfyYEOLr6LWYm3t3DcbRINPj6l/lC5Gl3j3sQUZuDwIlOymAU1Goqj4PKM9uN28wKrYtk/MxSHO4
7ziUYSFaMrs6+hDvPYXeT70I01WwP0LuAOxLiHM5TDpAUUTR13COc+iIDsGLiZmDELYRBFtOzN7E
bjzNhSRJ07AHCL7E97fvCBc6ltrn6AbvUCfivD5+3006YeYhdG4cyoC02Fbw0EPgpCSYjoK+JrmH
B6cysJeT0O3/ovrCwkPK8+xAPkOf8CyJzeWkFGNlL9HXTsJ15NlF5UIP25y6lmRwM1YSUvXI/6QD
LI/6T13Blz27HgYFaX+wxWmDPhvWVn+196dxuoGHBlOLLB9F/I08NVu4Qu8avaG9qGzut0EBk6Ji
pnc662USg5W7zhJb7l8bz0uV+McDk/UTD0cz25jUKt2xGXeEDgOErdaI9fvmlaTkXpu1Q5RtRL7t
dRyUVm9+hgZF61tqATQYBqfgLj2bsi1hTHNns0JGxTbk/Rty6WSqMPsGM2POUPfQlT8bh1GdzCBw
5sELnt6Hy2qwXoaskH2rOQDJbHX/pH+nh6gq5v7L0MVF9v05UXsscZU0AV5gV1kAGn0Plr2+TEhl
YLSoYAV3ZWtkL/NB+7ZdRh+4/N7Vxze32X0x8HUI5U0dd8OF5wJiCSgujEiRF/MmbPe0Evx6dgw9
XUgLqetQmimb4+2XkvUGhOng2zSgJ3llitFEodfVkZM7kaU1Ptei/is4QW8WFtQKSfpuTpDJpmJ2
5n9uvMvppnygh8Y5b0tGY8qK0BREDkhGIghHiI4oyx3mdHCZ795C6UepKtxxfDbHFX+YuLuE1INi
1BkwnTYBexrgUONcqXPbjxtr5dxv2Y7o/vyMphBdH4D3oXGxp7pmmq9rzTWlXRjOJjvciMU0cecc
tdJguUPqKchALisfTJaMYDhPTAHTkqn07P1tXOylpWDNiinAEMw65qQxeiB/MXb1LuFzGcencBgx
HfYeNCARLLrXGomCNvZCFjEFYv5kCyQF9dUhTnfplN/z5Kdto4zhQKrBPxyqsPrG2Lq+Tx/dRc6s
Y5jqLqfTV3xNlJBDYoi+i7WcjGEHuZcgrLKovcjHep3dpPEnHd9vEoM/shbPkO12tKOVqxJMhDf8
cPklWuaB5Y+jjbZT7Np7HZZ/LxvGjaip3V2o+M+7Qsj4kQ8yHNTelm0oh5Vlnj912676PV62qG+Y
lgetVgOPAMZjOI3zUpoXwPJ/sQ+kJsZGQ/KCfDPHQGtLpiyEg2FcPctp+l+uIxQdk7m3cnxs7SJb
eDt0ncaouHh08MscyNBOvVpxYCChFPorawM8sSjLhKx/XikoEocB+gZMW3adDSGcOsQEY25EIKW3
U+9MaMHnyKK2x6qz6YLazsyQ5CLu3kEBP+kSkF9vdqm6IjlnkopWSRgy9gV6pxiYWVkYq9kOz/vf
3NuYECOmmfsOV6HNmSohgJr6gtsKdHr6b9Yy94960zb4dFDxzXApnXdjwWdASQGSiHrgbqDayasz
oxqpeHPUFsVX/dWNLUwtlE8Xr/AtVt0y1+zWyftahzwnjsQJH4a7+QEQmYMLmqke9mH/Q4zyUCzT
wS92y+x/ER/Da6n5T5DYEWE593imNwQVRbVGedQRVSJOBtB5q8o94fiDvzwoXb1lllkdjogI9CaN
DPfrQ3e8PKuWr4njCR2yOp4I8q07ZQq8YAI/slceB9R5W4W4D9Laq5VHAw8yaC6S33yQh+o6QFxh
fWdq9qUnBtqjvCW5gzR6OdS1mWnUZIjlp6GVYBVIIyCh1mebS4qB3nVDJo4MKG/FN8YSIAJV4SPH
iVTYtziQvSTRajpk/hcBm95aPoyFvqBglzEcxNTjrVmreQuMLGdNwZ9PTKEyj1mmLHA3kGWRyAMT
ZY0XQHgRSTHaGfx27cJ14EsIxNvuOtxLeI9U6RJfjMiCJIHO8/Y6d7Gfvxcn0+zu0Pfc5kFUXMrQ
XB2sR4fFoSZNkCz5mXYWfDM7aZd6rW13SeBduc+qAOvVRjJRHIC3gZ94JT2fX4dXii+ja5HNEDPK
Ip29dRCbBLHdE98sPs0MZ4wB0LEZViAa9FG0OOSEzwTNFBO9kkq46dswBgOmhWckGPqWnx9VtjIK
JRipIwPcBsB5wF75H5Pp0o2nn241g3udZKjIIihHF7bGBORS2ZFQFswJDMzr/PTbjKgNn9aUXO3W
+u6EcECJ3gF5f3M9RZxRWuE8safRSnzyQbIxklAC1taljhB1IlhT+t1CuRNfDOtow2idDqDuAlNH
jcC+uP6ax0vc07FBCnAznm8ovyq1vTOVV70LMcJKEQv3eg4ZjnDxN4iDb9EDFq4OxSp19gigx0xw
+0SMiK1kKJSN7DSSCJFgcMZKN8OZmTX75+GqAKpVJfyHoCb7zqe1BbkBqzQL7BLfO39u274kvUTH
TrMfUiCP9ngVrTR8BSk3+9mP6QvTPrjIEaQDwoZNMfWPYn2mjomkdPl2W/gXprB4mnqSxWfQHLUS
YLPwqJufFewy7sigGecVyr6bEVZvkr39k7cbtxgM012JW+UxqQZ1QDk1RwQKfTk+GJ3pEukR4RLl
d7A5k6JnZ6qs+zwqpCquK2Wyzd8x/mWodztu4mwTxI7FuQvhqdI2mEAK+rixXRt3SjEBTyc5f5SP
E8Og7xemJNnsC2moN1kaD/favqF+BHyIiSy9sX2X2fb/FiTx9H0yS+GS7K7H6YFFXC4OJRsjXVfi
Ld7Gm6BW552vt/S47sOaiXmdv5TL65Xj2pjykdHc+ayGt+RAk3sQYGK4/GzAx+TYjEWBwd/B+glF
giad2aLqPzTHgVvKtH7AKgLLzRX+J4fgYV9eMDXxIJZZIM230clm1qxY4JOtHCkX8+KkcPYPAA1p
+s9OorWafmdFEBbDmnMYqVrJ4I6C54NvM1W5fSq3awjeAONscJMjXLyJOJobCYtWVlr+8fXH4rK8
91HoiSC/OcluWNjEfQlpX/QkjX1hjQyJDrQ9xijGkJ/VH6ltGFN+UuFEk3zZXdft4MwewGCmV67Y
SIgZ1+1+njuFxneZAVZ+i7pIR7tEcM2gRB3LYXVtRs8eFM4hstMm7TutKxq71PI/lyfqu9LAYNgW
9mSSYlU+x9NqpY8jlIHC87t8lSW+JjR/2DDx2Xf9XGESZoaV1XZmRdT3msKRl/phUJnBgrdfQdTJ
sn4p3ueBSATTAkwQZJX5SN9n/zM9ITLSKaYmisl+us5v4QvWUpkamiZZ4BjpVXDkesuged34gkTi
iinoX2CDQNa0q5YWsoKIuBt04RVocLyVavXS13g6TG4Xtj84dwSzZtMB8lAiKeH3xQXKKVgUqVJc
2GGJs2Q88NPiJS8XLs7VQal7v36Ex0L1lDcfSeuQHLRHlFl3Q7l4tiS3joiYzfyRPeM4AGPVWny2
ruPFJrdcUl7XN6pjoa2tu5X83szfiaUm9IVwH+5nuo4CtTlRKzjlug31Ng01HBg/RLG8rE4Gu8DL
hfL6P4vIvLS44/g83l9GmDMgSMhmO9t5xcOgWBIQT6FXDcGhuPjzI72hBUIKW45w9NrSHsN9D+95
e/D85tIC3yeXWTSfWKJKVwn14wVKWvI7NbfAgGZke1xmITy1EWym3fyafwvvxSvimi64khMytOu5
B4JYe0Y6ZwB9fm5PKvGE6M7SB6YgsQDGhwO+ZQNr7TP1pRn+hyJYBGe3PV/UPz76kGuL5AwlgzUa
25xV8sT4/dZHjd/QNhyUEQydb0UbHc6WXK65Cbk4bv50VCp2UiW5+Ko7WmxqIi01dLxJh9JncNXh
GL6egVZkc2kvSNT5qOFKP0dtHYn4ecQ6y44JWT1bIyUFw6Vu0nCShAeLdT/WSzaMl5sYu+SUbfHv
J1D88w/kD+6IDpU0/oDOwzTUQpdxTzZvIvpop3BlO8osP90XpcLEjqXiU/IOEbyWlQEuZ/HQ6KFF
5JohSJDWKO8uES7eiF3Gh9hEeZ1Vk+HpfquNxZ4C2NXGYd6SfL0EBDRch2MoVk+N2+Jp7lph7ym1
tC6Lfa4Nf4i8dQNK8gdhagVVTBAHI2uhTNSgBz9sPgCum0Q9xUSMrGDiiExbo4VA4HfeXjADYRMN
XmtiYKj8BUKhS+54++18ipp/46ntN8BnFnj5KPEVswlf67szYAGHXcBnImQKegD54w5eohv75xug
2A5lLSFs9RAkcfFrgIs1HFzHp00ywcN1iQr+6SsAjCxkmV02L/mPflotaBothMt4HKyfnq2O1nTI
iZ5gddxYByxQn8vIDKnv0O/UgrMkhhpScgQmaOQMrs3m0HwAE4lppGzMTT2xeDQfVwTmYLOMjoX1
xArX6KmA38Ap/+3gb0PPYpNSKMYQXD+ZykFQr5tK/4OfNWTMQo3e+B8LafFCg1eAKie07nrF+MJL
riMlWPCP8EOfpZRiuUISK/Z9EJww3BcR6cu14vLRdiq5zX405eN5ayhZzK4A9g03FJvK/2ARzxyi
91ca9S+NfTPERzz2wor787f4Bcn6ZttPQm4T3qwE1C+g5QQxlPInm7U4TDN8v79GX9i5ZhPX3lsc
vwJJ8BxhQXaXDeSLhoVy7qoCobJKXsWjhwPL/vH5JBzsUaOs5Aaqz/bIy75lN0GJGenwmXgH5pH1
9bRiifkSPPDRe1B6R8mzpHs8EXZYX5I6qWmNOdjxOjl9nOg7AIUMBRwgtlX0DVribUMF0dyu5HWa
POSYxw5/3y8vcYjOxZ5oBEVg/yd0OUtotL9O+eNIZNYXcs3UQ9QJ05/bYyXInc6dANmcawNfzdpF
PiN/6xURmMXOmUen1aZV6FEfCXpOZhyrsjCKYNaR2E/2whMfLkV06NlXSH026N4xumHpIJVfIr1B
6achuR2qj6E22rjbxb1dhVLW1m3dqnhUp5crBkicIjUblyr3snNvgLJ7tcQybiMkEXh7BaUMo+kQ
SnYq0zmzUfGYiynCOD175c8fLWSlNG3DsTYzeJ4xS2uC2VY0EOlnABxC1jMxRuveuQxO6s13ySIn
jUbiA+SEfbOB3AIS0/UxcGQDFwYyghB8hGhkZv/tv8sNqLWzjLIeV29GtgD/tMrUAFj5ZLj73U9a
MVKgnXMmrLfDYD8U5y5uVFzIKrpoe7Pi1bLDDf3HoBSjNCFXoC6M3I9BThsPOSYLXxXSjqmWNLC+
+Y1SMytpNdD8ET1fUgePwqzgD/yyY380CNB5IblZWckZPPXJMEuYaA/ge88EUo5K+bSd5AwKJLZP
AuQJDfIFIxBYnLPt/2rwb0Ui8V1Ibp+pIWPt3VOchXKnAGis67Zlwn8n63tiSumvCg8QBG4uE2d9
GAWUfqtds9RFdTzAQw277EkAZespv4UQRseyeYPJlx5UPbqDPMpDh5GC8LSuuBUKpKR6L38p5tNv
9c18BUG8zXprcFtT93vJ4O14Kfhytb/8+bsep9K+xo5qDU7TKTX1GLL2jcuwCoTKbSlf59+Bm7r0
I6cnS2vPxeramc52wvG6VUurjTvCqiX+er4QJWUAcR5291fQqqSEmBiRrPpnQVzoOq7FhzQaDcBt
//FDPmdhFqpbulu/hy+aK20BQ3yZVE92qC57CCAPGENN/v8rda3Sn9I8MTTerPXqlnPKpoKeKxzU
poVNUzyBnQzhSYm5fLgevY6WrRWDqJUBmYN08DewL9xGx27WylMGuPJe4YVs3d+PetfjpXLnayXX
pANdH+j0ehLYzdjcDJw3SKl8LWWVHwPmPkMVPmX2IG7ZFN933fUaSjYmieQrvRUqLXCBzJRrFhyi
DfjNU4Z4LhQcDvo6Z8TQ9LaMhlW1XIRlJmJjET7eId+fFHJ/xmaibSqSvDLnw/JKkt8+1wTaBewe
wH0q5h3YvdT00UMrAviQ2JFs1gCNyewKJCN0YpFwjPfSFa4+JS9yIPSYueQUkoyscE6hPRoudBR1
tlWo4CyWrCi+Grxkkhhnfx52hrqtrMAOrVrbUFRvyflQTOe3b7rD38mbTgOlYt2mrN1gKVWeeVZ+
m/kKHVi9q2dDjKBqhEM5YsDmHWEfklRcIx2Bopptz1ILZeoAHnl0Ev4UDAaMGHJIHrh+W+4OdaEG
w1jhiroHBdGQBW96/CKOtfRW0XAUbei3QwlUnw3/uq5XgHh1s81DtNFIwzz0tny/x3A22jkFocKg
wRGgw1xwhkt80j18Dc2a7EOpVDy3fvhl9L1Utv5n+PGy5ZtdPGauW1lxy11vgMHBHIvnS9qnljMe
NTwIHRD8A/mTSKa/Vw0Ib7ku4l3w5K6Cl5Lu1qqOhBJaGJvQRV0bvx+weCYDW+W8SIDyKXIDH36B
06arcZSljtiJAC+gnzFJSj9uxiy/TVWW4rD64INqp4BSfnG1b6i3xNbKoDkbVgz2SIHRKWZvt0vY
qsKxj5CekehL6UJbMPS0oiaMcOTBaL4IRxZJzIBwnQm8mwe1yTnyr/a+Jao5pTwN5qwNqelQKd+6
qR11jf5lGH9Cc9Eu8ObSgJONHrIA70blQWJqWtHTdP9bfI6lG53lupQBwZByjnI0WaDPbFDxYYIc
td/MbwoN2AtRlO6s3pK4yeR5dF63L8hPayOx3T8xZFAoiShrCwOFjcH4WhqESPOoUdXwV4WE3EeY
oIE8ji9cZ/BepGrDUOIu0MWS9dZ/TjznzsKNAU7ACWMShiM6xtNDTzSOnnqpA726ofaVN/CZmOJI
hibA8nqADM41mn7Q1LvCn2ulx/nvkX6LHo+QSjHLyxyqvSkWie+YDtIv3sn7dai5L3kFwy5Ez87v
PlhvF3pAIan1MCBq+Beh3QJ4rKPfrMDvxSWRFmr7KFgk/X4d8aD+yb8GRtx0ugl5DQr2BfHxkwyh
WUT8Clqw45aUA0pkB9n5fZtXLpZ0qKzQNphRz+bM2fC/RMn3R1acwgn2UL5Qhms0bTmO4NfH6i/W
g/OPWUoucWx41gm1O/6CfxntaghNc+BM9YNQhitLt3rGsIhaFjnExO+k0bJIDnN3GExb10GVNH+F
UiS87/VTO4GH87q6dUeYDRIFDNlsBteuT48RWwEiZyMBKfOvsh9PUarMZ2S4ax5+0hfEZ0u2InO5
wTC+wwQgyT63OyNORebrsXkeVCH2Uc39deYRL7RSREk6Q3ASfd4aA//t9x3MJ7THe6MySDhPK/LF
9iYIdPB536yPbHqHI1bcX0H/ZxHu3QcVXKv2sMeXyK8mPj4kZAomUQF2Q0WPbwudcgrcaYi491t1
hahLZ0Wfm98jgliDljDqA0etOMl13I2f/8JX9RBQgvRO1vxBD4zGNBIpFbiCHbQmq35t7br7t5PA
eHzqulp0NP3egnRHl+PcyLLrG+mHi+Ms6LvjxOL5Ld1gOW8JthjDOqR+bvff/w8XFeA8fZX2s4mb
o8ZQL9AfH0P50pQA69k+bn0QElOhZmjWREF78Xc3Y0v07xSj/8ppcOyfQlpXcfFJhxhNbWx4T/gz
aKVEfpliwaV9ip4qk0N39d1cumTYYsBq4SioG3x3q6W0n2wj690Jy8aC6frQL84q4BDluRRtZm5D
j6oo16VyK53VCicV950MYbiT4jbwxLLFo+oD1Gd6vV+jraBjd6jaQDbo2aKvO20tmgths19VbCgg
kdGiphz+RC8VNJ2lxn5FMJC2NLsjOWERP/sxn9A5SZ4Xw9TMfJSXQWbt8QBRl1tiPu3yVE+w0gk4
eYCpxarw3YL3zGcKKXLw3qU14a0mGJjiEsIDBu76C86a4UtZlOylgZDHyZ7ehqEnbpDaQhhVOllZ
PZUi2hVbClWtvxx5tSjVbhKs15mLynVxc8o1MeO1FkmQUuyNzv6kvnEcT6sVIElkFBzeY4XLxQZm
2eMGNIiAVLTseVXJWfMh3xAk0Baz8GQ1mV4LQpsWW5BLs68GO5r5N1mxUhZZwuSqRiVbgntGed1p
kjCRU4SsJT0nXOcBUt5LmCWkvaD1/rl4sVrmZxs6b15u61neojlPg48/4wR5/SmrSIs7BeHuGbz1
/2j15VeR+olyoVL7rWgnsVf/So5lcQXn8vfPY3SyNi9M/UciENRq+EFsHLypqfk16pfSIJBW+XB6
cVGQZKUZG7cshhuO3IXMkaunvpNkMePVijcFcvT7e+EU7Mw1kFlnJQZyR1v9LC9VHJqlVWpG8aKy
DqW8dJUVQ4LODB6TJy+HUim+nM8fXZ+pqVjwkhgLGcpGHgeDecl3nKX7XChh9dgICrSYZrRLtBuc
eqN2XQFw5KE0h4UonOT4PfofBjBX35sGAmS04G3T4ORh5U8dzEHdtLtQfHoJGe74dGIRalYuKC2a
UbH+ZmhTlTC3nIJOzyaUwvWfmUtMJ5m7Wliksg4/vI7zUfEbV0CTgluv1xbKSd7OtGBFm3lCNoOR
k5eu9ox56HpO3EFUoHLaUqqEPc7RqD/Al017oHabY28g0TUbX4E26ii8Dkr3h6fefX8GS07QICWQ
esNmnmy/A8z3kGUeicunVY9Wy4BN5e63plfWOtst1XQAwgHoyz1wfuatujNNSVgdiKpJ+c44StFM
acLK2n59uMSOO0WFrNDoU4XtynLxWqYOVKwnmAQypx4gwATSj2g0oiE6l7OD6Fr4nchxODjrr3V9
6kyxhyGQwZz/TzG0x4MoKVjbYqUcsyqecKN4gWUr4nMAOxTf11QKlpOpYtqfu56HpWXH72t2Ck+r
qUjqm6sUgushjE7ICi8MFKq5yc9JKE5EQKDFPSZ3iAsLzGJuqH9S8Eh9B1PiK2iicx8TNJQTFlxt
VBjmtpB3JeraEa0PB7bDuEx1we5lJy+Oz9vMGeaeszlvzyiOkIfE1/ofB66nWxABwuwW0Yzunc2u
DNXWu7wzyAERq3YAF6J7Ipz/7mFz2a45Fv3erzSAfFkx9r+QW+dq3TtgSaDXXPC1CftSDdzhSCfx
jHDf9YMUQJqleqJ+i/X0aR3ICMtlZsd55+AnJPZ+XhlNHC3+Fpx1ZUx+Ay3vJbY2wpnkWtXZftQ4
cyjXHKieL9W1mYsfgHTxA9vuP8pf4QtBkICZ+lpNRRV1q2yLrcpxf6Sm3NJI3ffFEi9kFSV5D4ut
S5lTUfskmmfnO65uGzCoaw2NeUkptxcvDFvDdNcIvjfHN97NhaVuGSv9adwfG7bpinqBEjXgfKBi
LDaZDCaFF0Jbc3A0hwKiM+lTh8UDKAsXpUS1UIWprgfeBCtM7OhIzMQc9mPqsx/e6Lqx5qadC5B4
GP/5/AaAuNZJ8VGzRyWwJussKdAojas/eEWGOu3YJDnjpMi8Z7f3l1xywli8yfgy5gfvNnA8fAK4
D84ZXPAqHQ41cTxO8AMPXt3pl2R1GIsFN0vNj8KIQ1rLYyB3qpRvAMSU6xtUdbqgSBD9cNYaeVH5
dnrcZVILsd2q92QGfzElNExsMTSwQKSBenp8pcNCRA3FOHoh8EfO3EIBDXC63UvYoMJB0vefHGYe
v5O0FBe26qXo/7HUjZ1dLnQrEzbUvDtLTCSggW/bcbqs2ajFf2x2t5R3RLbTMr2DcBmPiCkKw3j2
r+F2jhFssnbgmJuG8rS9h+BYV+n4TwYJpbxeK5/4C4BfANPb/97+O7BIzmj2SR8xJbGfu8xajfJM
lE2mF4PXTu4DHp9fcEz01uiBwX5bIApGSuHYNzj5WNU/JuWNlWq3pGx9Gy9HIPCrm2DrUsmnKQ/3
kQeoSNbJorZAOuZqWyBpuD7LUYM6wM7TTZj2sDwahB9pZNjQB35JBNp687HmnYO5p4P/CAcIAFTR
P/MDZBHpNhffHSGwtn0aZhFfKqmH1W6KvhK3whsdlDibJohzS62BiCv5llmRTb+cMA9ZV3y4T9s1
6IFGzA2Oiz9wLw1cCJ8uusvQCj8eVyFs9l+R4Wki2etP2KFEypUg7+kKzno9jjf4WQe1PMQWtJmP
+Jro/LqihCq2RMm/FrnotOJB/s+7q8EY6MAGR5Dq7Ec4l/+q/iEr03lHBAOgnHqtLdNeFl4C3R8o
x1aygt1kIqJNJ2E9orpWHtvfQ43fi/2gjl7iLBdENWeNmn1RelU2R/1TOCNwS/NV0JWXgtL1ajIK
wnCPicos/AjLcLbrFmhqdxUToLCTZBG4VPqMlSrYtHvgGm1B3T2SBVgfggByLZHzavbaaeb8PY5H
RLo1O/aSklK4T8JmAgri6eF5Cph0C/uRyMmxxAlkg3rWb+s3FLfNbXb4BIFzaXt9DOFoYqZ4JJtW
tGVHBYr3MtszVHJ8zD36D6k1qPQIF3DPGEvvw3pjk+ziHwGCfzXsGiHX5brPJxPF2OYH+0wUqXzp
AfTHbkPW9AT5hSq6SWgTH2q3iTiR0BthrOUUJ69n/KNhUtxhV/GnI4FEdkUXGBMZ3qjb7T9fgeVg
j4l0qT0LXInG9+UrJ3X0up8BDQDuR1y9wOVpqWOAXlRdPHZgL11/bI4pWbkhmgyeHR2q8JJnshUx
wJbWlgto4cYRY3sKDhbrKe+xGr3GJiGnPlicSUcoYQyRtmgkKfTPna6jucjfroHpQ2CQxNqpN79V
cOjs6GRnyP/C5yK/z+fFmN2q/3l1dOYU1SRV//MLPoWRcTY6/s+LN6xKGtG+kbv3FHsLUzlHvNTR
xbk+bJEWLPZ4wQUewow/x4vMP8/gWfJ7ow3Ciula4sJuBrKEaL6FvjexscZgTsStPuU/PGsTvAir
qhGoIhPyG2UXKE62nw1MySDTS8eXTd+8ceuo+aa0WtWu40upr0Drk9MSdJXfcEynqS+7fD+Gtze3
ZNj2eysp1INkUsMmdcnCOHBbhmsZlXd7HVnmX+bcHzlL0sRtZLc6bXAqiJmR3LOaSEQ7fpHsftFp
7W81bNHr3scTdE+QTgwADmHWQjTuOJkimiUu9Sxp0VnvH6rnZF1raB2sMQS85qZzU91u+XQxv5ZX
mDNGGLrEFykprzwKDCI71dE3Xz/S8gmxwOPLb+M1je8JAg/zmGJ7f0SK0EHv2smnAoNucOSRBJNY
O4KD2WKqnA7zTiPwl9c/iAdGMAIXBZDQx/w30wh2eZ/szgoINq+XE/cKnY8noPjxawojK8WCEpD2
ddoshxzH7Xs/cUXxPHN+i+7xQicZAsiD0AceW4a94jRWOyc9lecsnaAitix8HqZJtSbcBuWsU59P
YdYQ8MMbCCzxhFRVLVvM80EvIdTUDaYlwEx5HOUuG701i8TvJlxZaF4zcAn0Zg96683iqF0w0aee
wFzJnGR2JLT0YUwzo85xuCpcNY+AoZuBI8fu66GRrfQ+7f1pfEJClALvPhY/xbdBFhwd9oBos5E9
sG9L56RnP18NqNiDyUU9agcS1QQOdHZNt6nszl3ijiyd7c9jB1HqiWQS3DgMOK9vcoKUjXk387lO
IRLZoa+25DiEVaI5e4k6Qn2syZboRZYTuvrVMbUOAf/yO9++lk2UXIz5PHvNkDXnk8yr3jeCUeEt
zFgJFC7uPqQfIX0QxM+SpxDFOeb52Opr62pgMQg+qKvc2jn3C2CPLT9mX2wseon7byrXNYBxdsHK
dwCqINd4rT0+uhg73cTKQTsfBN/88NCkeLCWrUrbQ9Pw8CftzjJAv14PvP8Q28Z3RHemRjXDYsrW
dQyDIqJRJoKS9gRV7V8Q9ZF0uFo7L6BOtBl5z5ZtTo/WV2snwUAZ720fJVLZ5YPcxoUbsEzIs2S5
ltG75iyTvPUq2FKyjF8Zyi5J33LYJE81YpTe+LTd8ovva3XAfSPbpE5+ia1ice3rfH5dxXvklDZs
N6PDtS6fzu6X6fDbsRD2kuNnGPf6hX5JckkwA5MKL9q4bFsRe/iM0xZ0P6yOUjvxUl29K+jc22JU
JHnsvChLUypxClrQnkMcawm67eP/kmsi2cDRjHirwMAsaqDw0F78TQJk0R6cj11GbIrs7Xth3K9B
Gtxzj5cxMf4Rme1/MvOY+rwPay3A/DlnM5nhs2+8m3vqv3v8qnZYfSpCY4MRAepjG7tS16feDBjK
mt69mmBpowQvIrVerPJQh7b8Z2haGrO7F5hq2lWi0yyCPN4jQ47fCmTUTe99ODC02SxdP8XOH4GS
LfHfBqy1aEPQPr5TeHgM1RMbYNqtsIXbaRo9P2bdWq1E6NYguB5Y3JJ9v3g3vJGmVwRu+oVZsndy
ArpaNtUgsJ7l5xbdS8oWZOzgY+WwTtVhd7mQirfVKK6I9ZXBL7G9/6uVfUmHvdChJg9doFbzU2tg
sfg3o/0tqJwhZ17rYLImY1ANPtdut5LhaThEiMjqa7NNGB8nZhHQrocqdhqbXkCyDgDsPrZcQK2M
Fc8pduCX3MOD613+ZjaN/e8CFQVj5pVL6EaALS6S50jezbSfXVSaRT5N+ZMm2Hvimi51EGx3WmgC
BGkJON4lU9B0iGHRTJKpeFR+4u3wL5cH6gN/82bpgMk67csoyDnW3Ro2VPhWrTt9RA5783W92HrO
s5kBj7rLFSj9qBNzGb+kMPGOP2dAwrF195AHFM+xvuVwcsf2m0Kp4+5x8Hb5exV9B14rzLpDmBLK
DbzmIwNRju82s+aBGm6rizpt3EpIAC5a3GzOVEffEJTFk1ZWv0BhASi8gKqGTdoucVD/QIAOITKP
PFFBKd+Ya81jDBYTyJ7tNZZP4YQHb8vXg9uj9Hd64NN57eYw5wv81YjcKH9W2sAJyrZaoM1v/hq0
IqXxNaVIYGoJqv6CdY+zbbZRnsiah9Q9Mc2eRRyYu8Q3M2pMkjrIMT1tSylWCUiqWQQyg4N25eab
gpoDAq4Iwv3/wFADVH8pDxE2x8hTLzvsc3J5InYlL0JxJTLgVmdB58NqhbVjCa3u36ikm+LEBR6L
2Yciwby4Ty3RlQ4AC+WK0gzm4xjc6Klc7QHaSe//qTTb6xlCvk5GWZCoqhOBVLhWcbl8cdY3gHhj
mu7Lx965W7bhOcTGjxWc+TikJ4uEfqiezyBdu5WTVT9NtcbongiVKto0snWm+ivjXxbD++1i+fzK
aA/Wb3s/XRfOZ9CBbRkVBKRqUQVcrL77G2col/KjQqFgBHBY2qqbzPJQPXoxL0Ie1pLMTYlsIj95
XI+XCaHgf29NKj4WbxjkvtRaTiiapHsZMxF7mcrOGg30yJ3B7n4tuL3TW56I+/MMRDBLAogOAs98
wGUmZrH0S2K42qF8B1SJLvGQGV9we8wwUvoUkC8SX3H/IjukWkYm+/tC1CL8x1xBx9d/vcFmROQO
5JJGTev1RooRErrdjMThENnthXcFzYUcIFDZ2p4UeXmL7bPo2D8iWAd9e7v1y6Z+6MPakGZ+HeY1
cvrfLdqGAgyoDqxUf3WgS+5kPbrA8spwyU90NOzlOHkcbCE0pXF13iEXy5F72MH31ksBB9w94XpV
B1lxPHHxSFtpkREiIYv5gY64ywLxLKWmOZG0PIO7h/gbFCeYaa5wVGCITLIn8TMLaRT6Kb+VRBgA
7guexhc1cgRTi6Jk18M8C2InZtrMzxTVMx50QnDOmL5vPa5xbE1fqrpyhBQdL+hCr00msJUvLEGO
NfP/TU4Zh2E8gCuGYSb4yFs7rv4mJTe/uTtOYkLVYxnzwESM9O5n4EztiIyoRbdeiC9ad3RVZo5z
OW9F0zeFs424qNkOW9Vvz4tP/NVbrKmsYolcZlJF1Pk9+Ptk91pbBKd4pDixvgMateQPZUdJNsmg
116U8nc/cnFK7ofMvKWYa+ISJOsOgzuv9J7yeNWPNNucdrP4HhIbTxtyWI4PO9+AHjUU7UQ3RQQn
ZyS1AKrrQRRJndzlATR/md6huJtL2BqDjAx733kBPogzhIV4uFELb96l9I9s9IKbMpxIyM+VkgxC
JWsL5eGQiP13/TWv2cHqJPzsKXSyklZlCqXeuE8LVTMfw5Y80MM+W6KNlevpryf8RX0LA1GGgHEr
yiC9p9V3XEnACGFzxJojIY80k3a4tiYPIvzg7HJETdGtGNVbgidZS56AIx9etABWFSeN2vEebrLe
EqNZlQFstf54IrwkKx9ldYGr0+CLekZL+9rYhcUnXMBsuR3V4Ip08wH+USkG65nsY/8zWhobq4YG
BT09hzjU70u+Tq+mVqPSJDhPoxDdnxnTxZWRB6TmYAqXPPVctuSEWVUcgRjouR2Z3aP3iEhVhXFu
05xWPBoSQLMmqUTpqE6fYnG3Sww9azrVr+ik+Cu5OLRbDXsL5nkwFqs1dcf/eTFS4fnkdtKCb/Ip
78igipBjVIAprd/Wtz5vLQkMuw1I4IZXXKNKnNskaibn80iaO0QbBoq3r8HoOYmXmG1X88HWzjyL
cWXqpQqR3I2BfF3DSyBhZ0+Jl0V5fX3vET+eczJd15AWrehZnZXtAVQ2P1M6vNJqpTHC8v7tmQYu
Fn+vCkyk+yPGM+2C2htwlw5Rd79L2hjalL3b4LT+RYc8PuN2FOGQt62AyBnENuG/LZ+XONpvWt1k
pSsYffMbZt9hq39s+2h4RVoNJg+Nb/OXgilj4VHnuskEYvbe2a9OgvhoyGp2HvLw4o1PxuuPjclg
MHEumgGv6E7LDajj/iWSpBxaUdG5/zSeuoBxFy9iBTDnNfZF3Lwd/3jU6mStReZDTLS/uD7wZlru
INqr0zm3nWpUWJTl54aXuEzYMXcFY8HoiZwIFHgww+T5DWBUySRLGvrdLkbZPCxUCJogKGTQ6AVY
pSel6xmtZbIePklxcNxrUCcZR4MnYdqUhE6E4KAKu843WKrYvzunHIYwybaZ6qPzb7KT3jGe8lzl
b76IAxrEhNVXbJf3Ftl6lKxXKXnja83hEYvNj5U92/7xAYKXPvTcqEoATHmJGPuBxoCn0KBlRNPO
Lqu8NNhEZFxfxcVGsnt/+aZzqvXlVFGePr3uePhRCJAVsKTHkhwKYmL5Yx/sGoh80r6yOuCG4J1R
Y2Kr7RLiKrwTduvneA+GLRP8HHAkDJnhDpxLSqkEh5PQp9RK6eQDv0Q1wi/jJNx3B60VOg2iZAlR
d60bF2BE/wBuGaUSgWi76xQRgsQSS3JdvqLkfV6OUHFkJtBODHMbPmL/Walw88OXGztIXbRUG86J
3aur4QdEjv/gt5dyuisEFtl1oZLnunO71hiq2idjcm0sywfjjKQ01qcH9EbudZ09dazEm7Lucg8A
dAj22hbwj2WQg+SwSlcfrVP6j5Ix7Ly13vBeeUuail+Yunog4i2eplcKRW8rW/Xu9U7W/xc/wGFZ
sFisxYjp+VFxTFdj2EDK/W9wIoZeOT8/VAoYLuKRqZ5F9V1vCxYRwO9xAMgA9Nt9kEVimJGe2j+V
oyn7h4kYUa0cIIyQJwZfcX57ITs3oxs57TV7C0D3rmOr7HingG4ftB3rGOD3xqjPN3vxtEU+90Z5
zQwMlQ8lcqZVdRvyJ0/30bbxQPzpEw21J1WQlIQibU6CuzC4ifIb6yjGXhlzw/c4PUMkzWM+fbBZ
5EDomRn278N8KEvt7+wCMKQ1HF3bWTQ2C3mK4bGX2uGeqd4yQ3u41b8pQ3qwFdyA5ry/R/qOuzvD
j9/V/P00lMMZsfiadz+Gq7r+5h1hfAPUgHFN36icmRs5Q2SZN9MDej4mfL01UNr6/BAxXEbhseKL
a9DRTSTr5VB3LC2ZQ43mX2UTYuVk2wRo0T+dVAZvzC088L2WT3vlFp0C19OP83FfAvWu/xsyXDSY
4uJfRoPC8DqG0HEygPQMIQeFfGXr9DV2GJsazrIyEjuQnP1w6I0k8YGqxXLz/VazFT88G83jMLq5
6SioCCyKlW9/yq/K/CqdVsE71uMvaUHA+waVh72xYEJhIYABuuIZWR+PImWBuRH9x+tIRcB8UfOz
Ne9gp/XEkz/rwsmKGYT0OV/DRatg36sLiPYQ0cVTDmHEMPc1KXW60zkohI/dcjlBAhMuv/73BTa/
rCOnry9qVQ3UL5raFaE5RTn8wdGGbGoPbLsrQPkG+gi65y82RMn5vH16Yf/1DpELLqbnZABbTKRm
6IgexGZLxS77cA9l2z36yeZWMBosYEe4fFmrlFPwUSo3z3GC8B5zEuSuNhm1gqeloMTh4t7eetAW
lm+9a5Qq/wnYsnLlJffY8Lca7iLFG8MKF2TKzUW4k+o/z3tvBZQ6SFoG8T+8gX89vWUTzB7uV9vg
EwW/VWKbLBDfhqZwp9qI9j2nBHHrcxIGcaCG0w4hsxuaAbKLCaPMADVqFhRH9HkR+FBDpTVhHXYi
niEc3mJ0C93rwR7idOo5lLEdeJJmXqnlZ/15hRtgnxU0N+t1e/qCOWzkUmlS9j8Yj3wHrwX7+yaQ
uFicU9hZVF4FE/A4Bgruvx4aUcjNRa+LhdZhHcYxeYjE2NDW7Xs9/J87yCxRVTvEuGjug+28AYaP
oGA4bsM8Z0F47zR/bobzvIx4Iu9spp5rTNRx16rD0uV+wI7xQgwBfTOkybX7YpaaO1kHSEzegU37
9Z1429qRaAh28MxjgBGESOOTPAv/bnCKRAq1HcVbwFrlVVAmjdiimmLBsGIAf742Zp5/tzOCaxv8
aQcZm5s3Bkeo8b8qb/dhxveGto4UFLZZdt60hu+4NYpjtqwk7ckVXDRlKIkZIMP1yhyGfbcu/BPB
fyVXn3AHYY3W0JpVV0SRzysvPclBEqyxMP9e8OxcTBoEiCALc6bSyElSJx7kBV8I2eqviLQJmArP
8rKUhWkhAMfJNDRGjmNHlgoyaGd0ZbNsaB04WInjwC9D81TbS6sQAl1lSaEeqUFJv43751PwTnPj
dlKCK1sPaOOCBoDQEWBOXIDXov44Z6ZbEOB9FhS6kv8PFc/FLQPO5pgV//040bI346wXJWUJ/qmp
aOUGPB4CEZjWRGWENsXxuqvn9h3Z5W4flzCo9piRl3lADjYwdeY4iKu9ou396/QKu0ZLbevS841H
Vn1tOBWsjfRWxKzpKqf2egdMEdJtfdJ35Nt5gxvBHP7TP81wqaowlYvmGi+pjY0XDD92bjR7KpFS
qSbbbI2KJR1U28ioNcOG1EyAT0BAtvzRcNLpG0wtRUog/4Lkwx2Ta24VWNe9L0u8d9aM9k5khdTN
wbzlXGRLwMxmMuLrTFpN1nhxxBpk5YxRGvgZlk8XsclvGMCDxf/dW1zQxyyJLPKzonl/+bHOOPnP
uAwBuAEDNDK/AnX6+yfzM/ekbQSI4naF81zH3mka75e6cOfGWd4LVeL7+wZOatZd+DF8nJYEfLYO
cRLfyM0pHe4Bke5QeATYYf3B2rkUGXdvwNPN/NTV/SxyfS9TvrcrLlrKp1gwERKDKEcCV4smRe85
CYb2OYyOtaMc65Hu9pB081AOCAkm1R2m+WKyjkocvQmxEtZWepEHeLCaz9BBV2pHt58ThzBH94zz
k4i3i/U1PZRWGfnyvyrQs47kBNYfBj9gy9SDHP35Jcv17qIpT0zYUEvLs/goNyWpzfkGMJpNFMAJ
qHJv4QoIleSqDYXxJv1EpY/edPsCqZjbbu3GKZUdg7ZIGLAFgZ5zwjgD6Gmukoynx8aa60VDaaTm
hrDSYXppxITlHXEAAcPMxvPq6H42gSuoDF8hDbKiXqjVx63v9ydtAZ/x+nJtIYeS1OnpZugU1NNu
gaZ2T6cRVhRXN6gTV/Iyhu4TY75fHnl5sfz64VoUQ8fr0dLLPyb9ebdWNUgwuEYNxTpZz3noLWkm
/9opsNPVGK/mQ0oyaig8+aSkDA0kpqZDn2xIdWBxYwHGd9wOO3U5vLeZJAJXunX0weGwG7/UQ2OI
FDQHxJljTYGdkqYL2+hgD5K2aclt8GfeHLl3ItoOz9foZTiF9HY2mU43cYeMA92aFJttFtCpCgXr
gfV45ut5uUhR/urDWzDXgndURQwkoQciz4vnEuqdXjfL4CqLmz2sEUCtPN3zdF6EmrG6gtFi0L7z
7LuB3hmFrlYK5An15DTkrXWEDCyLHYUCVGf1bw3zSx3tePMnty8dPYyy7J8qmFk1MmQhOetXoizt
7wmHw+oOuxyd6yVPAqoTL137F1p/d6vnf+hU/kJndXE+oWRAUccda2Hl9aQS7wvISVMaU3RcgPv+
oAzwhUAbNpNGdGNTg2CPjiWbxb6l+C7hOb64o8MthOEGDB904tETb+Q02r0A1e83wuFXCTQEvSiq
extEo/YiRkZKwtJvsSM105c9wBmCO7jtKF3rN1SqCmzue05Pj0Dmyhc3KT/9aRSh6lpJE9bPb+C6
YvYW0iEUid/ZZJEakhJpt82hwNGxmVIGtY+JXtvXcRttH/GiWVVDceNjRt2yJ5tLX0x8uLZvJGoh
DI7aES3UZ8yfQCf4LUuSTrDoeMQu2nhQ07NTJf3f3fIr/FuAkAAJp6U3Zp48UZ2H5yMIPZFqalcF
+stMWIyPWlzW8DYJnYxJvg78uAjuOyGSezGslF6qK+08gmZzEsdOalKxhZRlkm6wI4jY2tP1Z88t
cmC/z3FU268BES1TjQ16vImn1447DRpJATdRIvq/f616u7qezLd8KHn4CUYpinb1QxkdmBsT4Ezk
UhSitw/tedjopQ1LIsYJO/mF3zPQcZ4QLobtXWBi3clMOz3R33jQxCvldma4LaeDRYzEsXW99gw5
718R5VIpsdqUrmeoHdkS11uHIRB53pLjSVr/pn2epLV+bYgrq0sfMudyFSr5isH4NmlojBCF7xnU
aaQAWyehKBHuR5rNyZFyCIgGDlmAYwpA+Kvb5Nw6268dLnqtjn9wdqA5A16vJ25Pbvnui1UEbmNr
7SDXXcXGHCSR+BfkMDcuRxilvYtcJUCtX7sY5atE4W3y5JaZe20LsAqRrBDTHrM/gVSjl7ksdMyB
O6KT/R8argCcbTsRBGw+oitiyauziHNFDwCBJE0ilja1YtU4x02c6movEFrf3FXdjGBQ1rV2rxnc
AKn3XRsGE15h3COi7h1ttKbfjpkM0kpwlt75KC2lmzHbrTz0Ja3JuegRcMgjBAUpzCJ82XqKyHij
F+b6VV1dKPkg5e2OOhAN1kDkp37KI8FOzokXjgu0+vaKeRT+AKqt37IiEOss98AgXQR6AWac2oxY
LRcWCM4Sn1BEp260SlJD6bAj44utfsI42lGSYHcVMQ5dpW4dvKboFUa6xSOzxxKqSUHELAL6OAUS
t2YtbdxCuvFqFa6D+SPiA9nn6zG+lYxpp14x9+gQ+oB8cZ9O+ByCxGaWhSxSTrbRjBHHLVrf8c0b
27l6tErPo3jvk2DZawiMC4IFYWvXQVxKPR5+hOEXGF4QahxWAVYCIeusJoZjZKZG+Y/Ep56J9niL
m/SK/Bp3h/EnvTO67KyzS+QuPMd8npqBuW88KAIddYv97PXzwlZ9WlhuQMrbdG5BvoidVNw7wjM/
Rjh+36NgtPlibCmjG/msKHxa99OBja4Eftc08D3IeLN2nBQ02mekyQkxOtlJuFUm6eVWXLgTLSrK
O2/UluqXkGD/6ynmG6za9i1Yj0CRmDuURxSAzgfhTIouqgsgXM3tZG+xl764tWO6ptqprBe9dTAq
rhwhxLKzcvOQRNHRKgaCSh2pwy+TF6/V3dNSOQvJTB6UxwV7RXXt6C0eFD7LDriJogsq5L0HQZvf
SD/b/k7y4Mi7F9P3cuvG0tOtel1e0tEo1PQTPuLj6HzJZyL7/Mxksp8PO9RyqUFHbUWy/P7NFnpr
KMFahxj1pQA03HB2o+T7Cg6OD9TBUc38eTYjPQ5P5nmz19pUg+MM3HD4aQR3D012cHGM4zeNADHt
AXM4huyjYdg9T/pkgFkKJhPbD8bwDO1Ywhr9+TiEHUrcaZP3e1MAXFGJMdKiaJDaTgtXthtY43qb
cZifr4g/eNa2oUTHmJp37y19IqML+3UobzLuzEDIP1uT24KvXAZ+rmLwPewEolP1pHmIN0Mw26F1
Ex49OqFvOo4Haf9Ck9Ij22Ljk9uBnVTCPALiFInBIEXzyRMOhO2C/QSzRmR1SaK4dIynPMsd0Ll0
xUUOe8uD/QaBPlvSc8w13gLiLFND5PFWqvXhQqBfGn3htYoR3MrEtsM1muFxpnGwGS35P7muKFaz
9lL2qHT2RHgxWRs4j+a/PBtm9Ut1P7ajeUv6qlRPlBgvH43JqenSF8DPauRnO4yMEzdeoaOFfsAq
hDq/hL0Sy0sIrxoZ/ABtS+vywcf61OaL8X771aSQUs7/kF3mLqB+h20H4JgYE6xJaXcDLUeanDUH
mAdIei5X1lIBqpp4oVl6OR9pM2GRHzPhLsCpgZZhjac29iHB7Xjwr27lCaLuwH2Ldft3wnVAswEt
caeZJ2+ix7W4+nQnKgmn2Wxt+DzPGJEjGHEt8Rn82yniRe7Ii+mf/IwJpLjTEU5nksZD/GUZ6O1v
BbAgViMDgntgkc389KLIOpi1hDqeHtpoEII9G8bZyusUfjheMxX2dtcNmku7is9Ikl9Su7DzsVau
U0QwBSCSmjm2e9sAWRsT11UAzKqxaTJHQ6P+rg+GeS8NPmVCpLFXeCuMKyWBO9Mj5nhD7yMbm03W
QpvgAATV2MhjpWj6pEBQHX5zLBWrFzRvmaEqL0NILvfMxXcdor03LIr2S0itaVMfTG6L+SvswI+W
s4smLgcgTM8101q9PV9AqQf0LBaGdwQ7XtmfVm6MLn6JD++yG4cOLa5Q9bgH0eZa2kdjCtNL0e7r
PnpohVld9OP1Sy/k/XlklbQmdT2jL4yC3eNdVu/7AbONbbdO8wadUjrNcL3+fZPTEH0rlx0ZhrSk
jd+xJ/BYzxj0Qp7yXfxlq1he0tW1IIrmdC6lAOsmghG2Cg0nBjsoQsnT5cFbb9w1cUNFr3GSoTkg
lcfSC7pVodg1z1Oz5Q0D8s7NKbeSALwgG+R77YadPB7ZoSvM9dPHE9ycZHzOusdECp9vl1m9enrM
6oxqvV1BXkRnBsCEnQcc8pG9RvannkW698thESBbB8wvhjAKFDIxwYObre7+YD0RAJ9MW2LvF42q
AppdrdavNKPrMhKz7zmnzxjNVgP0VoDBFu5Fr84U5kNiAlJ7aIyG8SCeQo7JcSr0fTtDbOWbywTi
qug8N5u2nXkeqt8KQTc7ncPncyA1fcRiop9lk9cAH4P5IkIp9Eqydp0GJDDC1xPPWTLHI9lO9aoK
uZAk6LCdjMDSKYRas4fiY4KRiQEMSorSTKPzuAxxML5Bx5cIlz2ZMr/TAKBpyWFWehOknzB6Mojc
MitQ/LnRJ6v3fBqPfEH727HBHeUusNf9rq9vJ5/53YH+PCeyQmTc4nbTnxl2GNYG8ifBQBRb3Kv/
bEd2QnhtGaSN2H3dpcTm1+F0t8anUUGYGUyXNZz13JbepC557nKuIBIbMezTD0iDQSGVhSdp4QHy
8UQke+ovzzAOUzEWZoL0TYVutIUuTHmkPdA8FNSPTBJSrx8F9FxNtJHFQsW4IrUG3L9K3gLF97bs
gp2A9NK3/Gim6wyrMs9pX5h6ZSSgFrwr+nsVB9hB4pTCwusCQ/Qum+D74Os1+LtWnG4H89/YXzJJ
I8vaZFBdVjwBrVHhTuCgOpsP0yx6QbypaWuYcpPZj8Fl6LKGWUaJ8o80hmMnpiVZAMWEsG10+g3L
2wwfSdFC7UgC4EskaCSzQFiZ38Locgnmtx9o1MpkPtWhiYMgdSMzuWv+Y9aBGoxQbAsGsWXimhcR
IgJS/QF5rF3heEPSbwv3Mwhf1/nb01nriSY5KZmVO/UREfi+Vul3+G3i22cIx0kx6OSzXsIPioCh
uf1UoEpJFRGXD5B0Bs/2dDaWtUnMNVzIovmT1VLFsgs2yMJfhipfAPhMNjZ1UM889ZBMJHrU8JbO
YIVtFzfJKajqeKimiQ9vvzOULQK0Qr+XL+Un4Mo6JEL44OpDSjMesALxpwtYfwPZBAOZRLVcmUc6
rPboAAoTsfIWy6OH48AeemnsP/VeaCN+N8rnY+2ZBndmbaZrc6I6cIYJAjqzSr+7r7CVYh7ABGSt
A/VQ5U7cb/gIKFDyC9HOetcLX7YrWOsRrH6Ao2NHFNlYg0ntA+UZ5k3K/nATvcJKwIeEPf+yTnSY
wu3aqQ8leoic4tv7IoAwsdvxBpR8iH/k4XEpN9oTokFapVQqioDjdkz+rGvbml1+cHn0o4oD/SfK
bplrw/+bLLdWj4hMWPBKo67l4GxZyrfCjUJ6qujAI9UXxayUWaB10iHEhYVys57iaVECSkRBsITg
298AgagGCKYm/JI9BSfdh2CloX5TddtFB2PgUEIpzO7FT3JPM33n0Tu6ejklkcSoo1Q+tmptEiWT
HjVnBNEo4Iov4dJeBjs9D6xM7cqiucGzPts3HByFtbHNLi+8OFJLNl+lRzTQNvgoKGIGDE/puDKZ
SDHjeZ3EswPEV5XmBAo9Qq/ZEHD8Rctdoa7VwxpS45ugyC0YZusJheygCLOkpod62sK85NZvUcnn
DR0uBYYvibklJKEaBpaET6/ic+6WY7HfXPtgFi0Z7PrExh8U9qVft/gAdVoEeSIoSGKc+jccHGRS
KetNX9aNzngXHOES6S14SZRq0dSsPBXIlXG/aamxJlVGJ9qqm7wDbAA8nKChprRCbJ75P9lC7xLo
pUUw3mJy+kOEtSE6r9+/hei44H2Rf51abqdG9v1vHKLkA+GcjRk6eu0JjGbzfqcuFEFYaAXJP0vX
Znt4I39+1Yhzi/QITF3etvA/g/nluR22YscNErbYfhNlpW1/imsmYyjo35ZPvzPY+BMI9Ati3kAV
scxu375e3gvPhd2WQ07IEN4iOiUIyCaF7hQmMaMGPjZK+npUxddcw1kySfK0ZnA4U8S9bAs+H/9s
YGrdKe27zNdeCHn9gWPFCTPYQMhEZ1zmGlyAwFlozVuQMee3zN54AarPbKcdANYJ/t8QhXfEZedl
bt/QwC1Vh8ht9AZPUGN66LnJ3n98jsiRXFoN7iNrN09wl2AtaqPLeiR6GD4FDydmDNM9R1Odp5Tj
248kq0/ky2NSaglgK1eYfCV5s0jBtQkYb8NYPZvO8RdhHuKuGF7KXmXwGLHpepUosv/VAN0+6zxc
wLeqjo9lMAfEoXVjMXto5HZrrH8PfwEMSP/urbarP77uAvA82nARN3a0Pu/izXrfKGf5GjTlPgeX
uH0lpEIYaBlsyWL1l1ht1+X/0dxm7In8Bh5o10DPfoWMeNv0ecno5z5tax9dnZKafdJhLjm2eEfH
MeMMdQP6QLlg92NmCQSmFh4wyzF9zu1ez5XtDXujYQWUFbkSAjw1qfJhZYvmt8LP3HXnm0Z+Hm/8
ImxYG1NDihI7pMdH9dYmxRPvTPO12tTmhPt5VhOjBLib7OndLeVpJyF11HqiAL6hsWRQN9TfACpe
znm19fvKbhWYBNiWVXUpPozMetbdH6lSxJQAaQ7xeHQdH+ioAIejFCeD+EnK0yzTI0496MgSigxG
ec95qItGYMvLj2yYbjIoFwWV1zbnjjgF/oifppxDxFZVFal+uOxGlbhxS30XMdCC7VGdgqzkXCUy
VuPL9dvWDsW5yM53+72CJuTmcH7n4wV47HvF+GBUTpdPHcBiAs6ZZU2jt8hh7gsxCAjH68chR+xg
NFDf95U0DjKyK6ndEWmBkW6SqC5TyDdNlzYiTErnwzC6KSUlDW0YZjCZOAiLYB0jeqieIeAQh+Ge
x40sGKUeds/usFEsu2/Wb7hsp2moKTg4GoluffVkxhyQIo6yI3ed9u9XFvO15ZPfLa994LnVpSmx
1sqIqkC2I6TXEE8EuVvi1ejTYgauVxJfZFce/+k04AJt5JLh0E4OI132mcO5Sjq/+KpQXMJZweUB
Yuy/9wPs8PFTDNO4ewAMj4VLi9owZ5Cqe3Bp0ZArI8Pwua+x4CTeJF/sDnzGQfM8Exhs0IbXM/Ju
nzXpJNLBpmvxRfyQSP8sGWr3qp6F2Fgu3lZ9ckw5HR970nW/7pN0xv6OcasvWlsW6XMeiDysVIZO
UIoXhRaPp4sA0LOJBsP19+9cttwkc8FO/e8OB1DgzVNmiKdH8CHvBxJRSKhMCZyGfQZQ9zn4yYM2
WAb8p1mAytEuDulIs300FyIOrYoL5Gnj02RpD/GUSeaMnfd3fr4tEXG9dKBuovlC8iTuMoumxFAn
Ou01gQ5qTL2W5wdTGB973eaisiyvf/q9AlSeOLc4t2xD5/W3Y3z0DLvWjjCtpY/GrAiA+7/Cumxy
A8GTopNOiUvIvxzY/ge/0R65zPrpGVZxQYDfeqtywjL7paMLqqR5qAkjP6l5zhLzKFUpVIDPmdDe
+xYlkDZwCvrKRJTdvKHdYtUVTe0osUwN8sBqqgoo39jiNSxUfa5LEktiEgweS/LwnBZvskJFgTzO
eZZJM5aZonynPYF8tBmrGQ+d0a37A2aD/RXGP1lC7bHHklSsv6tZnh5tyLkFej9ujUkX2cCymlH2
7coVSS272VhRRzZG8Q0hJja+9wMe61CpqDH/V5dzs0IQnobOjj9DTGBhGXRfgH4o909pXm2KglT5
qbkzIycrT92rvx0k9DVG+r2CLhOpaDTX6YmojYtRQ8xVIVELObYhquscM6oX94FphqMOKy4g5Zme
MgEbmwAjWkjrD3iMpxdbr8V6Jwc+2REqIGnOjYLCdsYA8Daz1HkvAzvBcOBNYoG9UqDGAYDKuRGu
tT4+MTK1BOkVDkmnyFe5DVXQlbHhNmVc8TdWm65tfN2ozd5vd+mWaIyRZwKLrw5+PjaTIJrhJkG0
GfujauT060mQs1JVTuLefRgH56J0SUbnY2T93BNjJpiBepO3F9deMD+FmugcSyYmEptz44Y1Qv7I
elviFaAQ0eo2NudVM+86yxS+WbGHYKdpf0DBiqL+CG8iJMjhoBLAKDPS6cA/yx4nAO31k+hv41IO
qtGWEOJWQs0hA3WVKDL3SYw5nI/fwEI6R1R2WsYKNfKQ8CnpSP8Vh2vANc55Kq3wV5t1NNpBBhpP
vOH79Quoq14ZqxnRI9VgV08Aplc4driec38Zsbvqm5aa8pAFCys3q5wuNRVMvLt2tVtlvj2SBGIc
GlOCsIga/Lc9GTwaAiw6ajpJRyPit9J6/uPyO2lAHIsWRqUgCiubWU3EGWip/ejmNZXuD4qB5rD6
WGEVKmNlxesICtPZlHBg4df3LJ0VAubgUpt3dbdY3JY6AUpn/5j8qkOQJwszdnfrcOB4Gv96srxd
otpmwMymk9rDIdp2aA6qlbIVoTGMbaeu4wOPXzE0aWUhWW4woCkPtO6siksgXsaPzVqqyumlKu1L
XxLwQnF0J8E4tiC/mNWl2ncyyq5tO6Njp1geCG03lT/Dz1LD9Jrk9OrYErA3/o7YL+XfM8H6izoR
v7Eo7gHRjv3T4aaWWhtPGqFJma3vuAblIK9spyt2T2NiVU4Z69v34JPsm7ot4dUMyYFmSngXC28F
eRk3rMqsD3AmVHqVPzDPXJ1IbUc28yCb5ObdSo2a6x2P8+K5eQobLs8XCIDNTkpuO9Ebf4lq0bNs
2C5MSpKPzBVQzBCNsWFZn7YHRXNeBv0J457iLq34yS+K6mN1yG46CZQ4/Oapw6OkWhylzdPiUbcy
gcdDthvtNFInDKVur5/t5DArz+QOw5xK2OwMaaKW0MEl9HNuTuH5DZnOWYnM5dM6F55etwg5b+de
nqDVg0ea4K+PyZSUyermqmTMvPMZvSol9aAlWk2nUqkxVdzdR/7+5X0wJEezCTba7Si2xhb2hN3J
vpODIx2dz/DHc/RIxnhHiqtX8FCTiZNAW/6vf4KvTktMrorUuDYcNumQvF6ukks9bZ+N1tH1GyIq
HDwG/QvFQHuNtA+LpphCYME4U2NN7iYyuVfLvyJV6MLbAWx5xyM+ZObjWQlF3I/WoRi2UupwIm3Q
IoEY//nrMcHNP168CtaOpH7Eor5sg2EQ32VbBWbfmjy3hQqgIW3wcE4GcrzJRamSqXndM6ixXnsY
HTKyXLkvcAh8PoMivh6fOXS6yvBOjoyMCT3rkDIQqBMfDExIAIexP23qsctdY0kpS9EVbX2M0i46
fOHTNoM39joly+oQrOM83zNsXdkbZGTp7RVhMR8UYHHC0NEkJTHYDArevClO2IyTBN1k96PzfKNI
INxYfXixuP087vZNWOEwnOimSpa8jBx4w6hfxwYJ5KXyGici1b9otUTAOxgzT0r5l9zIGk8jhswS
qoO3zVlh4g2Nl28H/3DaM6ZCAUpFbzlnLll+rssPtKgvJmNdvt3EbVtxJkY5ZtZ5iconnESfEkiO
V9cH2T57AIqvkssHrS09IEk31shoi5ya2d93W5WnXgiJoPlDatTlZngib3vzmPubGkk0TTJJl3qN
gfUSuNByYxGq1icoXmECWa97oY6y2UuYRXlaQDZ79XlvUdSEXbb0JT5FjRi/U9yDUfLqsZlGHBwx
JR3n1Ti2/urS8jc3DN1lKNFVcDIy3VMzoat4bVGiU9TO2DQysbBJTE1wFH4bqS7UqR3X23R4e2m+
mYdygqRnEXY9WZRikmhKkU0SwEj2tzMuR6u9KGksQoo/yGnPnJIWUWVUdwV7MUyMNkYEVvlXolsN
teIl77UiFcHo0x+pR6vq58Es+A6F5zbfCiVG/WlMQKRmhv4xBy/6e8zd7euO2IPoilPQpCh1WCfU
WdTdBpphVlUHF60oU+ru0V3s0xOQ7IMaafwTvXerqgq3D/JEaM2B3jt43L2LiVlvbo3yQYypTdoM
nYXp/VTbsEBXwvyBdljM0fP4fAYkoi+p7b8mF1xsIqZ/8WDjTe4wzHT5O5zTabPZLEPn0OCSNU8n
0zkGV/6qhuP/O2EbB7k7GVrHkd7K7dMCHIcOC/dVlUwlWjo6ABghWjgXldGcxQDMNwBEjBiAyXhh
arxtH+8uAaY35he3i8U8/2kyNtcHc7tMdWoGutEouWTxxR+j4uB16BwapGYn+bRfUliRxtgoU82E
PFJ+z4YMEX6d2ERiggKjREw7H7fLuA7jjA+X0uqZ27jUl1RTdq6kf4GNf3/Y525VO1fMJZrykKCP
dMGCBIywMHUsvfM0Tct/gqvon4zbt4w+F+oEotzIEPkKxNZcNza+1vIGJQiMRWL115McrJsf/D41
meBXIhiFAZAhSlgKd0sVPVH3OmQquKzvYeyMuEp0OsYD1PmukgwS0XhqoFgpWlf6ME4LN6LuHoES
+kJOQh4xPQFe2rPV1og0GIa2dj6PTfIYJAcj6p8Xpsmha8xZ/0ojRN35bH2q/IJpol+Q0H1I/qOc
vWsFq7zXXk+VddJyd0DFjTnsUgQgbQB99det7Aha5z4A3Nl8EM6HYqOWroYz2SvCwUynI1BNi85x
NA9KXu7+ckycD8UR8plhGkujRyx46EcanpcqPCs39/cLcqceD+d8QkT87H/YFuEdtCDK7yZfufdw
Kvyx9MN2cEd+KdJFMIw/YTculm/IDnefT6QyWuay7pqJDCbAl6R6MTWMgsf85YvG7FGuTNV4sQqQ
4bpthXjD2D+v3EUm3YFC3zOiOemX1L8p1kZQOU/mAfVI5SE0e7w1qaViHoo5sE4h2ug8DaUZfeVL
oHpbJi2XC3+HlI8v/8N9FzLkBm3zjHI90XnBlDGZEBkuvTwa+RZrN9mZA34twEOmmy6UBUHToPcN
XA7zBTDRHrRDy+WQUr02UBRBb11kcNy4YmPkMSbwAp40/gQSZ1m/0QhGx0n3LbiaCjABZRQ3HsiT
R4c9HxUbnc119kQzd/GUGKGzh/+YSUu/6vgdfu6C4+u+hKNmKCWantCRsboeNkEiHESu/WFSfsqc
CY2b4Csq030NONHa9Fq3Bs+O3PHg79FQzCaxlevHiFTBoTuslFuPhERz1DeLZv8RD+4tgOE0wrls
ynHqQqSsktbuBLTOiJ6LUuor5OlqgoMLdSW5NQBTbZxyBmGh+d3guYUSanZ4ZistqPqNA68UpDon
R1ATwqzsnPi4Q+r/zy5yE+OuYjBa/whWgn+BWXXtoQaph2K18YYORPrpgvKObvBM3F8AwFXf7CM2
VZR7NSW5t9rfv8aiw8e0aitXcilblc604cFe9QZ3jIKFk9XTvD+FyTMp3G3N1of9Sp0ngYFbvC4b
WlXnrP+w46mX3g6YjTz0eC4fhdydb8t770VyYNFpWhdO8H2xZ8+mhHMYbT37aQwCl6byJJsC9MIx
kzJDMNksvZMqhi/bhuUdIdapuMQA8+/Q7ahXeuCshLo34VGY7BHD1Xz6uc8mZagW23Hac1bgFgme
jtCjJWfpiRMqMwhlp+PY7QB8ITX8V2tNDaNOWh5DVzCuH3b7TGGP3lMLo+cHUHrW3t3nirLUIWLW
cwI7TBuQ6FYyNFWqtcu0BWatLyn9fJWIIGBY4VnbZY4o3N78HhE7rZktqwiaKHwT16Qsq6GhqHWW
0L6H7ehy9cbggz0YMHen0gUrHw0z2f4AwfAjEEr6W6E5PBzYTl0d9bF5xzi6k4TmN0fFa6/TZMc2
ld5X2Xnjc1EM5El5Wc96+aLUWtiVjT3TkMQbhG4OwtMrJ0b/TcGHB92VxTHfuqwQewEkHYRLnECn
fCkSmoKHlXMXCzxGXUWUT8krxim+UeR/V362H4/fsrnIicb6nwq7aq4IT+cK69xp6SluGQyzgfrb
k2+VovDM6nWonvbLh6ABoLDBfzHB2R491TGndQeTZhLlsiWAXCa4YQe47JgXqmcoHMyw/KpxK02s
zxxLLQEYDoDr2yE0OjP4oPxhlfwYSJa3vUlrCNOMNeiBufJXjSMq6LpRqncelun9lf+OLtYILis1
8KjXEPfN6cAPTGJ5eaz0oiK+c0PsK4USTBfnlIPqfn0LgekO7Mc3JvFHHUe5bJegfs8HxCU5WKIw
Q1tFttQC6a6i9B8jQbjgNeSoWSp234/ZIaxdhJ3yLlst0O9PopbXh1f/A5MIcoSQAxNEkUBgQckG
hdmK9WE1VO8oe+RbhRLbz3vdHDHxoqHMW+mhitdHu2CQuLME5FQtBv1N9D+VnXtQUE/hmEZ9sPgM
uaIV0QM2QmDJunXdcHPM9XeJI4uAfgIK+r5cyRIFVYyCmKMLyGp7DxJGP1FdUGiQwuMZnUVMIa54
GBxvI+3+BEdMFW27Y6V4snLisQxGvEeXXGTayqkwpAjC/4Zm89PW4NsxblPqZ3WsJj5Qv/DQ3RuZ
d7VRIwHV9N1Xyj+c1IzwK3VtWNYXHuipHUixax0k5nMNMgGJY6+IQSPCpK2BoOjA/X9b7id1u+M6
h9ui2YyGXYDrAIQQE+DjEbUid3lso3WHWU5fTvrfNl7e2b8ieJjvOLS7GDxhwOqMEMlufktIHicQ
QaebIksM96GMyeHS7LNloZUPe0NWZOZS0kNu4DgJ95dOHn3u7D3UUEfGCmc1NDBdzWk9/Pldj2VO
BQWu9DEMWBlLp1dkrABy0VtFSLsktcbZ8A9ef3O4RV/8SkuXkqgGMtEHisdCDnUNcGcIdO8tKWm7
Rrgz7TYKkCwxMVwVN0jmBUGuJaZJy96Z1/wJU5F4jWOqKWf7mpdfmZOv+3rflCpttWdgwszYXNbq
+bNwuv501OAxGDMhNyhtCePrji7KRrXEufjIg5Wqu/DmgY9TZUszh/rvC6tR1HC+68dLA2uQparp
EAsMeTAOZmxGlAUuOe7dR7Ks2EBvLehqNuj6p4igX05+S3d0hA2yPSjMDb9iongxa7rOqAHxlMNh
2wa4Mf75QKgE4LneLHMCjEsGs75r0ZOOfm531OfFU2IpNGQdO7zMLZbUAFnol6Gm/5RxhJxSfzC+
FgGhi2YwPlnPvH7h4JCNqOym9JmOoR3hO15YRJAp4oGniYDiijSBiR7KzQle1PPpDFjoLHWrEPSP
dtSb6pIucX8ZJMz41MmaH3JwdfMW/u0dI9v735/GWbmHqMotVZtEs8DY+RUuiHqc9pVRPEvjmeMn
eZJG6cq2qbISGuQQB/HXId+/T0ANPV845F/7gXifLn/VZliFjgGVpLU5iV1PqYWgvGTnHx+Uf7Wg
2Rscw6cvNhAppyaCLBJjd7WoE9ztMlaalsnj9FR8paWjlOVW98E0VTPWANd/CGKrfkocYfOV0Ppr
vQefx1zkf/w77GFmRz6NKvus+u39Ztwzoh347Hue1HuznvZa81jOtdN7JGfZxICzro6hljiUurW2
E40w0K1HugHV710CDvt/QoDbhZBTDU15rTSouMvf1g1V+N8YJxQGs61gbLuuqvq2Vb+0SLlTREQs
9VxKW/3KZPN+zlGpC7SSpFUgVRrqUDDKSB71hdzlrR1E1dLdrwsNpVAsyHBuCytnSiL1tg6chEWm
Vqs2EvdKSe8BpDsbLuV5UThmIxG5LqaUdfvF7JTE3btJV+KjEsmuR/YdSGZj+DxVoSG/97qJ1wU5
BPZYG1APgRxq5yJfKXk9NXwYDXdOxX8Ye41A/9c4DuUHvQWcNPk7Vuz/29cVwo6OCTUgjZ5fwmUu
Nns4ESFGjtFIpbgYlRPtZ4v1hXQMCehC+uMTn+Q8a/vr5EItOetIKYD3HeJARzaTvWsdblbvWdW0
iHfiyr66UvTNHNbTrgF9v4SDDf2NZrqusXrPwKNfe7xSaoZ0J3TPOw0WlOKTv/QyTSVHeOex/7gs
sYCTO5/JwjKOw5JFAQqYDydcCLPtFk8sxhJsnA8PBpBt7SJt78VHnXyXp8QU2Cl8hBzyoOOQLV/0
ea3pdvTeHhSqhxnoTOjBoQL2VgkCqkighYYU+itCl2cU/rJEO/VU1CMo+Vqv4ENv6yCz+R8WCOgE
izGAbex9uB9xrH5wAqhKQAU9w9f4Ox9vT9pcl+rj5w6qMPrZDWLCfwn5NZJkayX0PIoCBko3zBO0
aJYRdjuVkQOYUJWFHOvQOj3P5Sj2hz9CZxeQIiR33gEMVsor2rU3WT1rHPjejlFLeWwtIXl2fXVb
qE1GhXkPMwiwtL0dHjS18WmCRhHKye2BuJWaYPOJOwdSP90rQBRQwuB1Nrs16NIep/mTmwc9jyYt
I4pD1JQ7om7IHwvnbu/00kpR30K5Qom1xQuH+A4Mm8WktRpY44GiUDb6Ghzw0VstcA2AdAX9FFlT
7fY+XWDazqonlF4RxT3hRowV2CKnEk6qIci5z+9Vtwt2s9qkhM1gNZJw7SAYVLkanWbGmNuno7oJ
w0dx3Pqof1M3j8TqW7zPjwieekspbtGcXo/yeHSrTrJbr0tqqKujhmkknaagtVm3U1B9zLCGPOow
8rQcWyg6E5nEr9O6QTOY+T8YY90ccHU9rPJvPEZymsoBIR0lYvxqIyUQsj+w+LZ71aun1yQxwNfC
ul3HCHRDmLm74YIM8NzXB0SxjoDJFSga3O/NHyaQf4JdIdYr+xy6DY6lCXhfCw5RHTi3CUohvz5G
ZlXH2dl6QmSKaM8AB2E63AOEvEiKMqfaa8NQhipixv21S0panGn/GA+BHQoK/E+jHqHmQBdFy2GQ
cDQnqaz/OL5JCqOkCsl5ufHmsfOdxVnZs1I4wUiX4T8O3AylOc5W2GtSWW/c+gJ7hY9DGED2Epq3
+PRjMkNp2HBkk4+AU8Oy0Vk6zG+SEig61wWXrbmb8blQZ4osIvCgpA8FaxVfGeVRwKFYMS9t/7jI
M2R+4p35rMwbOVyfwIjCWFfxXtcn+FhUKFRXqTQXtBVQ2v5SL7+jKlTRKpkgtJQRpoyR8dUUEBoB
lymLwJqx0AKWb1f4KGfM1InXHM3b2WyMpZvKQAe+zrXvLwNDyRQdGyQ8jOLQW7AfTh+uJ8jXMf0z
gielVpdqk0ebJZFlc9pACzq816urXJqKOGYKmtRKUXnNkJImOPVZS7EQGwKGcN7cdX/GJ+mGBgFM
iq7z23Db424JLVYUducA/Fvo1GI0X+PI1DQsN8sEzhx+zxT2g6vC2j2Zhl2P/sxJ7xr73VQp+Uv2
lFnQo+kiLVj2uub8YSvDtqEzQrcX6beNVZt8zAHVO7XL6ZDouWGWPTnAlH9Vd0kktcuv28mv47tF
Dv4GJrI3QOhpaPPEKxf3C6LU13nD4XBA5lxm87K7Vi3lGM398BVfp0mDh9MTwR9d4GbC+LSB6bFR
NKy/MyrkglgUz2bWA7iTdUXeFxgtQaJr1zJUSPiK2HQhd8vR0M0o71LkZOwNxQAoXRqyKrgpTU1F
8a78YyjICo6tjFvCkOGwxdMEXIxDvu7+smEIR5jksrRprCBrUsiGiixl1GFKPFiQvtpjQVuDfg7h
zjwZFSeEBeGkK9cN9Bqh6hmslq1APmYmgLgJ+3LU7mXOw6Ko5TuLn32BqMXKzUX1RGeSn5L9Ne6/
yQi+6WCQ6Jp87+FwEz94PZWq0SrVteZVElVwt5FwaB+KAXdeKJ8EQhp0Q1KcM7JKNxQzLMNfMhXi
Gq0lLXB9xOIvge5zUEaZ4cTfG16KQtJyCrFj6rvNv9HbsB7InYjGrp9inbGrAdmqcP+2noPsq2Vq
oq+LmfYjd6tbeNRPm/CzGovIE5mbfOCY+CWC4p9qf8ZsTzB4zo0Hiiu7noUOm7riO2AfwZsPH0PU
UpKoc79Vaf/++ohX8Yl1Ken4HqXEsvWvHVI2VqlgaQehnhPYrlCJl05k9p6vIKK4zKtUjTckGRbY
WT6aKSuYf7MaAVTFsbnu8sWIBzZAkSu61ptR6pEkzQsILFoGD3UoAw46ssQebielk0R/RA3s8Ekh
LdE7oJzvbk4MsD6kqfmvtcRTpXp3f1ZOvOVW6Ls1GtzTXhHkCyBxUeXXNeUilUu30Yblc/enX4tX
JvxJnzaH+oiwuRXcM82gTkDTgPwE/a+JEntYtgGp+ZcxzqKWyW13YVRx+SA4xkgRqLWdWY+AWMQU
GQucI3OU0OzU3qQstlr0+OHJm3dO+vLCs/eayeuq1becPm7hBJBevVHItg872LO//afAm1lSJD+Z
wZT36R/eJrd1r7ziOn5J0dmiXh8r1juTg8nRha+JjTQJP3XYbUO+IhiH3Wkl2SjZQKkVied1OHua
izTH4g7tELimVk/+wKt3FWunYNHMmF41sB0ET9Z2uRA8eEYB3ypr6/Adg25xaErj+LU27iuzAzzF
ctvcZL077wssXADh6+/q5H6Kl+WchNIsQ2RPZ/kucODuBichcRHyuAdrNIT3sb1fQrQy6xhx1Esx
wkS3PS/iPE33w1YJb3mPPjWYEFEc6iYQ9zGw7NdVwUeyjnOb6oSzPPHxiXZL1xBzTznbCngsvf5D
XnJA4LDV2C2rFf/CRmIfs7DqUvPRKZub2RFRNyRpcO1ixcqEti0PSqx64q1m8JlSv/jTHmG1jGv4
TKkttXZIV9QQoMZNLm+Q1crqbc6o+xjdInz9fYETbzqImRZ1fY7kRTN+ltze/RfG+CaoulTTpGm8
1kFroYLfbcplJ4Xv7V5MDFa81+yZP5kYkfj4vtiW3ESreAFmfuuCIgHCrcYJHdspfa0VfzlHuiGI
cCfbt+K47wtl/FbIXkv5ZedX/CHZP9dr8qqC18s1GGU6ut3ZfBUqS9nWSD5jvFnLsexX0mMHSWu5
5Mxe+X3QUHRYGOsDomV8QDmuya036aDwkreMjYJ6ZsvwVb4nhMXNR1F4rIspmqwDMbhmlmx4Hoga
xq3XiHIkmKkFTfpcOYqJlHGtthTbdCziIfbwIWJh9sNopZe4msJ84k0nJuO3IwdWbUxW2DnSITOK
B9q8/2tDEU3eLCG7grq8aqVe/6Un3HM1oN632INk55CU+bCNFyxGcvBn8tCcxcqEO0FBm9yOYjMp
TkrRr8szEJirv3uAZG1BK/sc7F4sDx0DHxAt54+jIiMtuYUfRy8iFLkBcTG+wVS3kmzGln3P0VmV
+FAa/8OTNVe5M/BWqsUKZcRq1kGtf9E9N4Itl7S80fksqp/9trK5O2Rxb5zViMw9yB1I7diAhOp2
almTlm9rC2P+8yRP8J6Bo0gK/0H8erB2QBycdOdP5Gvm6icgJHyqTmywIIpOYYbsp41Zj2e+0rlt
rJObdMxMO/iCLvxzgYv2Vg+0rMT+k1+FD1xlhteUBMHeK1DHN2yFLMNiuQPWUYuCIwN9okZOv/ZL
zHfOnzumxowEp9axY825n707nOn3bcLH775oq3dzMPcJcL0BTACLdgB6NXCJQETJdBKYmEZz4D3I
LrLNd0mR1DHl1OKOIRUMUmRkKX9JXr7rE4G9gMM3bBIcWhpvAKSzzuzYjZTKLm3tP7au0YMhBguv
SOEwRuec+MhZYCNPoCpW2gem8esa/eQi2JcGnIktb4N6luyHmTyW82QUSk1fXhaZaXlDsRB6lrKw
VEEtYuSQWaJY2n6STgoYpVQ/e89fkJUuwmjdFNsknNCmyE/x84XK6Vb85zr28Tkbhw6Xv+F0dN4Q
WiwIfCOHUk7/xOuvAsGNHGKph+GTOMrCU9Q9w/1wAgLkVlZbA1OtwBisHaY8e7UeHnT/zrSJ0Mez
OsPojDd7aCoOjIMzZNpxxX7sa+gU5GxC2wTy/7DHeqAIU4dktsJHHKBCpH+eb0fzyKFphZXQGP6A
fYrenoeTMhK9pQdRYJUyNCcaEXeEgU4RlCLd7Bp0elMfLYbJ2JGB/16UFw+r7nksMOIjTd+bFUhQ
PWllFlUDjRxFFuKh9n98s6Uz4OKpAOa6iu+wq966AfyGA3XbJppph1HtAaKDdHDEEsaubb9SKLMR
2jiew5K8o3hf5NB1MqHcIfHNgN/C0gQXty0qZFvTEZ1ppxDaZZTUGaQWAoW7vSGZFavWEvH4AdTc
4XdnVqr0+2NjHAbgVsHfmPictq9GhSOC704OeUNIF3+72GsXQqxfDTcwIsMuPiQKrL7TK+2sKumI
yP0ueyNNaINBsN6pqVNxm5m5WcTmDOTdHyxSvW3UWY/jDEixswjZAMxhEbK94OVYFWTaUcaJ94Op
4fvpvzHqwiPsLIQ+IDKlwuJd4EVVh3H2BxecoBobVfhazfkh+P4+tDS0tRiWT4mW+AipVMKyH5Uy
8pGv/A8/Ay5eZ4QibDFrDVeGoSStjswhEXxUlr//FUR28izSOhD2kDEhEHfSXi+ZUGCiuCTbC5vX
ExWJyR3wbUCKhMEUCys1dot3dtZ/K6ncwSs9UBYS3l4dupsnopzpsj+LvT23FwPYUoy/ev1Omk8G
iMA3nW8I/xPZXLtoT5PBVyF8ZphcsLvdS1JhyA1XHYLRdaaBjfymGrtLLHwwe9HFsl9qifW7gecL
MA2w/6lvQAh0yXAvHfVW8s4WxpYfEHkwtxr85CpvRu6I1WIog4TNZV3u3Ucnl0Ql+9GkHUwRCEFC
p4Q1YaTzCoxRQX02ORPlYqfqiGTtZ0LI6LBrJYh2znE28RxWgnLthbGKjc29atsQZ0VbLtD1uOxU
2PoDYWqCsxqdpj60aql0+ItzcPU1QJQtl4ilt4i1bVZ+ltHV3CjKQmiInblk7QfXi86axaI++aEe
YKjZT0ItQbvx8M+PvmhNXTiU1Q8ahmdtOKBPRWZUFQh9vhpbYUVYVtXfl5SjcP9fxfTDl4J+phx8
CR1VipXoVRIQy9+6jjmOqqNH31rpmFRFNWqMuhf6f+FShFArVzDVebBo+mOTp0164wsI5OHPEa+k
c7vJzaGu4jA7oi6sJTqIFo9ygF+r9UizjavTqcByEzUV/MEYuqHFWuryRx3eDWriso9TwNFsid0A
E1vwAz9Kd4Z3/Mkp6dnlWf3IxBPlUVLmEqp/2PNruRkALvPjg1wcucqiKFdFW15GIPJY+xPDzHSA
SFw0/OFZKIpE5ql+Ps+zvXPd5hvmFhEjgTIE+HvWQTuSWIgQJ92PAMVpYMthh1jNEDoOiRaqycA7
ptDXiFsCQv5NMJYtJm7Xb1Kq6V22RbKJJyUPkVR0com+yXE2KJIDYs0mUt8jPR6FEgjSjP1nUgGE
peDGUR6OBmh0Ike+ptXvHzS8ZKgkq221Sx6B8V69Snvkfa8jP8qqCqePrPgwdB6kSv/yIhq3VH8d
nqaUXP/fLvOQkx1y1XT0xBwD6QbkA5yzbrAAva4kZmDmMLiyKbfDds14fe5HB9epwd0P1u97QPyd
cUpvX87JtfieIh/WopOGwxK7oDRf3X1nLZGgpBxJc5cb45gfmr8C6D/5m2CJs/kaIUXGblcrXbkC
BbUWtxknHkUSl5reyOuBJl66FDKDhjQr34RAdmS5Fw1gLnY+kiRuPwqfO75+tWJDQklezj3PtGPl
ipy8dIcUTXOGbvXVsKLelodplqkBwua1BSnt5s8ItX+nWN+gk3gEL1jCXp2syVUjc4bTqoAk/Zfy
OR5riBT973klTsZE7MLBB5kK+56xf8p2kzVz1j+qwxjVHg6RGkRKWtU5Fey2QA6cW8I+xfMJEGi8
m4xnI/1k8zTfZgJ/MVNVNPmUR5Av5Dq2NrG/FPGXJN+wi+ZbmqA0AjMWCg/78hJZ9h9x9o1uV5/t
k954dRl06iaY+eYRvXjCqptzcYAgH+gCmqMVI0iJ13fzf2yEAuipV/G0mhfSr1sRXk+zgFESTW6N
NvMg9G7mWXU6KBu+PoPr/xv+G/qnHLU6qGu39FlOzJedlW0U5RCdPwWhgj+uyb4umkCCamXF2mwh
vwBYj8ONPgM9awFYtHM4Cm35sr3FgzLolOqSFl4W7wjkW0XaofY1JJrv/TrGdEG3Mt0XC4rW8S/0
XYb1BrUgsBmSJ8aAeWI6Ewq3PrY8+Ev2hZGN8LZBnbXSE1qGNuVpzfPQsRV6ZdxujdmI56zq04DF
XGJO1J05XV2au9//jPsLiJ/jlzuzbZFCm11gUvmx/4tahyyUCZADkZogh/Vi9aeSQididzuw3efX
RZad7o6IEeqEs07UA8lpTSgiCENO09XtoTlfSuXNma5e1lGZ6ahTucj7duRhwLsM7WS2EsYMD5pU
yPKS8u2rz4CsxDflxbKdP1aybqd4gXLOSuYxJvq13G8b4xyMYBG3J/zBN/xgr2gLaCaeX1kpAllD
VeWeaSYZJU7J0b4Jw7dimlUHbOAyUyN8gvs/25E9RWzbLLVK7oIG+V09dnqao1k75qf0Q2FWODNh
PzKHmDIBDTe5C+M+5nx/ZEZAgCbrGOylV6q1Zm4+NT0BXboZpnWQgq9eByYBfXHI3hUhOLaZx1Gp
TbXULAL9j8i8oGYLVDujYsCAWbPT3+qkWP8xNNJ2jo+bZ9HdlXkZkNJPBM8DI5oprvbuLn50zd0X
1vHZb/4N9dw70jDSNn5Ze5iNpNuKZLWG1n3KSJa9dqr/mX/bPO8DwWvIzb78RfnjLeIYjL+TqZVM
HJW4r8DDmSx/DMZUwjGynunjDIeL43w/rUxJWGsvnJmH1XKKSa4bCZ4n/HNZc+0rByMrLdYj8uFw
yZ6/S3IAKAdGFD0funeVY91POLkYHNDwr/OJDdRdIMuWj0Wlo/Yr1TLApRYP4uW/r+8MSBWxNqSz
PlydAupzbqxRUXiInstoihllNUQIpz9j6zpoLwDkYcz9lrFQnYfW+FvkyPbldiQIX3uJaDHMmy7l
UEzdGuscQrlOZBrK8z7HTonqU8yiK6eTyxOk9jlVANaJXo2Rft/PXIA/nQtQIMHQ6R6BLL06dkOf
ChmjXfHQE57ziatgWnvhK2jm/6oH4CjGcmueneX2tHQKjeJCOuNEEw4/wuN5NA+Hxs5uotL92N4t
YjDod5nhl5oe/g6E6PFr3ErpxRtdFtfpMUv6cuQcjPZTdS0QrfCJk060+oorj1Vi+PIUeeSFQHKW
ltCcOKBAKWc92raHdCc5SzC+9LqZL/64dPHhmfFT4/e12/lXn+W2UHUXZVSze8epO1k2vUHwofUr
yJQrxGU13RYwI0mNQQBTh+mr3uK7ThF5lYhmYXpOKu/bMINHgRsbuuL3VFIUUOItKro5I3ywTYR4
Js8NDEsZdyrru+yRnrNc9jC9Q5eelenq66YfFXPvhjtxDBDCh2gBIqZwGHiOthwXngdyvTf7NTyV
mPPUUEbSVtXqodGpikgfEEhNdR7NNqDDx9IH5asFiNpBx9gNADdAmrMFZfmbpMzcY+Wf+steAzAa
lg+YeHK2uyyf+zQhDs1qbZhTfnHzicCSKXnG72vZnJvIxCXD/G/JF5CPlxTY0d8sOBfDcPIWJDFa
stkpvUq9hLY2kmeTkWOz1aP4Fvty4DhNQrn3YRi5zXjP8lqx1GpXExOQDfleYloohkCGokm34deo
+GKeNgXBmM3skErnF1j3l9MWHbCbOwXGd50ZkZt0OGOho50xIj+QFgCEjDzEn+8TWbvSLZcFu1mU
ZL0uib0XC04YO1hlgQngEFkC7tnQj82snyzWpN+bh677wu+/HeSe6i8dr6FL0Zq6BP56BoQY509u
33euxnsfT3JFHi4dicCTVWv5u8y4U9FnK0M+IeiLSES0xuEr/YB4hDKFStDxh9yirVya216b/qlt
kixZOUA+GgtlGTQI3SJZHcztDSDAEYeDgzi9zFY8AZV+Bw877SBq9DPecD3h8SS8/H0tJYWt/5B7
9N3GPKKk/NEpwFb3/MPfeXyN5ES5auMZ8gvT8c0i9DNA5fWl+UopLHOiam9Uek6P3nyXZy0JqeZA
tg/WL7tXGW0j2wUoGMLW13qSYVQMj9SKVKceSbkM3RP7Nwmzn0TF4tcyaMUSSNyBqo/xDI1xNQOI
s1QUVTxtomKnvc4rzxZzrG3VSGlSU0eeDWZ6sArUWvf7A0j0IdfUKiQxkJTc7AUYKtZu8eVFvrDw
ncpARL4txVTJT1/aD9I5QSFPm3aSDp/doXIKZ53lbHhCLyEsIEnsdSqhJpKquIysYj1ZqUiPVpPd
lloo1Rum57yeVFobQAt9TOHiwAe3EAEGdGmPlu56dkNgoG2hu/Imdri/eSUirCXudXohm7PWB7Qp
4C34VRbDRv3T5dK7pFDr2cz+36g6TeUcBku4/yVDxwwCaTwC9z/2MaWxTNznlv+0k4qLKCzInZQ1
tyOOsh0rPxesLbMVoCZpPi/A3gru8CzyhI5+ysavQSeNlUbm8y+GtmqMSLZrT8FL0nTgcp8BWr/9
5Mrhk7PSfi8EaLBBgXcZ/A64uDSKcPx8fo7wARI/z4MeO/Cix4Xj2wnow9mReBG4Q5T9QEgbV01C
kD79mfoaeU3VwKfly07TV9E3gL85E/7U+xelnU1oewkOVJbdOZh9MLaITGHUqE2EZw4czu04MmNE
bSIIA3Ni+SZ1+98cU16WFTqYOtJzoVKTQROGrqN6eT100VSPoeRrMhB6Sg1RGLDNd5kUbBYRJvLf
VL0Yky7E2Ak45GueNDPmNPqP9c+X1H1G8idvd8TiFcgS+DZum/VeuOURO/4Ligp21cdWshbn8IHh
swL0k6DcSH/JcCfhWWEoL312e+EPAZflfWNglvsk5hungUHnodUfnBXqxW/z2n9sIbYtYeSZn1qW
QRBkZROHgr4AZxat2kfimhviY2gwYHa6PYJCsOT4B9Vu4Im+Ddw0u9eAMo1WDAzLzmbmul+6EDUu
7U+37T+VUPzTkjN1maCA8AvRV/H6M5169c/8hfuP8XuuSr1e8ZGNJf6bn9ylVPo7IU6MWw3NKkDa
hqiuCfkZfPt/WA5Tropz0avwuW/y5ytDwiByVw7g1fuxMgFFfPhdEXrfYHdgbYmzsrWXjuQTdn7V
m5JAExBaTajC/frTN4JdppBMCmeI1028V6gpTmDkmg49rFrxQh9schlOkzL8N5gx7CAJt9LSa33t
U/2Yv8HEHbL3xRXVGR/DSe3b2phbSHpaXPti2IR0oCQX4Xg6zAmhVqgDol+S/tdEt0NUhHlvDzD/
QySi1KbqDDZU7C+lCToszbLyhytlQKtLYOZhn5K1ePJQVG2szf5VGKA0aR8Xr4jz2lEJjEEh6M40
Mbc1OSHc59MYPwqrb1fCxONPmQrQtLGRV1Xd3oaxSNVnZ+M1RnaTDyzB1VRjS5K/MasowPvbU66D
R/IMZO+p/wk1hIyEKG3qQY6zBE8RYJrjTus7wtElMJjYTYGqbL102qLWm6L9Bus2OvCJwafFNAUI
OpMBb3T/9L+rWIo6K/BB9XQPUYxBFncIdlFf5sazx0xv3YXM07udqaduWw4NcM6ztJkmUMHrYSI/
YMoxT76tfdFIGAzfdEXR0EW/ugeSjlMVnjJ4q7qsGGzPzQWn8tLuFrnMqK+qF3UJlXe9fOq/ywip
Fmkhv+5NN4psBq+T49jmmeQNHxJ/klpaQgaK5l2hXCBk/bXTDFSROUHo1U6pcEX39bqmWjmtj5Ec
fkbAvWu7v7oxdIWZxZy8PGHDXUdjrOYzHV4/s99XVDvjFmzYLAzz17OseJFwt+68xVv8Me8fhtZ9
VPR6VjIVyulIxaZMBBS0eTlp4ay+HJgGIoGJ+JuPT4FByrOhBLtDH8uaQk5YMGu++X0HxthZb74g
zVqkrwR49tsysOSrZuYBE9rKZGh9bHSqEf4mHwJcXiTPOVwcPVP0FKYLeNFEx8c6ustExEvfgJ5G
8NPto5fOWQMfNp9vwL/8lHNo4rnYtD7kVCUK0gcu56ho6wERzq1LDszlQ8omG0lt4Auk+ijf4mfC
2lNLDS4q+ZnpVmiaBPWrS9qMtybybLxokquLkSReFEtCQDdGqy9WIeY8YOxzp48syjtxC6AtQRHH
n2gWtUHlhFDvgZtHj6uXXF2DT073z33oRELd8adf7c9+sNcaIHmVlK0jaOQszPoWOsZJpkFSiZtp
Yma5iaJdXhBectKyquoimxJ9Jkef8zEuAGuOEpveh55fZTVLVElDhI5Ge8FRwAmQA7oKZQa94vQ1
ZzenEKdUAOcINx3cb/cKKocJJWerDoqKBfC77iHL3iHEPc/+gCl80sduEo7OFjsJGYHiPwLCBwaT
6H6zSHioWFr34TV+fOmHQJ1Fxrn2vhRM7XCobraF0d5/MH0oNpZuthQ1dCFrglsnKeNPvMfVlxD4
JKibHJXeeXK35WyIUPg4kM6XL7T5dOfdfC9h2rY0PLyoNUxFcSKKcGT4vEkqkkGY3ukxuhlHnW9u
6ICYSS+Sg4csKu3Ad01L1JXUa3tyDyS7cmB35+vZfxix7XvooehsZzzUOEXU+mB5oQerz2/akT5S
ilHyKPxTl6fiUT2uhB11tgyH9GQ8+gZljDw9qgpguJxBIBxx2FeiO+hX8YPz5PfrSAPl9J6H4ZiF
M74wR3jUiq/ADDChMJGTBd39hkPq6CZQHWMfSEyWGuqigfNZJ1+aPkp+JTh/GO5yUcpFrR6c58yo
e7U6vsEd7r8MT8GM2oUlDgLOz/uCzRaFLNyoFt/jai3sR67VV78BWa6AtdbvaWa8nS1BqnYFhIym
TtojnvzwEfLRXmyqeIvD7N0k85TRjEHCEYJHeNOUaP/7qB3uS9wLnEMDffsinpO4LSQi+/hsLPTN
JWNOW/QxMU6Vp2UjAuQG0BzQi+udH4AND42HEnC9bkvqMz9FKa2gbsOCvXu7DPcE46/qMvZZ8TBh
a3yNA8YcBtUHfP6R8PpuX4USWkJtmzSNVk0mQleOHBCguzrS7S7D+n4IXq1x7E+YHep/lO1NEADw
VA45sdkapJo9bN3UGqIY9o/e6DNM61MRAFKcNtFb1lUPbtr+WU31UnjmNgOgu0IVqbZSoslaTIsj
KEGogD3Oo+Wbwe+sbXjelK2rMXrjo/ekWpQ7gnSOcT6DcedwRlSRsAI6ZsxVsycWSuvRMfcUkAym
RDibsntkpYbQBc2hYpa9C9iNL06XzWIVrMsZZr98iU2vt7qfNEVHFSyzP60IfkY3Ntd3T3ymYHUF
FXw7xoWBqs5LILvBRhHy5twtWKgpBXQG4+jw2HCk03EzTKhk0q9DNMVErpxHEwV+zDWwCbCwZn0k
HEQWtOVpa9XldyeBtmjOZbo3u1lucFEnfxFwupPqf0SZctevXgrD8Q8Izp/jTkqdILW9n53RJh9s
RbKaz/U1szr+3GUtc06JS2C+IHFope+M+VTBmfjUok9wC7tGthv8lzzK40/FzDXgnzwFZ1SRbZor
rmaQsUQx5w4qLBRpttBcFLstmTfP9BZlryPE7WZ89YDa9UMCQkGeoj7gqnKn/q4b5ob45O/40uVu
UfKG6FKUsy7yfw1YnXgzXQ7/hxGUynfP/aeQLc162BofiLF2vQLu4cAXFw4WMA8UEQLVVBmhQJ35
wlIq5CXrKIvwuhTtkdXW3ySiwQc+IkxEgk7mAhxp1l27Y342lmyawPcHkp7vVyORr/zHzTR6KBCb
H7chNaGtrJtRLR9bCrJkhbl9e6OgHEZzjPtdYijqTh/O+IG2E0kt/UoHmvVpw3JGfi9blRfgDDme
jC5xrkHAJCHKcFHDJ/Rr3RngN7wNK1Eh2nuiAzxXYFuUoC2zHS9hU+++oBLwKaBjIKEwNLMDueBE
sbHum66Zms51EIwPytqwn/lUp9ltHg2UyLLeY0Q6u6C2nKQg2rDR9nMafW71GqaI24/8v+vixtDw
9Ej8sdd+ogU1H+9CEEOsKvgy3veiFwLjBhxY2mzklDlU5bXQc555E5ryLHwkdLb9HfzvjhCC5tnx
WYof4WQAx27sXKsL26tgpKePG0/kCd2VtD8EGieu8WIlPIzR9jo/lfvZSBb0G2G9MQZ8yVwoA/p3
25WeE6Bav+6iBSwTO5zFDOZYlxEgtXiIE5RMYNpCKmfpqtEf8mxtT8ozbCdYHXiCnGw/6+SZKka8
U243bvNmfdPYEKj3fb32pEWfrTLUY4xgQEvFOIPQhVjSJn4WcyNzk3nh9yTt3heUUw38sIbO/v11
elvqX/LYLuZtks4rRz85bSpSXC27HRdx4jjZh/Hc6Kn0uWe2oyZ12emqQQqa5FVczMC9XAY4KTea
wLe1EKR+3YD9jtSGL2f2SRFTzViWkSB4G+znAtk6Gg2qlp50cHZdnxvmNYhCL0czhsHal88uoFBr
BJrIe8B8evP0xkMCqytcUQTTn8TW7fThxbNbcGeVfY9bjgtv7ONfgLATh8WbNqbenID61sL+FNV9
tDA3xfsaQNPUyEVi6A1Sq7vj21qBFzUUmf/M9jY/VjpQ34MiWhDqgGjj90XlG0TkLFw2ALNqtirq
vKDbmN/qVepDTB4Ug/ZFZN9OfZBFZzway4wMW8DENxt6zwnWhTus5T35lOqDOcMKAvTVTZCFZkcq
MB5hodrDpQehk4zR+/QIfJGK7jKqL5RV1Fn2tvph+gKVCGDfQJEA+91VOPx236EEamIsSyA8EJ8Q
gxOKnVwhu1ETEvgXQpTKVIcVwWosl5Blvi7xXikCnpR4SNc3NyiamgYR9IHG8Xlc3gOoRnNkYOp6
33enGvpGzc137xH4kdx7ZPxR9Xqmr6vovtgJgGZqvEmrsL6HH/IbVMOkO6Qp1NyK947PnUCMhQUG
347FA/4xN05ak2coqbtyjOf77I8RfS6RjpD/HQIejjDJOlAAEEaflbwZ6WTPvG/1LUbjNMQX0nUJ
9QR/xWTP0v/XM7ZXZpn6zcGkNEoIoP4BxxAbif3LoRPac0dnFBS2/6NJvTmOcu8ang89ZsrLZk3T
GAt5kbDid2fdfmODw75ALdVlcl4+mF1qfcTqvqbUlUQRkYOzMblz8BcYiZxZ7JcATDanRWUUqe5Q
pN0BhZbrNHPaU7tc58mYB+crE+tEzBhq/RcqbTKhLInjEt5tZB2uNh4ADERuckoA+0gNjXERcKGQ
eTbGALhX6aMtUH+ott9f4NAsBa7+fgkn4Y4F95lPTwK7+zL82zBcxvI8COptOmSjdIPmQygD60WK
Kp04+TwDVAbHsTQDKLVBFPlga8yXAOxxR2N6aE/tXNAPX2LZ205W2ShJy+FSbNE5KNVgr8lPabJO
HZ2D/cfhNpcD7jNH1dmvAlvTqE7SYYQuq1XC+0XOmKfRSqoE/gOiacfUctcu0oYq1KgrQknPxgxM
RuOoGJ4WILWeGqiR0p5lBj4r51V7hv1pCHamWVixCWof8tGdNZbVzPTEmp1fb3oqF81ynbF4834i
QHoKMLjBdGYZxgoz7UZyRxg1N0DpxatqloEFIMwSVQJlYJcML7MftvMnW8Okz1iFfAl5ygVflcqC
/nrQozDMcHk9DVT7o+A9n34heqdKWRWwqzTHMtgNv9pdj7fIykDXZroB1SR5b1qWB65PEfZSmd4q
DQ4DSQYiGzPJhFS1GV1nEepFS9vjZqywsTRCIT5x32n6r0vMfQ9S0JRrwHFtu46N+lJmo8OQj+MD
o0JzE9CYltt8yUhAwnvBp1vmhJ2dHiJXxuUsMZVdTLcG+rSCkKLcPVkpVfqB9xoVWc81th3IHO/7
BxqWldpI0+s2Jqyalvpvcn8EEkncsZ9G2Zn3pK3F+WZAfuk2a8wMw5wQvO8SDaYh/LOS+DKmeMTT
hnFIlbFsu1plmGtYlCsv9G3Yq3DZxv/MAdBs1JKQjdGkdsjgFmHa9i3uNF/31gmID7VN+VRZqWzE
oEtQWlD3XTt8TaX3VyZmTGmV0DUCjUf/ExfO26Hxxkc3SUk6FX+94xoS7nvKhK6uGpv5I8I8BpBW
4ov9iPUmoXSRtNJYMyXAkm9NN6WP2MUdwPXUiLb0N5k7SgufPfiWCTpz2u5TSl1bSAE46eKQq4xW
e1ieGpB5BTe5vHfcnnZ8OoUrI+NDJ905u4WZilqfq+ls9SHNRnUpDgXLsvKIAhgW6jgJ38FjFSu3
OrMrsno5oXY5YUQ3F9I6U1dprCZkZE9ohdOdFAMPR76pb3hIuuI/WlK6j64+4SMitaIUBj6cuWh5
1+KdBbRQrWRkmJTxWrwoDOb1GV1xP5yvJqbC1GmpVOFqmBIIZdvPJ9Kdda9rJveG2fGVjFOt2xXe
iVNn8CYf6wkd5szDgZ6l45g9J28q7nu5II0pDUriSe6vh+M6S0QRbC36R8htqKP0wmUp0cAWa2nn
r+ipum+SWIjm59WyFRbIOEzHXv+H6YeqmrlTbQd8Oj/RWU8bDnzYA7o6y7SWhEo/PdxsHpXJPCLi
QVUJV0QE2Vmvv/jk5b31nI8H5k6gMiCEK9I8tukmVLxaLvHkiwq6tsz/CNKyw8Wrg7Ni6jusSqwl
NOHY51Y9sk+Ctz6h4v06JBF/Ib76A9xstJVrmhxTlOx8ZN5q3nQYBhacsVgg4G5YHzWUs5JrVJNl
3h5npDCCzlOI9ZAByzYSjVirYymJZFexSgiuyWV6Bhph186MnrMCGF6+dUaDS8yGekpJNKxcOiC9
BS4fnHQsh4iv0TbkaAetcWHxZAnDbwDu5AV85JuMpCF9TB/zb0TbmLi8QOfIPqXNq690jOP7Wpio
LseDUewc2SsEPyUh7U9KmzHqvf2iAcPxIQxbWkGcIkAlqLl3sgG+Ht2XgFiWs/1fcQ1SBUGmKExJ
Nqahd+HhkkD4fk+jkFWx9W/M2fl8l6hdDBAaLjGAo8haMWdoDrbGXf2cxPKV/oVH2TQlyUP3qLe2
Khi0G6XJz6GUOEi0ekHJqo+rCUzwicBeyWzVtGX+jYvYfitRCisw4F2aveIcfIKC+0bYxtmsegEm
t5BikWZFj4UqB3hTXSW0X/j+J/sW0S+yuqljIdRRI+IsafvkDj2xd5d1qmKGsFU3pQ1uxAD7REjF
MjnNry+p7MXVNGlWJP8UJ8BQgtPy3y6RlTCNGXLZYXsUMoGPFsws+S1mF/CoLK7OywNJeH53AM1y
gkF/FQtLAllo+UEuiFVuSlfFfa+mzGVGVSIXm3nLhHnEgBsWhw6uksXXp6ihhBf5C6xGkAiNN7nH
7CrnZ0ZKYqRHpf1cxviDRh6tCNmXsWaWqFOLN3vTfHoHpzNSVcK435b8jiyxrxvlV1XESeg6tu4n
8H/C4w2dkoWxUmPIJgWPPUEzon45md5BHuJ4uH2VXTnUHoAF0j895WhXTyKVlnzAHFFsu35OjLZN
jIWrqwDGrox8d9j7Z2cmDZljt6rRTPe14ithqQEx4r++JMILydQg3Uk02hQtWFDFjqWTQE1tkiql
vLmgFneN3tJtCMkSD2sQvZv6XBk1AoXRWSQnjOB1UxfLycWhpjxiZ6OBm2foY7T5+hajfurtmsq1
h2+rwKI5C+/ppu94A/7/qQLIG3Lp0c2HwLdiKq8HCl8zQM543IsVfp7KQTfP8UuGWM1T52zVqcH5
fjDg9SAAzLx5cmi/8r1ts9EA9UzGQz0ZhCm9GXXtu0ElfDvpsvozfXVTR7A3IQT8eYcEw5+RTpsv
6KeBV3451ljH3PY9JxDzasWwpFQa6zTziNr6dmgQ8Omjt9nQJORmelGe+IJgxUkn1X2yRvsebsg9
naL/OIzCM1uszgu2DZh3qEl+5hd6CVlKbNdHIHPmD+kVtkSRAw/0etqdDBhaGugsrZnaFZwUb8hV
Det7kZnoNk+HlWgXU223AmY+EflOqZwBG4L4DtoMOq1/oPcqE+Rc907DO/dpncrmyXCAYsE2Gz/w
VcjNUen6IINRzQwtPJSjT04XtRSZFyzX4vi11bDyfYfgnsUeTjg6gN3566CkDZGj64KaAuGI8qcn
OdXR2xGFT94FwIixK0YiqHykS9J1ZiyA7hwO+tE1+pcKQOjXXOJFVdbtd/viffZ1Q2ULlekDcF13
u5n2os/V5/wVyIF4vc9G4nAG5ZfAoGtchGc342IMvRfE0NC3zIlDEzdlzr3y30m/RRZcJLRQ2bGE
pfIoLjh6D6fKbtDNPVlugPgq0NZuyHH0A5M8Ouyb7UfpFtIiwn0SutSFKhCLQAjG8v38esfteHo3
7eueqKrzL+5xykXfSdTe/YIyRwHKfVMchgwuBsz7FEngvHuxAVlzQ6yvvofTZLCfAJEDrhTpk5q2
KOWzumNY7FDTr2FtX/XF4FD7GdbinziiR4BFc6o9bt2nOeM4P1fAAOtDBdNAqOdccqvpIQ54WDXJ
4ArJs74fwy2wTcVO8coxvlSOhXZlxzgRPQkif8AP1eSxCNyIZWPRR0oS4tBysVtjK67py7KOxxcd
Izr/3k0aMKxKCcStt1Sjd7FogkKXn5fpSN/1nDd1zyHsP7q3eFALdvfWnYhJLzU3EervyrUbga1D
XL3CTYxyS/votoNdYOsLA0RdWbenuSUiEEMw4G5TmKoccPDM/SxKk8DOgazwcLz9DgAOmt9LTrQ2
jdNZFfSRWs1Zl5mrWwUxn+IVAnVVd2JbzmlDcpOBqLzbpBtipsCwtCQFJKSsT5z1FdIsI+4wXzYW
UdbRAgUKMt8GyzLXaH8Q4VtonBX03bDuDVSaX+UOhEOCVvR1vf0yMXlTI5+tgB5ShcJHx+aw3su7
CqYXS4/kDAoRaqir+hnmJeJLPCMA3YP4tn1vGuhv+LvDXc0B6c86PYMfgkp8OrFH9B41sgbXlHdH
nlxNxxXzHl2wbmZIXSJbzfjNnhHCUm7T1BI0IAP3FpxsAr1VZlGXftJzZNVwWWj76yuebacPAG2w
ZbCxtmc0/VjwwShTz5UaSXS2x+FAfB0YpKZo8JHGQtvwqYTVH485ypqv5nh7avnFR4nS78ciZ8XQ
Rek20t9G/ILhnfsq5856eNrOaYyffQkUGH6gKrWajLYuiaL25ylJjzuX4jmnu5XFj/3tk7VGGaGr
FEM48GKRpv+IuDddUkgw0VZiXVJyI0yHZPq4kNwUhKfofnnkuEq6b5D+F9voiztj2Ycdc04WcaL1
KbpHXLi9kwLIuJFZF7U84MxpIF7wHBxiRiWK8pgoOi6rsernpI4BQO8cFJHNDnf+WzwBh/047X9x
MXXZuwen72Vqcn2eaP4XSha5SJduNE1ToRTWDVJrZZthHyXNHYSKFGHB92RiMcfUvN9e6DY3i7kg
MrumKCLVjoRdhV/b5eY/vaYZc6Rta4qEzyDdNoyzcqu38q+G2y6Xa4Drcncu/lhJHVF3rGBgYBW/
Kk0brdYqJWD414qehoz4TAl6uUbeolV2bA6ypG4TZmK+cmpHkbV6IxTHPKcjMwerGRkgl3rA1P7c
IDKOYrpR/3iLdm1LEspHuT0CPPSQ6GZTWHBxW2/Sw+9MPIImdxoqkcg5MoQdroqdZNL5T2T3IpLU
DL9fmAaBg2b8o5mSxPrcuqWbIzYEBwhBOp0x9FxxcEFKMHq59arlRyW8EYYb5UhgU+0k0djkEFAv
02kNEWnpb1f1mVTjjA2MD/sGwqaLRlUc6/lwUv4BCL+WGLrwQK60Lqe96QSlWdq2r10r1yGA4ouO
lvFTsBB7ylsx2aU4HX5XNYnx4PmXPipgx62WeoUQ44cJgffKOASiH2L3WRfJb89xOHsgBRX4I/P0
Z+SsDDgaUbTf+YNdDTXJNc4YVlQ65rOnTivCBSFIPnw7hU+oYyY9xXovQxFLDfjt1kHnIZFldtTa
5U/WxX4vf2syaKBICPwlCNb8zIiWXXEe+qOUmT+MczwepCt9jVwHPTINZShaTJKyi/pQzWfPfQ6H
5dQwrkcpeMD5ubkXFoX4W8EvDdrQWW67A00DBnsYdUuUzLsottk/i9Xjiu4f19qw9KweWu1Na0Eg
n6KJihDbOcO8CKSWOIm2Ez95syoo7ejMNwrxae+9qVA29mMWKXlM90BOp7SKFIIjOaOOFGqg0W8n
QebrvQl/GFLIv9GpM7Q4OwxskINayvrm5P+jAebhs5LPksUon+uxTGH847aBbBd1YCqYO0WR0dt0
9aDbabjiKMoqn5mhSEM90WS8SGQqGOA6/IIuT6RNgOL2CU+TYKnc6GG/4rlNXr5EAOnh0PzLPRCT
Iv7DoWnDEe0GE8z7LdIF8WCekZt0MyifaWqi/ElWiHY1Mue7O+grZO7wjDlKcIyx1esUmFMwjMqL
9rJLu7PYMkrSFrFkOluxacL/URKNTsU1XupdE6iM7xnJLdPmS/W4zTPwwlbB4VXF/PaL+eTGKl98
daUoywNRy9oPQfCuHzsFBP9Q6zPGX2a4cjrxJYaiXZO7ekBSKnR/nmbcGrgH1CDgcdyFZIAou4SR
rzvKxi85z2UWTpaYMAbAcrxKny1K/Mi7+M98VNzaicK3DNdK5RHKGxk/qPeZph0IV0vdRR8z1MJU
oN3nOcEwQP0xclc9AD4AcU4Bxmhc/ODwhPvZtjsw0FeOkzoFAVDHzfOXJuqaapnm9bH6mbH8eOnn
Db4R0Jc3GwVxlwYycFnDwz/KQwaYbBCwc3Sx0B04M1hbee+2Q7pXndPOkaV/A2JCYQCsWtyeZQ6T
jP2Vgu6FrADGQU7kPnkeAPj20eiOO2XGRZdBOCmwlAhraWAvoPvCVbmpr1vuy3eMxF+9wsQKEeoL
kQ4CTonUIZm1VhBb6RizEZ6C6e0mD8mSPJmKFv5mAkp2mCFpbV1xKMY8QqyL19v4kq6wVWQ/2zHW
rSrlW6Flv8aeJO5BhsqbcbdC0A8Obkb1DThG2Akaye4rNAtQexXoMZau5iSWoQ5mmy5Zfym+HDJ3
ZjcAAq9lrFsdMOpSh2WjlQYn6Mq5xIjsXUK7YRZLKH0Sialq1dDXZP3iuWAQQdaM583e/3hyDxSf
0zjMk7pjJ8zeRFHMx+PBPdoybJIScvsjhh8FbwgYW21rRarX9pQc9RbdH70Nzjpzp6hp8ziz1Jtu
XzyQ3hmedQW46KW8xk/JVFBIFv+adyYwy8SpezQtmUdtBLWuFL8l1BCiouSPEk0+xWAzxr9q3aIZ
OVnwxn0BZ84u1olkIPEbzUK0yKT04R08BtCv53XJlLW/W7mQg84dCD7Hwg+sLnn2kDVoqxJRtgSt
Rp1J0gmh7iI41A3Vlz9ofi5tuHdnEzr4Mt7rCLnJYmAS1mQww6dFz/+nZfyRHSDHUohfGKiFzqzt
OO+d9KzRnRrMoa4Uw0ON4IRx1t2KFtE0qIon8/Y1+gvqZIpXfMxolrMzrVfetji4+empFTCsL3xb
CrR6xTu6B03bEZYudxairLnkj4w6zYdgLAKBNeyHz8WyzPOmKxSdsP+Hz5YtZga++XPUEOxH6cYz
pjjc3j/Fm3NmgJyVmRG12dTpzDCF0ZEETtGOIHErpKowpRoihe+bz0suCpCL1Z3/IiX7xOcVOXwX
4OEB2cmAsq2muFa4FDskmADawScQJVRK4tkEYV4R+R1BZy7PZvw3x6eYCsao4KBHREwYmi/P3Ge7
UCmB7mK/JznuX6UIG4HRag0VPASt16BrsSD3E3KdRG5WUnfwGIxRfh9qPS8FwQlxqGB/+kzX1tD1
s5ew1NoYPYdEQe7/3hBjnFMeRmJOpxHp9ftm6NJXGbmupmd+FjMThB075jhjKRXcgMP6icsUZ6fg
bIMh0lYzVNID9rnEc93ksHNOp0cwWi6IBK6sPpQfYL1n0mEZydZoR0Hp+HOpepnN5y10FYZc0/K6
1dRYOg3JG34wAqwlnd//hLOKkfhuXr8SXdrfR4124s7PxvWCoUsbDoH1nnty9eZttyYgE376FBB6
McnUkCXtzT57z4PizjlXeEYbRVgwhn0XDztkXW9GnmPjD2jofYyWMKKVH4Mwz8zXblOC07p36KIR
5ItOheIzXeC877xyJ/TT7CLdL9sVp7JEKdoPNB5Zueet94+dNutjgSp2fJo0ZOnyXVcscg4aHl+2
QAf7ZzL8dc2X+5lldUDtpifNP0fEx/o0+2A0L8y/91VBQ2UHZdUmtPTSvtALAogVUJixiEsFoLCH
tdx6CCP/s/4nVtb/plOMWx8+NELSHn0TmLIFM9QbL6K3UlvReSsbDj0w4TYK0/j0w8vRe6k+yhwT
SBx976vZrofaRJ23KvzrTNyNdmo3Eh8gzqqyP1CM2fdeD66ETNK4B02NvLEbJ6teW19tdvyhxp9P
44+Qm9E6TxVZYGYCbDoD882S4+UE2PHdkiPinFEKz6YqbEUZxP+0CTlnIuWcohZMlEmTyPDTiu0p
WP2tguUreWfRGgJFvEtooPixwxuNrI2E6PgLrJtSFZRl/z0L9LRpTTazmwEHn7KCbz5vBUAS0CyW
GdjcePjqAAq3dBZ1Jka+GmOV0R3J7W22UAzAqfk3STIBmSI1MZXxEJ8nw2lUCd39W5zQU5JbmkgV
ebC6u/QW7iy+Z7WByIfyXZb7Nx5daHizug6teJxnrHZJHJxzjbTG5PCjvLCIU7NMNRlqSoThL8iB
oA/tgZyvh/7JZOwkvpztyZkLrvdL7wW/xdntE9lsSadbrOWDBES1Sly3jZi2D5vNrHI7c0SCOwu4
gzHiFsooXJUPUBHKqtPygZwhCCqVHwTnx24WOxlU5hR3QyJrRcO2nIlBsHo4YMcok5DaB8R+I2vw
ifU4DkP89wsHfWnZb4PNQO3EpG9+8OLK+QDM9EBHwKoE9J2jt0prgQxjF58Vczy+whieOuv1jJHh
XoJcRLp4R60ysAyaJi0njylAq6PZaNcsxAn4GAZcrhq4hEoKE1OzbPCIcrrHQ25IYP8Wvh/FGmts
dp6IvBmh4LBrhyEMb1M6IoduhnWkvl31un9Yrb3X0lOAlPZfNsqejPjb/JeWGAjyOOWV+Kb94rmC
ejsFl53A40NnOtHtYVqEajbRQi9fi+LkumsBryu9QPhzhPj33rNl3SSJz305UQl/uQOmPCQUBrFu
03tYorVGUlJPOVDGmOyDySZigdqqJ+8KTbJ2ejpkIFo5/bPwWMKS5gIbdFG/IKLa92ZCv1imUlmx
zZZ6GZpjUHxjK5YuAz+zJGYL9lH1u6b3XffLgQ/a4hvo0rT23wGP5o9qvb/IUur9TsC8U1n7FQb0
qZsG92KrazI4kIyVcvDU0MU18rJv/rgGrmfzl6f5By63UWyJyfE0M1GNQYfhG8M9Ih6DONaxpmAu
+1Zwsk7H/Yu4CN74Jr1F5dj00ncWWip2V3y9CMp+vLCpij7/UZ3Bu/HujTONp2w0lrbmvf/rfxWS
wLGIqZfiJdhyDSP/fGgJzK+FUxrU6bCvxxXifh8Vcw1r8A67LOFQwLbmfi/ShGGlyVoQR68BwpyC
UCnrZwzwNO2MOMEruL0utujAx3eWA0xgi5Pu+Tu7+Ahf1+GUT+W8fSFGh5Z7Pw+aB+YpvROfZYDy
ZG492QzMDxckAwRim0RKxlCQWvoeL9cMeabKQtSWO6TdN/on57x2ppi2BiwujSJ0wRgMGgQgI5Ug
lc2kq5WoWUjrtVwbZL+k6i/1Yv9cDUvMbp5+42mURplbvQVSuG/IRoqjgCw0/mdRM7eaSjM5fhAG
wUF69JLZtjt0NIxRSjHUdWs8jCJPZ7hXRdmp9zscq8APlQLkLeoILIl6RfD9nWxbgt8Vzdt8a6FO
BBzrVSW3OO9wmedXysCaLs4PPCy30FpRqiyPuO6nduSUNGeyvn2YA26uNqByQC3HsVHi262R5VSm
Gr46Mls13owx4eZ65ZkiNLC9cdfLjRkjRzVtR5QMtHLL+bX9b4p+pHv7qnhMyG/OvBxuu+nzn7Mb
l3oqCNSviY6v/JjB3LBSEE5ZxbuhlVLJt5igkcMdgMdZBwgWe6w2xJSIw+GgKhYrI23/ImjvpT5V
+TLM4zclbS3jO4pdhBMAYHrs9PEdGV0o0FUgQg8+hJtWt6vRvikql0tGAxtMr+a7y4tnwB9iaxAC
oBCVE+zXMMI2E/ogBcq1mK8nML2zdX77ms2oWOya+xpWdpBBoCMHyciEKT5t8vZyGoPGHXAzggSV
tTmXe5RXu50Fd24qwyEaggS/v84KqOI1uJ9WWj6/T4QclSh4U9EpEGn4V47gBeO5Lp5xtJ7QbBAR
z5CJ68J8/xIVoyTLcP66mIkoRkTtxr/5Uh0eN6e0VTAb+5+Q6489nOUODLagSbOnVf3nxLcb4nX2
YHYti1DubEqDYMOf4OzXRxiEHmowF0BqjZD3Bo95+Te4ypfxAWLx+x+6dWn5EwQUy/5HWgZG0iIj
tVMUisr9EH9NIEsUZIHAysPvlLv1dRXSIU7SAsPAII3X9Kn5/1MI/iYZmRd8EPjxb5GPFvpfNDRW
RC3LwBHdr4cUT0A94LpmnKCw9dL3++gYSQpmZKKnEYcNPhFHHrci5gKv1/17FfwAYzThkqHBg7lL
FbFE+0J12kOOPYP2S2VRppEtjjBpHgeYEuoQK74sinaPjOxnJf2yQJxjNnK6SkCmMiF/F0Lw2hf2
Q2nosi5yAcjq5EfHm9CLFCIRDlZi03qOpULnOTcXiXg/mM5OEv7t7vWrYyDsHEPkAMD46HgQV8Nd
soaUKuwZrIck7ztplRe+8FgwPLIRFJhcgVWWeAwAHrKdxW8z5maV/PUuUU9qaYI+0MJJOVeRTjth
Dw/n7rrVjiagZVeCy9BDX5DiN0rziFZV8mb5t0JvzGgr12fMhObz9OE4L0qEVZ///ayQamJmKwd6
vpjIYDc8pKaOCg7A9YjwzQP87qcfBxeP2iP120iALj+1OU0KODethGhtY3dtIBq95CCAg19GI48S
mScHwxM08IRrnPT7zcZqmksRTyEVruXjj0CXG3rUkJ8VCR/aIS1SPhnpMoOr/oyFjpFb3zrDHrac
FFfL2b9V3J/H2RKCDYU/kpXQd5xTyulQrlyoz2sBV4STQJdzGn93kD4PKM5EUQ5UWIyg99AFKk1r
jVgBNBYU24SSw8fZXpqdYw361c8r7NMev3E4M2MfSDoeZecdIODhcGcsVB67YC+21PneeeFzkfDr
O4ZKZ4XGalIKseyju/2msHys7UTwU4O24aLVwyLupMYiztnviBp1OKYx5+J9b0RURYcj3Iz12z92
wThHePNwf/Pe8OsN63R1ZI2SN3/KVp1N+Znq4JlpAjV8nJJ1Z9TsiZf10jFIuIhf+1npnn6otAYw
lHIRjl+lIQkqkZrMh9a9/tSkk3RNzqEvzrHZV9tPQR1Sv9hEjZ8nm3EqIrDKcoLTsMORVNEriuUv
5gmodHEcLA10zTIbKdCrkFZDCyYbzspW8ramD0uhJKxtIyy7F9YaBp+gL0cGsWnHSvKPDSDKG7hT
+tMEEWAbLRa36TAnH9m23BYmON2y71VuFkMCAe2qBOygiGbIrWycGLkTRHuCFgLlblxCw4lmP8sG
XiPec/tgguWSm2L8qqXENyNUBJ5XWgpCUkQvMsmd2GvlUe4PUtzLYjpehGzLE6kAY2gQwiziTEQz
qwJRKCBSg6ObzIxnw4agrfBkK/+YHG9pcEulWsUD8NgHBJ65aLW6ZKdXDuT24SR31ZrXOqN97jio
Vkk6fGBapFrjCbf0OdsXDPYV7zFLdtdXRckOaMHulVgRCO8AdAgqe7fTzyJg6lxQ183/K+g3qp/C
1EswDNWGBM4QLkvXhdAT6KB8kLmKuhpgDazZUgo6e3MxvFOqsmos3kOZA0ozbnhsjWTXyLVcsahX
yjzjluuI8CQdwvf0fpooWC6IdmDqLZ9nPAmgKU0+iz97ulJ2CLaiCXFXEqZNjrZnP9CpotMi8Mae
Yms6EPZmaWKQjaJePMFvTmxmsa+3QOgZETP9HyiLeUpWbn7WrWzi4P4JbAVBidDTHgM18ILn3QLO
QBVTB8ULG959KdczrD7YG6ri12BaTcjQYuWJot2ISvkoY7u6nAIqXYZiN6YqE7L4vX+UlRYjfb3V
lbAFMk+85SGfP1ldS3VxRFxbeswxsIiDVSsdytJyCJkX2FXQPcyLUY4igiWU/+r/SpKNQ9KUT0Xm
X6vUbloAfaF4Ls1n68lS5RLRc3G0P1fdPhbrUZ03nI9YcoPjMdDmbGE05CwWD0GzUDYf3dFRIdgn
ZFY/TJlS3X62LJj0c57TTVVv5IgXQCNyunMCCjtiRhrSoPXySzQZYUB3ilC4/MBSzKsDtdT4BEKE
bdf8nupSBUPj6S9hlqixLyGKVdMuhXZpD5OJeJzF/zzOii19cMtc2C58N2jibJ7sNNej8LFKxMc6
3ZXIND+MAehSAqg9ezSPnf3C+T0e5JM4eeZQG+EaJyr+VdxRwIa0YHBhV9DNefxY2NnM7bvOmtjt
iHxhouq+OUWVAdmSjFMcsDIgmOCl64yRBNHGjmDsq+1FyeBRi6QHTj69FUu9x46ohYia7DFR/Pv0
2S6wFCc99z/DsL2+lXlfYFNBWpA9T6eWC8Z23/JMmTMrhAKxF7fX7eQ6lWCIVuys8Bnz/kluFQq9
S8EhFrbtPMGaLTPs5Sn3CukDE1rkzTI9sIMREBFF/UKpbE3BUyz2VaTm0QqoQXd0xuCsxB2JtwTB
MqO1wmC14I68HiUFMJXpo7xp+4BoVuAxQOlLeG5vxbu0eU+r6YruQjKuXr4Nd0LLq2veICfrlrAe
TpIUHMB4J+dihsSCql6Ce3iFP8aCCr8cvVaRUlnlIkNip7Lf/TllWtFRlpJhNlvTRduJg7NpZzp3
lraQCNX+jIAPaeT5F5OPwUlYjA7zkXFgwwFKYXIIHF3JtXaiRfHZwpkXj8dXqj9bMAfyl6DVU6Bc
lVQVIQKlRB0PyV9WMSQiBGq77zbUCVa4xc9l346xm/RufFXACDyjVYOekbAFI0qbNyHhWJJyWhPz
M0t2VXDXwQdFLbAsAFT4x7UMrzD++j9pnmQOx9Gq/aZv4JsGJvA4lTqQqY2R7kT+NvMCz9AfjQ3C
bNNOwnKOsdU5FujCgJlcVVbkUKg64RFEH6cW27HMnTumLI8gysspxmKNYG25eRaMILF9g5vi39MC
RkhMf5Dvlc94ev7E23BSoXfjs20lYRAOpiJRNKYeXxgzvfxpp7nb0NsvouyjQIqVb5Eo/vZa4L1Q
j3LYk5Mz384Zs6ecQ3lJOlkDDV0o1rFK6S1H2cOQAmZTFEYWZq9vhsIQPkgg2Wm/zzDCeIlWkZq2
CQCfGnaTYfwn4LYDfByQWJcixTG6E81m2VXlUIsaF/zmVPn15Z2CAbugA6vcuXjr55hxhJloaTPM
fOwJx35nGp8tAvLSdSPo2NPVeyMQn30oCPnPB9C+5WhytkpzgNwNSf/fxx9r5aIHyMfft1Z0oGbq
Chktx5zdD/tR5Vo9DceL0iXpwD3T/Ey7K50SApbFd/2f19mfOyuQzp/KbL2k4nqpxztbBKM0VH40
tD5hfrimECgh7aj04WSreFK7pu95OFUUdL+2Uvl+jXKLiu5kxF0uEABmEoUxQEkg5J2pI7OZxZnU
COhhngAJhFPWS3tIC98eczSrL37Qcb1ZXbJTaHLUidGzHkvYNmu5QKTx2q3Zo2kcVBao2QJZialL
H35Gk76zmZrJ0wXrco83NSbyUP0WU3PVdCqN3CsAYpi9LvKcHBCfueNNsBWda7wLAv97w7AtzwZn
Sjo6fecGu2+XCM0fTzbJy+MwZ6xih58vz5wHePrMHiPV1Ch2FsfaKG/64T0WXU1RjDr1IhWRmcwY
cdkwvbfu1/xDkPA/ipHttjENuk4xjvD5WxpLd91j26mJNlLI7gy/qei0QUO+lMLB13WyCL/LWOJW
sxqsXVp6QI1er+/2hzUH15xYVyWMKpSa1iQSu1EWWkX8S6fxcJOP77QZya9ozg+WgXZPsxp9uloR
rMKKhSL6mONPV8TGYrrI82uI4xnoeukl0mvRnI/ALhFwrTRrVQKB2RzVkfsRGlLUipc7U7eukM+F
hB8lWG1Vv1JN8waeeFcIBp41r5e8h11weZNNMyzhh2M85xvyOa7vbrAvd7rPWhyPFk7JbkK3iku/
m2ydHvNsfLrFJiua0lhjM08XE6eMdm3vXs5jRW3GXYk7j9mHBvn6PAHz/uEip24/POwTxbo8G01m
6J75VRtNyBBi2FlRCK3pAR+FWwV4M/B1RoUCNUvuJjJAp4ImzzkDqsCDsc49SqJ6HkAoDEa1IJQS
4GlNmS//r4paw6e3OOca+ZL/Ncq3V/6vs8qog41337MFoXQsgUMlieHzvCTpxp+K2UjZTJSac4fK
j1xEHo1BBoKhxJrBnQcjGSBHmOuGEfqJSMf7RfyY55TCQIeupr9snAlfjwCASS7Eg2NNissgje4+
MXgMH1liyYCgO9dkyLVfPIrFcodypO4560keCfjVj0+7ATFl2s0+jLzgrC7iAYBStB0xUBzZCu1a
ucXRGY6qblObe79P1rv20VVFq/c/VcIcr5QRE2WNKeMJd9UPI121N1jHp7mlmXG8sMB0OnvjAFfR
kf5D3NMsJ3kC/OwiyQbxCdHcpuRJkIF/JvQgZk/JJ/XyZX/Q2XGF9U/he5m8wt4zpIkDE6ZJiiFv
o4bVpSq2P4OxrhLGR9tizeSzw9DIJQ6Y3nbQxiOd46V1qrwewsFE6mjd0teDDjh2vuV6p6et5WNN
7X6S7ZaCUFGfgYZERfPdPczQrOTKhNLIqo8ojTbjx5/UX6UFr0Si1o/qLZgnWKLynYCGPLrsJPhZ
Fxfb5Rdfx/LAYc2sOKiVTxHmu5qRTALyWfsVvkger3nFHDyaURLDrRxuygYw3lH1L0NmquO7Ijbu
19ChAVhk0PQClKeYK3yR7D0clGwD7s1p1uYhrQY9xDcQnAOSrBtSgz73K63WzHNaJTyR4MITxY1v
X93z/Hk6onZ6kpvk8qmP5BnPckNs4003krVKPZ5fDmLmQoKk9l7wXAaKd489YfatLev08QJGo8eN
F9Fxp1Re6Skf81fnv2ERoI91rSblsFwOqMf2Xm+xys5PIhF9oeILeAKAqrpP26HBDCCzO4pFE8kl
LFQAvVWO2bduv4Hc2ypz78S7rGL4LBglDljl/V7NcZUkJIG0k6fdmeAXQHW4MzHFzNBdgoFGPLFd
Slq4FvMJO3qnB6CdNZWc29N76tQER0CeZpLr+9rrdj5yzffacgH8TuKPBL0DwvNxsuM78njJlxGB
AiFOm3x+oGqy7lhhJwzbU2h67b7aCI4LV2YwKOi+HTBMc21esXzvenBx3qnJO79fmY2zH/6TH2cs
buXZ9CXqjsx4Ep4wDasCzRiUfIevDa4jK05uPRjeXe/hczBYv0+sF9eZ6l66aIpin2y36wl+zN/u
M5A+7Ws9F21nY/bEZMQG3GoY2Vvj4p+w19mBpt6c6uR/no6ZvRF43CQi0rc2Yak7FOGQAJ+EapVS
CoN8Y3owPdWs5LrhRZBNl4CXaSJnjL9SPJBdLk28OPT6+gdUjfZ97ey1RnAZD0HS/FZNB/mBuSnf
Aoi/pu/8KyGeCVxucXuRqGn+e/1XxiiSAUwQedAfN2kXXH/QjAc8YwwPz/MHpxeoTX3L+x+ncSyT
UcZ7kj5+391/0qMiioiHiMd/Nq80YNd99UMKf+kvui21EfSL8jKLwi6zM0Yazy9X1JHi1N1SuU/R
wWejXxLGeJTvneMwKEtT8vb+nEFr94twYsnr6jw6ADzAm+61kSAd3Q0JwbRhS3WV8xdZaMPmMHYM
93sfQcyiVVXSq4Q2LznJpPAMWHas4TISN9dA7esw7uLUx0rBG8b4xGC39wb4Q+CfLHFI70n1lYXx
cVMsNbCJjy63jMqHDKn6z6mcK8X7Uq6KqJDv0qVI5qgIp0dr5DMGLdkM0HXpZC8+O8emeRrPl8FO
sWDT6jnXAJhN6NH6HgB93+GkLE41Lp4Yn3FLnUTVpUkhAvj6+Isau9sA5gQDCGLXnlHlf6crbUoB
UXDJpZGkuwR4+VbM0qPN1O4Dc2IxFZmahZFNMJSolGwc0Tx1PGYF6qypX8rMUn1vB4XqPHSw16Pp
Jk1U4kAsZFjpIEiayf1To9aX1RV4X539J7wDnbbno8RxM/w0SFMKEosbpaCzOQtD39U44u8YgzJk
S5rLc7OvY1IoNJ+II2foHtV/BO5oy+jRd2/aAM0IWnPCQvS+arGK2mhAsreff6zCOwY0T46wn+KH
X9hpL7oCiDSfonuAqmM+lseWallY+5eyVE/HguL+Y/qAToBcBBpaxc6cDR+hiSp5JuwW46GbX6AV
OurJmWqXq5aSYyH2iVvt0iPlHJn7nvc3pUB3sZemEJwCBMFQ4poSSPSbpp4RfpZHGvorvw9pUNRz
Dvmsv9dNmxaex576s5LwGRLGJDuM4b4o25M+ezydoz4iOsQf5uvw828NsvqtYzqPvco6ESbYwsMN
fzjKsFBfMww2t3kXhcsE37N59uJX2uU1CBYnf5UE2NgNeNadcCumWqHNEG7Gc472dOFgTpLtBKZ7
WUZm95Xgz6v0gACwlZTH85vE4WfF/tK/D/1Dmb64Va2aVHemqKs4SSrvKez0uE+3gZs/PAaq1cC2
VOtUTNXpm8xnk2mCjVPHANQPROf1uf9q6FRiZMoQ7Q01Gk1okKmt4xk2hOIqwbH4azlIg9hp4gEt
Zw+K95LNxQOvwasLosYdv5N7WuPVpV4KkXL77A45L73aAb7dA6i3ydQlkXYiU1aWeD/ueRPkH/v1
Gv8UiEb/woBgmm5wvt+um6BrXILJTmIk0kBtpZKaNLGe7RJdJAyK9RcGZROSf13+1Ts4GOhErNVc
wBcwJ5nz2qXMh3P5sXXy9kspUfNAZceovSWdMEvaWQNYOp4MwSqmd+X73M9n9QEHGgbLHHlx8m73
KX14z0Cyicq+PwIiRFHHOsNvSD0ppRTHhwRrssfF40P6ZTD+Hm0xn0jZfhyerSVO86DFTi3GktRL
WgLobldUmCXzMEcdDtGgfwrHPIG0gqs9EsKgKq67Y/R9XOP5XsJr+yeoEAX8BLbqS+4ilzAVy8x7
PnoyYWA8mftq4g540HAoylBMaBi5BSG44ysUlPavtiPM0Iv1uIkNX92lQFfaM9CYIsm1ELg7xVxR
rVzrrIG8WrWQQMR0Qxf8wVH3N7GMa6Bpuz6mfIZ0N4E4qJYtttcyUCpYhiKkk8duM+7GK4s/YQwf
4IbYwh2omuvE4XfKHhfUxsoJZPPk+lzvafXMCTqxrq9cQsbPb5MFTu0FURIAA0vwmSNqma+04Li4
ENNgHf3V/SaN/Es3pzMJ4jAEoYqu7l0CVViPTLaqzhINW8UAa9pKrcPYu/NV8taqRYUGiiQxwAvH
T7go/WVUJO6v5qx6wa1dITTW/iXjoJEoiy4FHO628pJRw2RcZREkiS1k5OptvgfkAaZmXVqdLGSp
dPAZjRCnmPYC2zzoJ3lqdZBu4aH76My6SPbCeXA+puXhNMoOWyTTnGy09ZZShwyiKfQKY/O/qv/G
iHZ3wvh/iF9HsAnBjOkFjic1WLFTDumOGMxSiEz+C2WmjIKsKBeWAjz32YZu/2Pe0QpzAtyJ8Clk
tDyy/e9108zU+9wdbxgfKzDFW1HmtY32OEyjDEHRd0pw8hBR8Qu1r3x9ufoekqfjBqn98PazoMl6
WGlvhPTVj5xkbNeon41E1OQS5Y/8Nv/JWeEmGGWJB5eaFgf6XrRupRCiaiSLkPGJ4i6JovX1Svbs
Ajdt0DyhOw1D5Eh3bw02SmkD8XQJTl9cptdo5Yn8O3I4Zu1aoFxZyU3q4xIdLd+xjXUhUvilGzBq
ckwaWIshNGuCwPlmK8cAbhxdNYHSGW3Baw12Q7V+ccKzvbJUTgxolasMPCdtZlvQI3w7HPhQr+ZY
EB8V195xiOkpRUYS18SnNW9TLEUr/ODc3KU7mzqnu/FldSfsIUVZ1gg6lHlEKQfHAmKGTJUvcxKa
bqbhsDCKYC6vlXIkCWcxufLpKI3zSip0DmtBw3wQyzN7gHG9uaqmA0xQ4/ScYwKRs6BeuJDjYkwN
h3j0j5uBHQiq8+UOKsXIOFK3Xv6DJsat9ASil9jgKuHR7A0xbAPEccCGy+RjidV9HL9wXqGuQxgg
i4h+gjsVckmce93LPBbGmJqnlN1fgPS+wHippwBF1/H2dxQJ68f6xCN9jAUcqx4U2/hYTB9Xy4Rv
mZLf1vgpu6o6PJ1tK2KVdu2K1IZDcWARaAZ2vxh0t5N2zMPw3iCtrR9aQJKI00gs7ZZDF9qQ6N4j
ZOuCnyz17sRwn6hCIAQDZquTgIlNtFMKqFARu859sVE0khY6et79oYwutkAzZjN1eQtDBymqXQi1
j1smv8dN5TNgc+ha2Y2qV12WluVotwsnsZmAUginK1oKkkOWEVFFEMMvLmSFNCD9Jeu3L+GH26xO
ssmgpwyJMqcFMWdGiat/dh1S/O3WgwSVPvkpyubvoztunwGX9aIKSskTFjCz/Dt1HNJATIEZ5pFE
19dd0yhj6bNuRdRcE1BRX8+hjoRsttvj7AKC32oT27gc3PUigKrgh03NscK6knFVHu/XgfufKucX
LDdetfvYCxW/iI8rR7+4DwoHlOWYbWuj/xVTJhfQ6uxWlnLKWiJngpZNJrW7mVjkwf0pjmvmL90V
eYOpCGuJmSTrakPCHff3bHj8s0Az1x5nL3TWQOQvqdMj0jKJsctCVlMuRu1wJ8vEG4nGBRd8i3BM
JAOYk62tdVrBQYYguKHmH5y75SpOSVnS89cE+hhg9nmB4VMSuRakIMDpXza8DvWMYGaf71J+WSmu
btOhbKqbtRsHg5xb+b2f+xsmvQwRKRXjnHYGD0J4H4YBhViS8o2/Ux6WtHLkn8FJSL+MT3MQk7OK
55hrWCFQBLW/JmSDDBBvniAiwE92lW/GrXKeFQPXOvcfrZo24Pc7ueTYRYKUqJdAl7HUtBKt9ZNN
Fl/NCyoY7/Ye6y5t6Hpmik/419rBkruHIU803Hgjbq4lV5B8pmDXtdXEbplfBNhBlLSJef5JWOkA
6wCevamDUPjS/EsIyvWaKge3+HOKUuTyLUj18/tAmxEnHHXtL7HrVsBRjgADRo1yL9li8TBIAt7p
ARddohmCOREiwgPFvkUVbohv7armHP5tfvBa2DDiD/BTSGO8Ot/Gw/mPPUzgIqRE1TQyZrAoox9X
VmPHaaqDVzb9rRjHBk6Lasc97GSwO6AnzfRXo+jjPwHARG6fE19dyTdFU95r+iPWbfg1kmX0Naep
kU/g19zD03tI4+0yuQ6MtLqxKAWxD96VjA2MlgYS42fhEjPzuTRCG3F8tVH0JgknV2m0BMIbtTPG
kZUFN6Pzpo2Nn6oDY56JzBx+5Rr3IKuf9LViRjgT/aRzlvDFfEbSWZ+FXU90rHt3/GJ9xFaOvnAj
jtMXFNT3DxjUDUE5CBLXLsqse+0keLItiOe5plitXoN2k/8d5vm2UbG3V9asnXxkfdTtQ5AzWC8q
JhefBAkRI/8O+WasR9yfTmplEcr2H8Lz1vzB9sc9+3t/oSJ9yT61ebpC/u3nyNWzIezT/HFpWkrB
4HBK/JeQCHplArtCpCxLXxuF3ghvsJU4tW873uFzIjhEUKiD6wZTePrZCIqZejjy6qi7puOzsP5M
DBG1JC0IRZlJlzbWy531/5YA1PqhxE21/K3LESRTTiK/H7FLq1vi5tpXDUFQlzF1vmNCVTAciqiV
PUIRrHWjeBXbctA9xf1boWt2RDqHSx5NSH1VAVS/n0GKnc4yjQTK+njflmnDdzdVhr0kueRfD7j0
gSOF2WO4FRyYAerlLEg6+iwj1Uw99coNwxBI/MPBVbzfLY460nhoFTF9v3LrTmDjgarIuQqyr0dK
KEeQpg2rlw4tsmZL6WtGUYpdDtck5GAVou1i4mArvbDluF2bZcC0+91xmcLMhYhS0mg+fIg1uPGx
bi1I7sNmjcVWXXiDXjDtEmy9vSCstCW1i4usqSGdHaHs6fm+MHexQOm9I853mXreNQg5xkvNWu+v
ef39pLDft1skg7WFbn5ISfnH2ODeDO6tnMXS+tGP+OW7E7YfVlA/TBAtBVRZLylIeyhQxHKuI53D
zRUQlhRCJcqTi8I/WNM6MLvx7uc8WjPshsLZAW57d2/TVKJS1wdBTAEvSnAoXuMWlCmN6W/HnhuW
Ay7fFqt84KMeMrVaBT+cEtOBNT3AozF8gG1rrxd29NjA6k5acGfxKsBw5taI3JkNvU9wcfEmgcPj
glaEXgrPqeKLZh1lxlPi3OAWYD9n/uBxw5ng6q6WPuZSNHjrzZsmPloI8FUbJd5hKwpf+itdJx0W
oDMtUtc92/2LsNy7BvYYR4IV4UC8dV/8F44jGhKlCJZHzuM9I8Un5/zsQ0iDg6AEs07/yJV+cE+S
+/bTfmkfMU9ml2nq/zF3nA2d24NY/tnN4Er3rwDLxpE3R27u9LtuaxpTFufP3YPd9+3d+wjFKIxd
hS/vOr0j0IZjRGdAYWY/cHzpHhFMJsiu2FIBaG0Hx1aFyM2vlyTexkEfdNXPO8BkMb8dc+bKwbxm
CKqFx37Iz4vz7RSCXg4A9ZZWrthcQ1pfJzHXi6i64l3LMjTeNttGQBa2BPvw5GOaceHPImESvqbp
blbsbkLqEMCIvH9vX7uvegQ9/EGba2IJOwjfSYOm1WAfOg1UemMU5eJshNh/oisbrlWXVrNEjWnI
7mdXMGSLhrZ9l4mJm8kyROTtrLMvT2URW3OEtG4WF6GFAUiW9+G2JR+/ADuPKxkJ3S66QI0tn9qR
harbM9dnvLJaX8Tvu8EJiOrSjP6r4FrS2uxP3KpkLK4J3cQ+2C73++OGuOPfx6+w1suY+4BTN8rq
YMHJgyBglPh954d8OmQkCh2iPYYeYWrhEEs+YBjoYalvcEUmjLyxRBVycCtgGBL9cV4BEGrnuZKI
7mKAYXQst56kMV2oTOko++Cwt4CYHN7vjQcvVk8dx5XWa/wAkiMRbnv4P9fizGM1+GNTDOaG98E+
Eue98M2cpYJpZy+IRk87te1IiL7ZO6rbQ08eiXJnJhZ4xreTRov/3Uz0UpgAmDb9Lfb8aFLr9fo5
xsc9ESP/bDKgwYdHGPGBy8ALmkcgSdDIDjNSEOq4b4Y54tqGpaJU7HMXJcoJTy4TZ0zsbIPpnhdB
iFc3JGTwuQKdraqPlqeL7Hda6WUbRM/7xHWPEmbpjy7VaDzZ3V/IuSBCfMiY9AL2EhclF4ZDCwG5
L2/aritXPj40eGnnCSgBgDpD20NHVxkZSJ75GARhklzveYZ77J7dju8TINuzYPRbqpFAfiT+7kb5
+8x3Fa6iEPyJWN+ZBFo2UnvDnUzJCoS5Q3Ow93yE+JRCuDwQAiFLUcQ3pK/FGQn2gqOxqPAu8oy6
uQfGCnOQzkQ6lyu1VA92zY7IRX5DyA6XkVPhQAs6xh237bpCmDsbqyNIMwfS2aL890iI3RsvCb/w
5kJ0rm0pkUSgoemK+FFmYJtPMJeeMT6eyQD/7pI3pKhCRcD45cwogDjBs3iINt8HSWT8egb50x6o
xGJdqAU7thDxlHaWQVrpZdGlLHKUfxKe487STTb5ffKTd9XcPsQWIvDTTbnRCseJTIV/Oct/4LDS
vBtIK9++GMKxy2Bk/Ja3qKZPoDHQVdsTB6eM28Au+oJXHppWIsomasVgLs7OdpGwJ3uaTlMmJQYX
0HyQ59ZBegVtcB7zt3mWmXs4CYAR4Wrljn/yXPKqrU1kGmt1RgASTCseRwjP/KqqV05BTTz4HPJ4
pzPCQ2F8Qw1GLNBN6A76/M23rwX0SICcYrqNnMqYmMo/UHI5IzTnRYvOM33buJp6SDpDBjgR/PpL
2SBdawUMFhd7xT6Nk5uSjbWYvrEhOu+1RPIIYdj5V95Lcwan/stkPGdAZDivyp7ho51116t5ezbT
0ho/2MrnPlwfFuDtJu8FjjIEebcGCi5i9V++aGd0EjH3wEHt0cdE5gUGq0TDpKtMhJZIGPdiPseN
IGPOuJkJEG5jiAs5UCgi+DnWwSNNjZfxG9UEGVTM625hUY+7n+qNqsTyoOY/hLR0Inmm6P/luC75
jPNLPOvbSPuLDLZ9HyLtM7LBySKbSvS0i/5b0MyuFR9Wyz08IT2i45EBPxWuqteVs7LcqEZFYbQb
jtUR2BhgYaSdZacrSswhxfZ62TL6BVDYPncuGIh5jicGevgrMJh7pE9xmHIKkusgngsNvAa8YvaQ
OjUE3poJRrVoXWhIf8Yzp+Te83ea+OjFi+sKFLDZHxe2Y9FFDcKkU51fcmwNUfVJNNAgGbOljbR1
+IZNkP7HVdt7nT/d8Qc+yfDIpUWVWQQAM+3vrzdZwNpX07CeCXcH0AIZYG/z9IeBd9Jffy2gcOmL
NPqoAhfXoa7jb2Byz1R1XV5Ctk67KQ/sdyeC0pbzGQKWE8+om4VvZrArWT5hqDqrQDFlLJCp8DdQ
jff+cwPg2HvcdRw6huPBsNlRm62Yg+oxLa3oNm59EuP9tBE85gRi+z7AElRGildL7kNll5gTI0Vy
Ue9jQLfvINvn97QSZMvLz5Lh8fGKfV5wnfuIYKqSJbbd1+FSbjKEpjb8vHrxs6sQ4b7D0wjG/7NI
0aBhgxZPjHFiV71UH08QkI1oReFO/9X6wBBBJqtc1BjefMuEQu+7PpP+ThHuV7/3hUCv6yrbFwBr
pBUe1YDApxwgO+IX2aFJGuee5DpAD4sc/HZ1BfpVlmmqozMDJKdK49YDCDisd9J9KjQbKeg6Zu8t
HHfSvQfSBOeb3UVbIlxM7VN+tNNUAnYxKOL6H8IGdrCgiVHvgx5Mq2fv5Sj4fAj+n5gHIYN2tF9w
LmOODq5uBAzzBVdhojLBt9ZAxJYl+SBZVDdwAdEuiaZlSQMGMBjVyuxazMMg2i/mS/OoiEkpRZW0
5pgoUL8qQ49vqemHiYBlS2EmqPYCVHEXNsGMT8g4hNfJK0erpW5LVg++bvCw5kMNjuDj6wJGDZ1M
4KzPMSoE3cALNnxvCw/LOdGskoBuWiWEaZnargp6gnNrUUxCW7Xd5idpeV2dDhVHLRo8Gq6NjbhO
U3ekl9kjfePMe++zzOo3GXPcVhciUvg/zdzILqvBF7jtmOW3Gc7YP+6C70+Vv77vKacbY++DC87i
yCM2K4chwTf7mq2xNrHC2+6M/JRJdGtL/4Oraf4CWdorOfMIumLq1UcpCnVH6+5AGJ3EIqLawcDH
fnkvINPqYsyXG1l9v3Qw+UWhVtPSa6Gk0fDlDix5CdcEKXu8dOUVB3pnhddPT4Axy7ErUCJ7Mm+9
M7gBaWz2aFFh5PNYVwLY5PeHJYWw4ivRkhAuy0O12W/Rh6H0HZYXIMV13ROQmQ4IejwHjQpVg5RG
R3OtzmZZQlALoqkqUrcaZ6cd6hSQwB/tRwAIamE70pjhHgmDs6xxYcTkBaN/7venmZFCfyKgoVTB
nUBvCF9UP6gw2YqrZR1TCxYTYmBMUGszK5GQVsRFCYf2dG918noFVP7UqiurVlBpBNuxdDe5WBTq
srADCsyjgfDp2IHF/COulRcYG8EJAeB1obuVSEmOxRya1aKT+09HafMm5CEX0kizRgDW/Y+yXjdL
xrUQgdkb6Kiugnz/MmxJic8MaPZhol1VJjxL20py5ia6ALZkZznahiFt7qOT7kTe7eKbq7SBhyG7
a3R27eqFNcMVw5ZOE//DIEFbk9y3yh0Wh/7sZWQ+KZr4gSF32Y+I3kW6DwWQAqjVu9px8XpkvCR/
ImTtijN9pUJKk2qvVKGIHqiA+oHNADK0AOXAphOO6ASyAwReDPiJOTqpua/bYPbjKSHGjkrkl5TS
sIOKjydXLKH6YtPH9N7ztBnZB3DfXLSrPy4+7zaaHWenR0OwazGn48K9M7/npErajadp6b7fmj8E
ixhQNNdf2Cpz0/AiCjYimNu/zo48Ow9CaR593c/bRTDOL5zbz/2HMOCVuUsySj9oX5Sv1svj2Y/O
JQobdyxaTgJXOnlHV5GmwAaN57Y0LkiJlJneW01NC0Jrb9gUZZKbhrXvOUQ3UnvZ7SBJl94mK4wS
AmcUDyP8JILUorc2c2dEFTGARKrykoDsOEZYTpagRQ9a+KEIn1iTcLo8tLWjhcTnB1xzPb87PXxF
D92LEs7ROD4QxqYP1xJkCS4UALBkHg8ibA/upBmXVRVabx6FIjGXtLiCkUSJZg9QSWIv9WB9Ay/m
cEoNrUY85xOmVgwjIxsRzlPH9QNo7XV1K+ORtXclrsLdimSqKz9cmZSGhLOwIOk9e8YT19aDbX7u
KUSQ8TR94bM4mWsJ9KvBAO+8xhm0GNDxBotC3sErWH5xmqHti5hBQAA6o8yXu0tfXf7jUfIfE4uW
Qn7/HZtZMgBaFukfONolf+15vg/VrG5Mi9nd/1EcysPCcGjiA0SIuORnUBSwmk4okAJBt/diPDsH
BEGvo3iKp8KxWNYk78BC080DvqGNJsopcDerp0O81NBhu9UliemPjXoBEzun9g1elf10DrF1hIya
FaydQ0Yo38o3QnJordSuCEQN9ZI04qg03Mu8xp4IKJzsjRyvkKu21EGEyQW2/3RDvxGf7ZTDL3fx
B3rYS8FzOLCpguGWpHqmaYQnzMMIdb/8E54bhqXiphM2LlHkJTTKysMcedbzTYj9KV0wxSagRQA4
p1Lj+zyhNZBzzl5q6GV9IkTlfvyib24bpnowE5Lgo0d64SfFDZtMQPNv+bHuoJ0B0aGFRtwu50g5
ZBN7A0v44+1lopLr9AH4HpixJzhuW7ARllQcvjOiKnCuMRuIx2TaZGeqJalSqMzN4wz1YjpAT0A4
mmTF+nxw8NJyqodXpkGLGBZ60KNfQoC0Q11ZLgUmLYtTsgp5mmuZsGBVXF+HfeicvCwv1HEoKWpg
IKQV4lW9k6nPKWksVqjAC3SbrUgyCI8GMh68GmE1G5t8y4Fh6DX6JViHMosPs78riJJdmJHz7/9y
tZ9g7oTle/qI8IP6PgQt6U3cHykw7l8qoYIatqSyH5DN58swjyW8Sy1qux0mc2JyDtj6Rz/LwWbG
KJ3G2HHhPTGd+MJnJz5Rq+I7svKxyGwlR3piZwooWE5FupFyKO37Nec0VLNVKk6+xaDtMwWUbYru
0AKKSgd6Q+oTYA7Q8nJQ9UEfIeMCcXOHJRtHVYdHsY9rLBJrraaCxc6PSQL+1zpZaWoUEtt5dnrz
q7GWrpRwHgy+1itk7rLRHoixyTujkY7o+uZUoO8RvrvzDuLXQU3aZtVTAneja8yz9vE/hEdTJe+a
GNieR0Nt55+nRzKqf1ReKZvIOVlA5bPjUajo6XPa7uScAxO0+C8FYbl0/1iWzreguQCHdlc3QNnj
2vE3wjQu5RPxQJ2sZzhnN/Ps79BapXfRX/epJNn7ksQqsn28jNL6Tua2bNSvmz2CjABnFQxbNyP8
FNdtV02D1kSJ8peKZ7YexSP98GY8uNQEd+P9jmarYyIhEnJM9T1T6wQWqX1Car9XasMdnWg/JV4+
g+jVUO7y+Ff6CIiM5RtiCFcoxmbq6a2mkNd54rTjoWovjo8K9GqDfdrfP7xLOlTVwHFkVsLQUwFF
KsxedWD+06lXdMr9HZgt0ObleMvxsXAWyyyepK+B97jm4VJIB+vmJUKMqg8u6PZpgLhbkAPYGqxY
8LZqVJiyRJer5jeQodBO1rUopPdYfx9587CAQdnXUCHjKNWWYtCWOTkcJbsO+3XXsGoLp25IhlfF
a1ZmAysVNxacwvvS01bA7JCPP1frOnyGvPxXKciIz7hTFlygngxinkopy03PAyaub6AEInNA8I5Y
n0/jxSuTFxgcuzvYZKCPPJ1E6XKEt89IBrWLukv1BAaQ6v+jd68BTBnH1G9ioWucGz0KJnqJqCvX
I0UdueIWZH62ZVgJjpKpobrTMadE44FIp7XKjyj76bnvnyPodzByO+DQgIB5PTLK1PVeW3Myh1RO
AuGhzHJNdBMQAumRsBHbMfqIKMvsgIJTl3bg50xL0GErvKUehDfuv59Mw7KK04gSP6oLtVmsKnbd
5y33cxKk5bQCjtmlNpo8liC6QPj9mBtITlvruaU3EBAU7QYvfxIG1/yNW7Bu26OzPJARcx6NcH+U
z35mVP13l15dUCE4gtW/DQyTh8ZagJUgAYw4lQrt0RBkdxUKKynPFxld8ZOTPpNJ7jnNiCC9ZB0w
z5wkAgTwhqUlqzbwNuiMuMNaRr+kRGfdugS//zTLqrBGMuscnKue/UbToZpvHQSfRistj9YUxXGx
6/DX8gET7SQfJgnzaGVrgIKOmpIDEpElO8IrOA36R8r0mTZqz4mHMDtwi/1AaEMbZMZ2mgjtjHOy
IH6GT0ToNlm28HGs1zclkF4rjhpi846k0VcB7DdfT/ZKn8gxp3VU9fB//zK1FjEoDurUWeM0YPTE
PYqroljXb5dCtRLWJtozDUgYrHlKg9Coe0VyOjwgi9H6cAY2bTBDm3n3qoT3gKxKNXFuTK4oe4DI
YRvoGmgr2DzjvkarNccbMhLVFjHtAjD31Pj2aEGOflzDJczf/vla8virRyT3d5XUzfopgUHUuEQb
58sE3GrbjZDKuDAZq/DXR2A3CqrOLO6y/BaIW4gLaAstkAKpopokN4EnfYrxt43YzZZqiexiJOhd
7IZiIRU+LklRp8vJ3pmz2OKYbP+7BOyfQPy7DWqZ7mjsT0lhV+3fvgyIXFXOaBhX6AGS9XS+LpZc
g3DBwtM1fU/ewJcPXPXiSqK5K1T0opm3hUYj0QagFWQpGdk1MngvOdLFnGMr0nzqvC2x24FtvIic
bjj+XgF5mivM62NqMYLzCcWLbhTb+Z0lAPP68Az3vJErcF2oF5F+krf0wP7yQt3Po2rnX4NNn+wT
swpNIV937D06FhxEUDuEUoSPl5A+hfnnMGchchN8wwUVNTQvSz9SkABCiPWUKwWEh864IfWkxAsG
mAj2tFjslZiCeWgjQZhL1SRS7pl6CIF4sU4uwXkrENbRw1jgQEiFoeM1jytlxX3nu5HGhEw3oIFe
abb3x1hqCj8k+FFcm02wT/tuqpxcT474jX2JMEict2iA3dCDYpa5m6n4jRB+jn1uN9pnmo53IQAr
2JOQksHmvq2W0YkVQt2EIZWxOhMVuVCcR2gQUa4b2LCjk/JWuHzjxPe4BUPr37vWdwpcz9fghOaX
a61YK6D3AL/7nxyyScUCXs3zQLaZdZ7t6oZ2ejx2FtDPQ0Teg2rNoylvXZAVN5N3M3rpZO0GZR1H
fxxZZnoO93WTSaAPishWVEuEiwzDjIh5h184gV0B+5c/OriAlgyUTcMtbqOTshJ5HnSNVhjxCXKi
BdiW2wpfK0IZisHBste5g2c7YJJZwgtcrIJyBb/HfHlpGK6t0hEzhaZF5scAM+Tdb1TU7dqNpYXp
+xWB52yv1drUsHKj8MMszpe766ARf/t1rSPmOt6Tv8DV0Dk8ruuNOY3gR7fvk+NzLfRl2uka/QqU
XDSd5d1KXInu2Uw115BIQ8cVsey7iJJw05fOSRrDxOaBf4ZlFqJ707WOwkGdJ+1MbmWlC4jiQEFD
mtKLMO3Bgxm6/0SQj3Kpmmni1/kYoHCkziUZU/16RuNi5W4TIspkBfh+0d3/9jaVIjB8u3EX2Z6M
Y4MN6noJ/ZY3cdafzW1Kky4Fx/rxG4tlwj94I6Y5lIwpcZm+vxf9JVqF525DCOiZYAofZwvZvlc2
wWUKApaQRRUUsfsXaoTgCEO5L++51jbLM2mGfDBO8uoIG7R4lp7dAO6CMwgXLhHe0BxQngQh7CJK
tBrBT88qg/lEt4KZEWbs9B5JjpjQZ4/sSRTZiPSNITW4nW2a0GGmFblVi8S0ZVOIpO8W746u+tm/
ulvqz0kXoZt2Dh6eRoPXNjHcLa7mCInVjPgF+HIH1Ss/ncULTtLfqtREE55jFxNAcodZyUxzD/K7
iA6DgC28etkx9heZoAIPXEuYDK59U+7sAstTw/Ll2VL+lDMnfWPyoh43KFGZ2YfWwqoIErRdLXoE
F6vPcGGFYtvsOwaNiDOECJXVOpRy0YJXSz+ivLOKzQSyD7oDD4/lRj50xKhQsj3oDV9tj7MFEBTz
8r9nzj1y9Auef176D6otBrQzx94GLbGrVFrbTXlSKytVbNEE+2psytKPu1b5EtE52oJI6jxxQah1
m3+fAXx0v89h476acSr5EAb6/Ooho5EY5aZGrCmPbowydPFlpzlpp1oTwhhZycurr7oe/StXspn+
FN6YZWT8qzG3RTDDVggveMZ6hZJYarR73Zz2tiADaP+7KIMjUfhrH62DL+ejf7VDKWx5d4a3QA9J
q9zes6E+MkfIU9GqyF7+2bFPiMS3jrDETYu9xV6cqP/tb8YDFiBVuKSBDS5JCt+WNqf0Fvyt/PN7
WQZpirbaAKsYdG6gX4Z9yGu4gHtuj+RazL02rXihRHU3qKBa9XZG1+wdPIj2/dbUkFgEaCo8rsMv
1X/r6ps8748vx0TDkeG90RI422K8QaIjVpH/ht643VoalMP90LIhpWrrp/nKLBy2uFgw2aSp9N3h
uknGWEVFbhGx+9DhnNEtamF84T1nQmMsZlrjMPW6ZK7pCgX2vBleChHkBN88+Nm84ltHNiFy3b0+
af55IWhMYeUGXufCsrL7nfyexGUTbUV+xVxnpTxgZ9mW1EuvfMABxfp9+FieffZVZ0Du3DeeDYB2
jlSxEcWhyMo2IK6299u+HJldDP29+hz/hqjftY7jSerqqtxGdmL6kXjJA0tl6Fy+mEsCy/Xsq3L6
bQDon0meKPzv3gKLhYqQ0QCdkVJ1X8XzALRSPLxl+tTuB13O4vMde03clDOtJluW3TOiMktoMvV8
YAKYrPAI0bYPBKszIWrNAbfvuF7/IKGbflF9TOmX1/KXbPqXynUUkTmLvF+TBT7tMkujLPziN/98
EnOxRurKR0GDMqOkHLR5waVHm6J8MK6IXzboaIu50VSNgqxzE3Cdzh/bw+0DZp0e5UmCzzeFtGJI
ssZYh48/jU/vhbmrTytPWASbmdt9TqJYmFDqUVVR0N0B03OAPIRzGcvSsUcNPPPdwLOEBJUyLvq0
Z413eSNwKULcxteJpSmJvKMnMQ1zVP6kId+v9iixKsnuUqhmPhzKxmiRHVJIQliY1w1VDDcZYWQa
WB+YfuANSN5Amo9SRETolAVyQ6iDXths8n99wuPLTVD/Wv+krKFAkfwyFlQ/JLczgMg7TtI1uEIt
tzn4FTjISotOtYRzsK3VHtkAGVrnRpCa4E1JO7lbI7mk008fdLqLNmUqLROAPl/0q9On4MkCh14a
bXzePNiryEK3jDRLap9k+l8cLBWswhAZc5DaG6mcsT57ckFNyljyWggMc+ul3qkO9TuA2nEwVcsI
tIZ6u7Or2O0mFsE4qdZz08BqLMBzgGQi7GSP/SlhVHwlJ72Njn8AJLl6DyFd5vL3WXeyFifV8p+a
QZeUGOTgiPfK0mfYf7Kg1+rIsIpHp5gNqquFecupobYRI+/AEjns8uReRkSQbckV/76z/Q3oAqJS
VsosGh8Fi0NM3YSMVAeucv137kILbrYeDjc+gAS0WH/HPhr1hVuAO+MYmaEIia+IAU1rkFlTUnCC
uwfmkjGLwNNAHoCFLUvA6GUdGM562gpUUcxADBRAB3tHZhU86hSkY08Qf3DK6T3x/U0SrdHlb08I
wG/ibpgglYDUXaNe5u6NMY36OVQpvj525ZVVAoYkVD3adjK9nCh8HUtnJOB2VYhUiM1Vh3C6PQjp
yUpDBvKqF07L4Tf0PnhPopWZc9qItYb2MZdqH/Ev3+ikb4uBdLTzrgOAw16w+R8kW+ccSfHSOQ6H
5D3aypt45or02FdCyaUi/r8X7WngrKIJyvlouiVBLrGgPKAxdycvqNgFqXz4v5exIzvb4VF+qn/I
s8ElQh+8PYwnmRPbLULzZyxPD6WlD3qN04Kct5Tdqc4uXgU26bwOe2MO8x6vr07hndJYue6f+V0h
sRDgNsBYr0kuRUS+vSU3diBqFstmQs//6eQM+KXixeST3jl5u3PfSkvjVEwsjX6ZgBQTbOfeuALG
NOn9fLQdDauXP9t2xNFACYAH9HBvF4WNwbt98KRciG23fK17hXtwq0AizPOyHKmS0rco095ydYkl
rq5gh/f4OCZzmrygwK6bM3wyDkxPUxSeDpJVHbyKnPL+C/2vzyWZwFDb/S31aLvH7I5ySa2pNRZU
eWphdYoOSgEfd6NnxK+meqy8UErXiS00pfDldjzXQdoPkbxl+VYVOY0kqkghjl6yTYGTYlvjkBD7
ivn9qIi4bKvbSpBIqWdtUi5DvzlR4FwtzIvjeGBh6B5KsMif7UrOCGXDAe3rc/ld7GFKkIxSzCNL
5JkBMWrfld73yRnPZj6U+z7V0u1Vbq+bBMKOF/JU1bv/JeZ26fiQonl1eDjdmUMGxyoRJIIKvlM5
zfaokFbmTEf5cXfZwAv0x00Yen7N+qdvD9xs8OBizuxs24YUlfotrzTiiAbWla/W9hL8QDQ8z6O6
7Z1dBos1MvpP3FsUxkQ5mKNzIH/kW7qj1zJLpwoUQmLdRhCoz9G5chd4bkSs6wLvkkwjAYUX25zr
crCCDT05AUU+sA3nRh+40TSnbasmQtPugepQ+U7NUEGm79xqj3VmprN+e9VGte2JCG4TWPm1skQp
XIgLUuEMK8sqJkibRJRkm1vbRBe3R9NNTEDdjmRU8HXa0b1Zsu+rARJSXTU+kFps6gaGSK/U4N/+
tbVTGRgiWmhpENIK+LCA4AznZW4sGK6Z9W5EFqSRl/8aEIqzi/tB9k+Laojg9S9FcvIa0gpXlUmA
u/MQ0hhW3PrsQ3YogjxVO71u5zc0u5QyIR1uNK2rJAbAMiQzvWCj0BkSqRaVQZj7rT3LSwv0pIES
eOCOlJRk2zF5lpv51MHL0XfQOtWEYVjCxrrUvj1PPpiXtmYNU4bodC0mbfrwa47vr49X99BkQbuW
CHVCO9t4y/+f376t/uzpTcO2BV/zSj8RMklDAQprU+ol344qRZA2m5eL8U4w36d8HjgsLjDuGWsd
9WrJ4GuB8/F+oxMatgHzhwL4O+Jz0CikspV4FWi+tpko20PTIrnOjTsGFGSEaMxl41Pm7O5FsOsQ
zVgwTD6BVQdQbJUi68fXB7wfZiLvB/NzB7PQruuRWKgAClAe01b+DNVHQuoivaTyc62iHkXes//x
VQMphij3trEgFE5YEwOabHyPoS9HFln62fyYGBLOWX77pY1+7E7GOz8KFiwCwSY8meZ2w9lU3t5P
gwwqkEdiZkWhmWYIH+6HfOtVf2hxsnlUyU4rfAlWFvwZgtUKbvUclYDcKFBZOcTdwHVTnuC5wx7h
ClIOnHazGTajZmzI8NlC+V5rf2d9aGJS87MrLcZEv+AFHJhdBeLvi14Joxut8PeG0JZnFdTc64j3
68nQrz3XWMGlJzOFOwN5kH0AgLsslRexQ/VSjZyfmPvpvvwgQVcs9uGvAWqUGxt7V+VFZovlSgun
4t0v5zB9FA5mZdFKrCjBZFCFXeCURukE804i3GvaSVqfLp145HZRa5hzPwxCUFvgz2lkDn5CxSFQ
DGN3NfD9x/BWOAmtLcVq5+NRfm8Rnu9Nun0n6t5mcIaH4MCnqYIBALzLjSM5H+4sSFmRLVhxlk/w
4FtTYt2cc2ZITtSvNR0pxOaLp0lGJXfUqhrDGPTXggb4vS6E0L2roViOa5OYmoqir+s4yDUwdN5g
TrdKiiQOBDtA9fNlAesUIyRY9kYDAUtpm1eTasczghl/jfZoI2ikzqVdIKbxU5ahVRi3tbwvJDxv
2oDQomVX60bm9dtaVTwXdbd9qwRYnCNViQQQWZ4BnI2huROEhNfZeZYDc0b9eYY3g8a3OinPV8fi
8NYAZnH9zn0xOiMqfWdCc7Ox2b4fCg5yqF5eiKzFh9211i/OkdCt9TRfgRaiClE/dIxO0bu2q67a
IUW7WDqhKvH1FioQDiEHB7rEPKYkGVEYLbeEi0XIv1AWWk1Q0wFSO8n7uFgxJll0gW7MlTW7j0Hp
v75ju2WXVhLFla58WbZqdLvCMKS384wapGF6/nL1ambRHtgx4kUS8wJFnFAQmmPoDRhchG6h3JcF
jHWQ4X98z6l3lw0jrZiTF/rNTuPdTd9aX7dr791StrCiBF0k3ycwp04vJl2uYsEDwlMaINby/M9u
heGNHy5xeY3k4PUNJeL+og5QhJY60G8BTb4fxBWkegOqdXcXjcVIFOlKpIj4OipxmshCRpQ/M1Or
I9vjnBSfgt2V68XYnFaZ8MrKGGLlQCUa1wjG/TtpiW5oCBrduqnYXZVAwhu4cjQn/0pYLOrEVVvK
MhUl51ldeFeN5cGyU8NB68YaiEbbhJL6xjZO8mKBCL7ccRGHoJkjpLynruLZV669tw/ZOoobvXrT
g0k4mul+SCV/2c5Y+9QLfW08yKTu+ID53Ya92oQnYfzQAHnciri52tLFxVaCanLNLOQm8LwZ9XFf
Paam7coxpOcJULdGjiSPZzMS3GpjUrCi2U391OAp6TrmAOfUSOr3QFFG/nR2lK9cVqYOliqU8Cjv
/Vf1rYDUUoCdpyvJog+FmJPj7vEIn/TvYpZn2rjJOhsPyg7pOJBv737DUBMPHbtNevpxeJ2Txagm
cjPFJkoUdq2Xvf0FlvGEmkXkB9Fsl+BVzAPGF2JisNp52HC988YGmCLKjmcIsqf0PlmE+4meaglM
83VtWv81h8uNSNP+q5WjqjK0agG/EdDT/ztM5x9IQzGfHECugt+4P+ZSsG4dTRhqd6/aLrw8iRXP
rCG310blQGi1E+oUOumlm7XCncBK2uoNDLpUBqAYb+9dkh+KpleZWvo6UHRFTl0mE5gOOsGujq4G
4k8XDSUBZKC7g5nHnsMb5TlRnJbrC4Hn3jpcyaxOCrrgOqt/s5HlJ+9oBbts5L5Ux489S8r4lKnW
7qa4MsfqZ+6dPQz1VsBXOyP3f1dOn0v4z2znOOrCeb/BsRQ7ZEtsfpub3Qk3M8eCBuWHVITW6cbL
HS6d2/AStp2OIeM7l7srfOhSxcTkb2S5SnhZQp0ufbUraW4SXsE5hDbgW5K1uBYiETuq8ObQD4Km
o+qqUNQn2jy9/kTBuUP+FwQ/lntptzCVBVYfEXybyTlW2FEdtUbDJ6/xT2925mHbDmR8aRJSDwKJ
zWJbAIsQvAB+vHSw4Z2bUCqCKeIL9KUOttxnBO6F0TkH7jgWykvC051cKX7gfb37M7EKxQnNwRRo
s/vcu6f9iUwrIMSK8zyRZVUl7Ov1szpW2iRIGaMEM+7za/Qfd1Pk+Yz3sukSub75OvdZ+BadfgCu
grW7fsmVRzazpsxFmZOaV2LZYN8aCxXiNnBEO8pq5gvYnirPRm7I2/VErcqWMsAh+80Jr8WzhxbE
PiLSaFAZ8m26JXigiHpZyIhaJCP0JnUD372tSeGhX5mKmDamM4Hi2xm4iFnr4mHWlE95msXxQFDG
G7nq3pkBIzqnYDJS1jxhBNBqF1b5pGzB4jtRHKUyckwy86+GBCsxhNiabC7tu2xLYaJvGy8Qq1f/
EZMD04UJ/Xwh/xeLo+Jt/KdICtMFL2rQG9CX9gMMOckwtqlhz0mOHyVNnta67uMZ6t1APAEm269d
acxnuVWe3X9y1xwoykzPtBKLQVjJsarzqt4X5LC9v5ThsD86imGIOV+W7y2kAJ0e8xstbyMjyHDB
5ZWXjVF32QFgv+HDtCGsYc0SvlRQZGI5zUFgDxlId2pGAoHxT/KvWNfovv4HBQvuL/C7JXXtVE8K
CXq8FjL1dwWilFa+etjR6PH8H1c/KPtVdrDAnoJfJZa4V4vlucF/tB/s4CSJ2UHQ3FuA+TkllMmH
kPP+2LjDT2TwwuS39FbFfeA7sXaFeIH5sRwg7QG/JIezOvaghpEKr2gM2XlaP63ef4DzX1N+SzK6
5mnBr4Vxe2xBheOxCgxhL5vKowHf32FEtmcXMRKq4EOHZ2WUzT/E4x+PD+CJrEx3Loy4FQnJjje3
i59Bcr2qjXE8bS24TlJMpcN4bFJSj1wBD4P4TlXDNP6Zauqlw4lVbty3yjC9rg04q3fFTeS4N07Q
vUBQ6esKej8c2+RpPacWwvP1DsZPTvnVYvJcyFEX/zMNZ05YSck/pM80dFiqEuzWbBCsV2llyshq
FsnsOAFIYZFJhnSHAHgfEK6IWhPSprnv3mHzgouGioLtw/D3J6beTC81IvKbuZVGn0A4L0n2y7Ye
vO20H46WX7hvs+loZOHSMMAwnp/LMvIujo+u/MUdCAY0XmmNWTrJsjyhrNFZMt0k6v9dqa6KcjoA
8QseicyitZbuwuDz7AzHZxMsbQtCoYb7kXU+05h4eg/1SgmHofxg8dP7qrUt68KoFy+My73QUrrq
1meH91QVulgB6HdEc1Ujk6BE1G6J19RQ48cJQ/x2FBPfifLoN2xp4/pnYv38Ov59K6k9iIzJtCVV
jdt5Mi3kf54tvSC22vtlvwkEFU3p8CNv3lZVSchIqN7AQLliEK+oi763eAO2unDuP15zQJ+p1JyO
2oXjybF15EqZ+HrfVa1P7cx8GqgjOgn3oSujS4+87Rn/5UJ5zHAbFlPReW02aCTCYDM0PDu5Dh7V
dmiCksYn9WUNmEXK0EI81v78LxDGGkAGsDqjQlQa2d2V7g5DrVVX4s70Cz3BPSPJRUa0PmYXGk58
qUZhJn34xzWKNM71/0CxXOZppk04UuB0/0gXIkVCm/oqPSAoRHqmb6QbZHhW6L8Ep+Wh9IPmpGbi
XU8Mba30xNOuBZI8heGY5km+n460tR3qTelzhpmOdVRC9rnIirFTLb1vmbBh0ccUmH2xQ/Xgipb8
TCWamW79MhIIuiJiv7yULfV/K+JZzgr3qqpqL7oErXnhWweY9NaXZZYdtalR4zLrRMPJPajMBHJR
Qj2O5pLatykEMuUAKszNNAC0kYOTYeChE2mjf3nJV1oEWqRMbVLJadTygPPBgUGu4m7dnLQCnzuj
EIHwzEZWI0rO5poysHOqFDludWENxzP4G5ku+fEufDnnAKbOmjbe08j/dpC8cbjSbYoIzr07nFRH
q/xmpTY2k/tsJW2F0NexRTsi32eLFdwqt69wuZW7wh96JYpztPG01WDcErR/GGjY65bqxD45QSrX
G2zhFzn3POOxHIb1F8/hKYn9RiDJ5ZEILIBfCApC0IuQ6oB1GN4yqxmbFILrt2LUc3VGIhDGj7n4
JB+jyoNW/OY7rblDPX2Df1Jg3lmSxPIg/kky9h0mGDwXP+rmBEqhMHgJ6ub5kMsIiQklLL6+hH8p
yezTooTsl2+19CskI0TLBYzxDNLBkFOX+Endn7niMtYYU74ThqfDrQsRH/Kj9ZspXnzouEk3gZGN
p1SzgX2qQdP0xeOQ3q11WD0k3WrFjFjHGaSFeiNOgAytfRGczl7qZ9OTOMEPzW2Vp1Dw06JlXpZt
dfU8rAQqpERM3zYE2OTTrY1K6G25MqDc6o5bAtzC5uGjDFTHXVZMswGbcW1kAziRz+ozfnRw20Xf
on/VyMaxkJSwVtr5o7dqd8hrqgzJXR9H7CeCKdfSwTqFcRW5vX4EJog7QILa0GNOjFoR8JZisv2t
43A5ZY8EFyIyyrd0YgO7glRv3yWWa8iUTbeWI9eC901mp/lYm0NkYoeNQPdXzp35zO57s/SYMbrp
DPsjN9HUDCIhSjR7CVTgmPVvA/jECLRwmIKqrQbQMmcE0hgTowi+lPV9WY5+YnCmWVsWx0msJtnP
eBN8yhqoTT8CYXwrhGxT++YJf5CL+4sptMiX3e/cI4nA2+4WUnfjgUAQDf/4WbtObPS+cB6y5ktd
sbXxWb5ycv+rA3b+/uk/2942cjOLKbpjK3We4HoEcLlIlvyXNopiwKXPLvCDxwv6T2Ozz01jyd3n
j85Km9IXBu9QSBGMQZWnPwoFM9BiY5KKMDJ4C5MaGrcCDGPpVB0YZI3xiZhZ7UGXQYN05iNaZ3iO
LCMpTNKQiyaG+RK8pDNM6oWf4Iyw7OG06g7kXVoy3SeyhbvhlUVz07IV0BRZZuBR3NFSx27SgKjd
ncqq+goJEfisBCh7vEFS49pxS9hfM6foYbvbCxwq4i/TlEBWysEHrDUbF4Mh7WJU1bBn4D/fTzSL
LXU/1SPqG6ckhYJ1HK/xg19hBGCum9yVxSImSExLY0z7pFz7zF9afu92ijAh55i4O2mt2T6hfxGA
XzfDr82yWppYOT7y2w83FQyMnx+YoKQ/kzbPugSGUcpSvDopY0eCUoO6jH30nsz4PKvzDCE+IE3I
MUl6lgG2SXLfASUACnBgyr/EPxtJGMA+ymK0sqGKLvxIPA0UjtRhtHKzVHqbQcDAlEb7OqA5s6di
PDqAa4r2dHX8GtpwDG12bKHx1F9hziKucWEcTRLcWb1jC3oF0tbob1B+7QZeKChNfkTiaRcMIvhq
lziCvn6O75d9oy+9xLKdFvWDBvPO+2xTJyV+jeGA0Bdg559rXmXKLLnvR+LTkwODvl9FpeTAOOs5
yF0qsCGqXp346rElDTzqZ6NqooWf7pv/2GEsHo/qgJNDJNHsrKxTDSQls6/7xeM/V0ap0xAc8LDI
Xpb655gptae9EIs9fEgCjiIOM6gOaEKu+GIEF6qQvmaRdlIZwsJjKyWLiPwPNuZmd/5bOpnmsIwp
RaFFhOw3s9B0R3AYp5HVtVyQMB+K3OQrarIOQRjtxXl58TcaIJjGAK644hb2EHc0oY17KBfwwVx0
O5TIEOBYGoM7urQzUiidFYa3CBK63NdrvUt4/dBqmA4yhyW/yjXZaf0owuXRNhqwBjmIsbu7tiAK
CcIKNQFcW9qFcPBBpSUigLQifgAUDBmSIMQuvU47QIZl5v88uaS9a3tbYKbgAhpU+P7L5FKnHz2K
d+PhIRdoRcx1yaVbSXu/OUh5GFz0OYS/vL9I5hhOefa42GXs2+bQdyN+D9n1KEYEidGOJLIA9Vh2
7mnPd9q9tgB36sTkV4qpwv2bOYYSK7xDTzlyvYGfasTkcJm6nidGj+x8lHsW7ApsMnVNe/Y1z3wU
EN/PSzlWJsXiiED7JHUlFspODMw96iRV16Id8BlO0NAugX8VxVtT1Xos+GGqvfNeEseXob/OTGAU
tDMSVMgdsHQpPceciHWcSaN/qJ9bgMF7qLyxvUYexIfRxSMnDTw4jEjUhhiiRKcR8+/Fw7G2GXPr
fCtdpiX6mW3Re7plZ4NGn/OVXeFNwC3uuswa5mX9s15zgjTqVUchkhVQ5DZPDr0g7vgg8wvI/3ey
o92Yu98zg2jgmt4XSoFYP0A4UJamr3lUFiOGzAhEK7DgItbAqguZ0Phz/3JmqTahE3wyXQkLuLH3
zw+tnsvCH/6bdWO3svDySBwxcST97Am+5ajqYwKuNKjMiPNaPTRu30dgdKpUl+E5xrk3O1mJ1/6v
W2zcjhIiyGu2TfX62JlKeG0KeLEH0vYlevr9uSK6sAzeW0p4X5j1J0Cn9MwhMkkyKq+mRSI2GoLD
uyA2HL5MmHSkzgafxZVSUn9vmlCvhSCR2nb0M4UQn0MOeq23Wi87u6BM5Lnr7+5Q2L2MQkTM6MrC
adW0AjRI0QAVhtfK+JhxWnruLP4dnnnHdP/UNx2vrIWMm6n6o0bxPlJ3tGNcW4BHC5QaFtWf9wPD
8wasvW8woO38uKvwjusyWd7EGUk0UkzT5Ugv4lyRqyrAfVHZlZ1RAq/Y+X0W5+AMh3Rzyj0u+PE5
lz/0AA0M/TEXj1PYVpXrjHoH9VXBKbMBoAnQsaoGVX6ujLM8bjjaMjdeUuuHZzRFTiEEhD3I/Ymu
bYWzJhp8QY6Lb7SpRSpPZWJULBUC5bqDbBGxdHYSZLDufnmkpABx6TkHkQkDekkTk4XQFA6FKKEC
mD7aijrqzIWhUZdqI445V75+ekq+29fHcm8yQtAeKNvZU+HO32/RXJa5QIP1fmso/o53l5NldtYV
wR8Plvh2vIm+rxaRHwyr0K/8xpCZfWRYE0SfSfuIjBSxM5V2YFRltT42iRfXBNe79UQG4RY9KOBU
Cljtktfs7nEqFgai+zIpP4LC2X9APLUTPMfD3u4keozpscZei7PvVo0cPBZoqMsruobG9o4mZbby
ZdQyGRjMcH3FpMLIbf73MfdoIK4Vj0EvbMt6qFiG1555DF73F7KLUGC36dunUXyZYXkFOFgawvHp
OCLm/3Nfzv9JuPXpC3wttRvzq2OF+/CgiuyOV5HaDiWSKFkf6CvZpW0SW76aq+gUaVGWT7d35ug4
1+Kd2bjcO4dl2CRUfavyX1cVpYAVympNrpSz/cYgqwyBaRcX6wtXfvf6q50J4ztMsBj7DEqxGLJF
Chi5bxo2rXddVTppqyBzDCqTST3r0mfnWRZJ6IasBGAN+95nWGWms1wPjwCT4RcHUYqc3IiuKdfH
f7Ulsb5y560GNwnM7RlQWKQ+9joMO8eslgu9lIzaUDzDygeUzy+ISJ0iQQzVDTyvWDeSsVKRJGYg
P0hddOqy+hHqYCwFV9F3RdYis6DJJZS2xK2nX0NTSIYKLhL4kDDMtSR1CZlwXMcinuN6kGLxyryI
qVqBpJiZKtnQb1ZvbtJQV1ZjPNKQJnB77ubqEkx8SLnSQG4vDJJ61w9jVJbLgcib2oKWoFT2TUHz
VrvGqaRUZVWMDt//ovkeZXdC4APEfDWknj9W+uHF6cCw80/DK/LHnprqlLdRdxk4ae153TBrHiGR
zPUk4zZHp+q4T3kptArRVOTQVOJZA28wuNIdhmS7rYVO4NH2smkrn0ULtE1Q26/FTm/DzHBOynrP
vzClXcCd8SLDX4Rv9QUDuz6leOP3YdBozSL/Z5PzB2HXFIrqEpQcXQPmSKPPQ2CJ/ZNmysCuvLBv
sUA1fo1OL9+LJrPhVuSKGjzRvxruBqZm5opo0P2clXiTxGGALiUOwpEUjwkDrqLRDCaJbgnCZ6hu
iafnc6PpihQtZiOJuNY9W5I2Azevktv6IEMsGYDrAJByxo8MtdbBd3tWuWp5TvK8eZJA4TGEPnJb
QSOvFS+FVUjsDH8fmUvlK6dSJdEhB9H1QbQA7SNiwFcoo6S7+VQSV2zVJ1lIQOUbNfxfpiykbKyt
XeemV/Z1C2aVoy5inTMCBYwrgglmsbL697vf/X5mpXYXmNkopJ68NySDvgbxnTFhkouzipEW81Dc
leg5nv0F6+alGHQ+jf/EQn7FAL+8MgnSOkAZP/TH0rXOEnMsXh/tF9TdcjwR0JIl7rkG1DndQhSP
E6przK0i+AnDpkqT94t2ky/rFvVgONCv+7XpZz3rD07pwKiZ6A1H4KJMccl/i4XDyFmeMdmrQjzf
k4z3MYyvKslRFn4cC9QiZNDvbmd2H6W1wU5AtFfyrrGNVxGQOAZsrU5k6L7O/0qeDxCW4NWnY6/q
nxA19rAX5uwA2/DgK5HFiuDFYNuXRoZDcNOtVaqfj7FKbaLM/JBvBAPM6ipFqUYr7rYlYdDVJKJj
Ck6uYH0PkTj+ECinnkrTa5BSD8het8u+3lRzQEPw7qLhTk2F/f5Xvv/uJOkptwLsIM2WP9O4zl6W
3C1e9WTyuUkApIEbK2IDXIwJF3Zm9yj8+eNRL7xo1p9eYw+R3RPY4BqkLhCZltcBrjl9DpmBr0Lw
cPqXzWSxy26pVFOZKu5hD/McQenO3Y1N18GEHmPbitqDh4UViCP+a+iyHTzoGxrP9RFGoJAeGX73
OQfdbzuKwAK0r5et4A75qlers8iOzphVf4XJY/gGtNJhL0ywqrFq78N0nl+Mg0NROP1n3ZPztPk7
DUyOq9gXDTULqysQ4Ik73o1XbdbqXfuLRO0AhODtD1bL/y2uTNdbWhz38GTjo/t9pWgVwzfnrRrl
lQ7BcuOU9T/8F5RPvYdfJ4XiGL63lW4CE2pKX8fy2WhTELm2+jOlEghC0tuvx6IO528NUsCRkzEr
u/4rAHWSWU+7etDybLcM4k8ttp+vTdMQmLO6elI4LDrtJwVGnJQ9lAPZLXajZ7CCVuR1+obdU/jC
0SYo9lWsZd6N3ClcAg9I83ULkkHsoZ8w3IrqWZOOs14VW+NlwE8j3PQInXvimqOlMBly3CmQBlHj
AU+261iWcx23XpfLg7Za9rVnRQ8oDULTvqMJc5ex+GCmV89lR6mXZs3UtGTfqaBuyyVnE8wB6ehI
Och0w9Di/INwVHcGypfQMHvPU5U3OYrPcDN/cTYnb0OOA4JPh1Wh3DVOrRHSAdjeYEqqSc4DP9MT
SoRtfAmpl15t9Lbs8y4QSOvMuavPybEywC6G90B3bgX+346xCjV3l0YgNXYKBg/mPEOGATlNG9Pb
KGRHABtsvWAZPNtUwYdoISYEkQQCtpyJihn7SkUV88M9bRRA3qRFD/Rv/ZmqijUnq04hvOjDvRMH
lOdaKQq8OHR+7dwzCbphP7aNzig+wAPKVt8IAN0BPhIu2FIvjdDzX7EZK62Pczjydlg4pHJu8uUH
CgAySEY4SJ9fd8/bJf7UxSkCSnouCdmtd9vExS1/M1cwGiVO5WDWpywlGiVp4R44rRiKReF5y6H6
42f2C5oyCU7OaIvjXujX7+tNfNUoF1aNPzxhtHQERi9w5Yov5GGWUmxIyBe6XPoR9Wxuvyi4X5kM
uL/C8Mbjwg8lUZLZ9YYTrX52j/NIsKz7tL8zEVN7trPIX50yNihZl7YhIGkR0TVeOwSquW/6qYvO
vOc8TxEEImiZx0cpyR1wZhfQ8Sk0RuKTbd3iSUH/+dJpMCw/q6UCnIUXqK9IuNdyfT94Kn1NmmEL
e/CYsI97W/2v4sZNOHY35QaBCbO4s0fUARj9nrP/Oc5O0rqjG9V3PFoU9yjn51mm9dNXNPqTYF1S
+LVQ1SH2pEwr2JtDD8bmrEQA6xFNaMFaB8MaC1hbYH36ZhSe3R8diRkHBV2QPkWWmNuDADgzsQOG
+xfE6ZZuSY+KLkErSpk6xz/crLFCuiRw2sA7pHlLYBf5i0LUXlZRw1yQWYxljQRzganyivRfi/i0
Von9aBlnTAECIhNHbeAylkQ43kCCTKQwhtYLDrayZSOzRpIutn1Raove5ofM1bQ9yTgZ06NhSSot
+SsivTGlylrGSZkJzRMljxeJFJ4rWunoHr5Epjk2d85TGha2Odg0f9Y0TnySCeTB69qgwC4UcJQN
Q4sTI1jwSs0sRYuN39C5xxDeyqnig92mvGGU0FS3BkFj133xb1nLHUq0k1FnO6E3L+Bdq1wbtzQW
WyHRQCYozyxTHD6PtUhgbHMuX27A4HMidnMjrDRp+r9QxEVbf7WirRu0becZJOEhCCwLic1pONip
X4b3mc+6/gDS0qt6hbr/BcDr2UYeGaF37AiV+r9fJ+k82gHYwwp4/EnVFXdKTyvxkyY2f5XtK6RL
JdoM0XplcdVV4klCaJm/UnUmbBisQlMgkHw4lTgmESjr0xztHUbHMGy3E8FIpCzF2+DT5qVLXZPg
F9YT2uqC7zMqWPYz66RyQsPtm6z3P7j+XCahqCnFrbWfyMuNXWWSFTrSO4FD4OzwtIulXfWUOzzH
ps+3sRDtoq5Fn0RrFG9FAtBILcZ+OA2SYDqB9QnemJ+J9E2MSUApOPpCFuRfO7EGhMkpeNpQCxVS
IFVS4jiJHJsvhJuDRkE8FyLLjMJmrvL8uV4QQSAHGiqGRZnWh9BicgQlZSEldW4O4KBTiHI1o2+7
lZiCv+IhiebQdQfyzXFEsGLA2ovZ777lieKs0qjKp4lRFlv5L2pppe15AHaV1SSC6zF0Dhc2jJ7t
Jx16wDEKfXLYPYCpifk9hgUGJUpH2ADJ6lLngNF5Cc7GSA4CF0p2yWzmmq77ISPUw1Zr3wMA8DgQ
3+n0WD4DuuLHe/wkZQUUZNQdPxvGx3xlGqYbcl4ioqGN5TCb3VqsjpWS3cdszh6rvlntNmc3/sWH
8lKpHEOev8iLcr4m5weD5Ky+SR9xiXLXT4lQIZbYgQ1YJ4wGN8X64yr8JAw0xeIWSg7VWQmgdhPH
t7h8FoCBqi3Tqdka0wXkGpx28iRBeASYiCnmg2YStXnuteLQQTkBQZnzoBQuTgvHEQuTw4KWndoP
IckwWNCQmmytcK2VTAErgyrcCpsIK1AJFzMk6FEhbunHc71FmQ82ZztdobCGbIm/ElZir0JZt2Pe
qIqltB/pv8q5qbt0qKN+uaEdy5HSfq3LjJVaLSoZ6CLNbB/pdsL9T7Yn3cle2IDNJ76yZxBZ9yNs
29dSt38wxqUoW4T4NxMRR/zd8wZE7tCVds7bhTHak51zxQwKx9wz5T43OaBPr2llU/Vsy5WXZ1zP
3Jp5mpYFYHX6yoQyV8vCYNbpgUEZr7YtIm/poyOmjys93Bo8ITDYMC/JvbfAyOxdy5lz3VLSq1KA
lALrfgQn8W/q6TLnM/7vodFv3YJqG9D+X351OPRrSs23Hs17OJBlsw8e4wzeaCP5ASjHCSNZYB9l
eLM6mMd1IEiLyeDYlu1RnJ/5OCH5yzWhmnHyFds9ftYdMFGbhrcqXM9h7PXU2hSRUP1ICHZfcrFD
tMUZ9BOW3s14huExCbRJGOUgRGUwe0NvTh5YP5GWYf5MzLUNjTSfIn0Te2GbvuiWs8F8KBy+HyPs
Cv657OJ0pcfggQWwaCOwH+KdlTOfPnONHEoH0pXWjDXdh6fH30nAwGPzF9vdN7guOldyDV3J1FcH
U0eK23HBhNqkuol56zwvgu5rpK/ndI8mCfrpPYwONL8oAOQw/1qAeosDQqE5jV3TXRiqObRCoPSe
TMpt/6S4C5fOm5ecsX/QTXhslKqlInDEhUpiL8pgCroemjNJgA3GBPJAUg0HFl1800bple4iQ7S2
S/Z6hwh9uIj1tlINqXj+H2svCTsosXyqI7YKcrZhFt8GU+5D2AZiR1XUrQjCVK5pc4n4uG9Lfogu
jc0F0vZBgaPrCRG6aT6GXnU/OiP/C2IIK/UmcCpJLiegehcxhd8oBWegB3ODBvXsk0tHx//5cjsT
9tX9Tj86EyB1om2d+2T2QVQmw3oXh3JH5nUatgL6haAnyODHfGuivBSsmhiUxEFU1i1qfkoyfYga
UPey32o3PrgFJJ/CsT7Ygn5PU+I4texqX1lOf6c0EJE+tkA+wcgevkz9BGX8YKbOTWQXlSHXsNNi
qU2R9t2v4eZ3+iHQxlZio17T2FFdCHV5eREvKeeVkAVJK+xB+x8vpbeRFWT+g+eRB1vbzwccbayX
CmK7DSU18FM0Oh1cWiUvvgQ/2gNyW6bzzxNGA2XpnCnFhZ+sz9NlZWTdtfVS3FRlxn2ItT4WuPwM
XosLQjqBk1A8JkubKlrh5O83390K/ZrTfNWtVipCHi/KdaRnXmwbkG8YVDKnScJhCV+1Y2zB3STV
hT8iC5c2SzKigsRJKAnXLu16Yv8LxvgLAD0lJ7rvenUrJ32Bj82H+2pIJCCm5SNH+znYHYxtt7uE
LmtwOEB2u7v1BletqoaWQdKPuM0xp8Qxrz7S91UJ98LKUB4wZYIhLTVnxId7yniku6QWRA7LSFl+
mWan1AybCfQ9VTVq5zg0HXWucWmW3CyD5DhI8ZQjUcHatSOQhd/hMZCfPH1aSuXgsJ3mHgv44sIc
pv5Y1lna/puSGeh7uJxmbC6skfIhb/6lZ9YNY8Dba5OiYXmBO5up1jYSpis4UaiRYC3m3EqbEAej
D+lUSUl/0Ay/fLj+7KSmSjwPdZ4uzlZrRZnLhUskGIV4SOEZD/zvEvHdq/MXK9DWbklb4eqiZqAC
R8MKM1ecXjdKKdB1X3dv3TF5cTrMIoII/Zz82+LL11C9NIczGv3qWdf8pR5L5zl9LkmJkLyadaYT
hPYYfq30cEGEbgGyktEESAA7uvG9QQxgmrobQo82NQyTRNJpufX8VHmDK8scXVu3BjkIL/2DKISh
j50Mb9NgiR88tnYuqw9VTLACQxTubHhluXdS35Zd+nvQqn+nGbUOV0vm3Vz5pqpT1sIso7EmCWXX
N8snQVT68QlvtS9xmh8P5Hu+tyIihkGoYeII8R3wEmOo64X7dEVE3gbSEx5v7pLpduMsRtobXAdt
CUaFErvkjDPhJOP16twtV+X/WP6d5y5FnNPqtlcNmBpjOawI4/5yz6Jb0DVtD6xfuLgi1HJDE/kb
y01b7bnOG7lL+Cvg4/U1IaZ2mcD7V8c8w7BQ5JIiToU4Ir7PwgBRCuox1oswF4aE4Qz516t329T7
D/l1nb4mn/0B91LTf9+h3f6QayO+frkqydjcFy8Cefd9fmSMqQR0dm5E7yRdLmMiu+h3xcD8WoW0
DrBL6VYPcIBKY6lIt1m3FgUDH0gM/56THFqsamZAS3v7VtDv91p6JCkO1oFoYXZzYDlNvvoKZWH3
1AQOeTRmeE3XteN4354kN6lNsIEULzk0+2VltgIOL+nHE6192u1N75x4P9aB/582iQHXvB+WxuTl
504a+bucaQWaol+46zlXpLZOy4Wn2TuHY5vFP2hCMtEYIbnJDNogRiEVcJ4IfAVkkZXQEL1B5wia
8rK28r7ls97JdPKbrcgW9uiusTgSbqfYGklwTRTpYsQOIE2uwiXFAoMVamx6Jp2wIBJwH90DwE2K
TqGHRUwu3ovulTDb+DTak1Zh5Ua55sbAGCzc1YYPnrxea/8IztGq9ziGTdolqV1MeUC5xF8oGNjc
hI9ChhOXGslLE9cENEKJeXoTFiEHeSbrSqmAQoubQDNwFvjcv363ZqKJUZDOah6ATEpsiapXAVRW
yZev6Aujw7oyEJrktdnAMfaayE1r4PjNSUJfjcXQNOJpwUi0nbN2t5s2R4agURooR9FAE6Wq1VAp
/hhx/qbeTDXS4tyApDELkSQxo+PmWJcO5KIaFw0SxgxIK15H0TgsQJjLo+8u/Qg1uikfd069uOao
ov9QYqY9txsIdc7kXhcoNPUrzaU6QJZtEsNwdxjRf3qvFHvfIgnJku27jHU90Z3dEBMvj8b0SDsV
qGmDDoCosht7d3dIw2ThxNB+cejJrNwqsy3uXv6OR4gUlCeRCaR0p23OceBcGB4/qiok7CjDVJZy
e7JUx8guC8ytUtiiCPMWTkUJjXzX/zvNg+hOKPhTz3effI7mrwKnXJlYUEtTO/Oo0UQ6Ne5/JNHo
dphxjyOGt7dkar6lD7nCJ84iEHmTwI7TpUaVEweqAGAQlVS6EXb+Pu1JMaLXzPFzZ4hENdw9E6FA
tjCtBbNoGG8uK+/3/8SbCC6SgPvCniEMpiZaPKYDCpAlVOQeWk/A6uSe4vD21W7xGaQRWKkXkzcr
76/iiG0m6WoCI3qdeZmcpcXZ8k1DoL9KOrdSpHZVa5PZsIDTPGgiWVnsC/TKyBiBnkBKaU9N3e+L
MwOnzTn0UpNYIvH9zL1kIyIduywgqpo7EY25/hw/Xzs7jUOAZ5vr3QEmNjTJGh9WoUrnHGTu3HCp
KhpS2AGNSJsigETEGrHgWZn7i5NNikFLRa+s1MYwjyMEeAD2VDP1bs/6QLYFBqFIyqIOvXkGPGVk
do4RiPsmkLldiPjqvMltPyMFASDSeKWQ7NzxffST29uO7Bt8eTganipdUr9EG/cJCxT5A27wVNTW
0PgV3C371/KTchJi7i0PgA4vTm/VDV3F2YeWlit/khdEiiCeOobwRiIYzTBmXfBdGCEvpexHHoRY
p5ApT0x5L8+7vZaEBIRa7dmONy93cOKCGKhho/RQxy4IwKKIu9iv6ZrVf8BJmTX08na6f7+bKXA8
InUz4Lqkc1ifJhT6JwmrMJQcpLfNoPhmV9w32XXJaTTsXycbHF5/Szjs5NqQ966hyKRJ7kL0Gpnn
R6IbP2DM9JhyWvRFWvpFfL3/NVFzHHOLg1FZ16gXfeBjlZYe2Iw4JWj9RuWW/Pfn16QFR0QOrup7
tDrOuT/GcRal9piR7xWpsXLo5deFIBPy63c3z5o2iInEuEpeRypKQozzPsydkCFuq+m9Sq3e9Aia
5IioEr9DY19QAWUbL5krUzM5CGz2CTX8U2ij2mr4DBXvAjb0CJZ9wZZsForbK7glINF6sb5OCJjm
y9Ss5jyWR2ZcVhrsjvpwNCZ2PvwFyX4n71LTLdaO9sxBYOCR50BgK+/0XLklnfsM419uo+8U9L/2
UIufK4Q1H9ZliJ6MBNFQ4eh3HTnHjnTKsu4bNa6168/3zsKWQ3RIV8ia5FjPKI59DF/eV04fQDcI
6cZK9JMVci952tMt0tJ9B25qWvRYIvwrZvhKJyTmOR9r9CfdZ0+KcDNNV90PbiWBrcCsalUT2cYi
3YIwpgGyQiXReWRzYqxKu55ogYTUHGBbMDi8ZXIv56KDKXTG195hwDa5U3Hi3/tihFFLiIkxNDIK
fGNiN5HYI8ozFfABF6eeooc7SZg2n7+dvAoMDmKEpE5Qjs7pJivQ9fJ7wR7MItKbWeyjKAtO5T61
WEb3idrSU8xZt4VI4c2hVEFsNBOkfgmjJpuJuYVblFDwxKwiNaXlHOSoRNcMqQHg1+6g9EwIZafO
60joE/pBp/8K4nXidc29fkxqQMg6An9Nl6QMhbvZ33if3VufoC1VqkqNg196r4YwxXnx1n9TcarC
YbsWjpcm84E6CeSsczi35Pfup8tkBX9lP1y5Qpm6Eo3C2JqUgZ/xR0wvbRQAqE+9b7qTRNtHUjHO
pHy6YQ4cFDvopI0cPgqGgrRxcILYy/1I9s/NIQsWlyKKmbHESLKhdL1qnxQErUOoJJ/ffCuLWqZh
B6g/65PVXAlMinCLdTQaKVcYQwm6+TKH0W2xBYaXuPPIbXo0vsKKNQkT1M2ze1pG+GCX9RioIL9p
l3yNR8KOeUOdWfw8K9y2E6eJFvvIU92t1gpea/RPaYNOWIYER2/VbSyZxsE0UAisheWHadLiFTuq
5GlqfBAoY0N/hW3Q47xkEHm5pg7n6SrYhuJOwzpp4LtmUxm8Yg68LVz/ptNGrcjeU/5OFlEzzKeG
eSaJji5vn/tTybtMdg1T5k4U7bmpnFESlWkm35NCTB7ydYpCCvnQWFlbHz+oFdukiG4QGRa8cb03
EFClEInj4xMOrHlWUHNiJ8SFTkAiHN5H2qFPzK6gGN7Xv6DhjrGH9v4NfTJFi9w1puVN/yhKYC0J
TTtJDaKO/Hgb6R9zxN2E/KAxuTnhQlu1wZl81O1LSP1Hh71TdwVfuGm1d6/06wz6lXJJVAk5wy5B
dsmTVQzrWrxnvISNLh0LTpMKkKyHPlKhzxYoMD8i4xCPooxwMq/tQ5mn9gUZWwh/qEnTn6Fq8ccc
RGMA+eT4g8vsfOzjemcH7BuEZ3iWfQzyokKcS4ga4WMIISWoBaupd7KprbwZO5nMRoWgYWePFgH9
lf9wJhfyfvUwmCXjRAbxeSkLpN6ig8FwP1oz2Dk6P9LpWTlidnHWKnNk3yEd/5iUA+UHnDbEG6zx
eyXZPboV3BE4ddTOu2aDCtgZAQHxaHYl810VZatv4yYfs8ZjYPSvsRBgCbiZjhKAPMqiCYadC92U
q32B01TvrC+sq4Lbx2uJ2PP4aMGci3UXeuHcXae/lAoTGXxVQQvPogt8zKwysauOXs23gLAvlqcf
WWl+TRNUOHtVJK7U4XINBOZ/ybSDO89TS4PYT+sI/G8vjQJdsKnAxI59hnECC1+me+E8/Ue5GpIO
/jIJIlZVpz84QydYOp1D9JDhArpTHwMy/Rx4EumqK60ZepXR0S+b1liIVpssyumt1ngqwQ7b1lqU
s8UhRTcGY2YhdGNsbVIr2kktg2tc+8Joaozcti5ZKBleP0/8MSFU/OuyPtFBq751a91Yaa6p5wHH
EeUa6Yjrv0ZiJAIg82j0KLR5Dyxjq++qmO+jE/C4RU43pIvZKNOCST3fn46dDRAsVfnj92jS9kGO
BwUucCZeb/mEKs96MBRzPlB2SLyjhajpuSzBG3bNKCCK0XqMfpQlmD/2cmXgqERn+68+HdWkHvv+
4coYfxtrkwuKc4ypwl4a4eHMhuwdfEHW9Yeigk/JfxVsqCQOVEEVmACt7okcD/K29eUvsqUzUom0
q/k/B7MBJQ075iuHB8xwzODodYySYXupjaJufQfb42MWFR2Tl5n90D8auv+kn4S6C6UlDtjAcLP+
nP6tnyqUStlozQKDR5jYZnUocQgyUVn7yeQLCUQlMRfpe5c1jj6Et+EjKbr8GEU25HoVZuQbyeCb
q4EQJO2lzTc3Nr+GN/jmP8YIBlQUqm1eDHCM4AdLHs5sUewSV78ZXxtO8ZymlPsNW2PuXq4dCsvc
yfd7tUjRzU8x+ffe68WoARghKQAkPe0igIJofYGGWNujbxygHu182hLddxXyWAdh/N324DAjBK9Q
J/sTkFaYSBwlPCwsaELA/fPdtZpihtHbyamlvz6q9LTxOHfxnsUuoEB/ptSjEeswwXsaNFG6zE+z
2ga8kGCkKg+TdB/IHQRpFmTGA0zy+Mgvi1CGe4AN9cXUkALVxEmRf8In7CR5fcMNeUWIDze9BNLj
G3WcHVVGvIFAY5C2Yt4KH0yWWzmySyxro9tTclYW5L0/98P7Hw2f34Pz8nqtvS/h1BJHxs20+Cnj
20m1RnAW8sY5H1pVkaQ6XxynXG1GvJ7CPHgnglhvtTPQqvxvywdX0QBly1EoZYPgm9lIaOleFg33
YT7cD5vmRfa3pMOFumeu8orW+9KdYRiqXcTeg93/nj1YtcUqiF/Ts1rtJVbb4yAz52UzdDlAstXp
fem2H8AWpSUXQ9g7LlEdNHylnJ6oUnTRbBsc+NUZGyWI2Okn92+rPS1wvr8tdqVLhtFG1iifVUh1
mCLYotJgZZF4Z8nl4SonmpV8Dneyeppth0qQO6wuXwE0HhtVzJm2tYfQ2uEcSYlOcb4LMdI3e/z8
hCNF5pVkeDeCVAhd+XzLEXJfxYEDHTiDifbQh4/HLMnXn9RtBHmys6+qQdkMMXo2xRKhtPnnLimz
6r2RHtmQ6sjLH9HPxfoyT65z4uuEBC/xv8DComN7Po/n+wZYbpxRzedfgBro78RKr2DNmHtoIpF3
1VH0uPDKPP9O265hiKFgUY62apoxsACgm0b7fx/usp7myBvsHzlkIsmpbACCU10Fd/XLJKrv7OeP
t+0P7j2/eK8abRsL1LGcc9RmHQqUBBA3DQqRD0F26HDWyJZO27PPNZ6ntn8f3/7/iIdfP2vMEoMm
SU1pgcN0XCdj+lueXFaAlPe7ipaFLzmAnRLacMM6UHUFk1Kcgzgs5Tf9ddWIaUI4N7zF/+4cmIj0
C3Zo7k4N5pEbxfLYnRS5wl08y1JHEvqj9P/SHOEZT5HaHPfzDNCnbYgAwX7uSF6shFsxJg4YLZhd
nwUmyWGgkE3IYfhI7iecFYx/b0cowj4Pi2X1Z/7VV6QaCdCqq5PPpa6WCON1Ieuxyq2wJo+Spvxq
YS/OjQpHwOQPOA3UbHIUohQqmxWAW4ifISUHhhj0BUnBX5Ah28sE1qkhGrGPTzcqUxdmQWxAqdBd
3eugHeTahoPTEsxxre4VmW70X3Q7YoIfWVoTscMN77qIEn9IceUESHB7E6B3E6wFi0T9rBT5utWA
cfOXQR/lDvQkzdJe9IU/oRWa4m/wtfStmSovfB40TQw70ZoIJS514xJHgVMo+q9UrI+DInp6k9I7
EBQH20ZZEx7zrioAi18u5UR33JEwdQYT3ZbUTouiO2wMeFxyVhDGZ1rSLwbig7e3mZSKeMNHau0s
7pWTsvUsZ2jx+InaFWPFQxOW6zwfi6Z8fDxNP6KJAfr3q2KUCd4sFqL3ZdOU3Fe7+ocN6vKaD0z6
GHXOubTx30elH9QTvbn0L01kfvpWI1VcnXIhMnJWKOgxD9K2b6/qtEf8xhPP27zioGwOyE0Eb4oy
N3k0T+TNEVx9sS1nusuoccg5kGqeo4T2XXd4yJbejiVyyotbNKYnoYSaUlz7bskP+t/U25UGroTX
l7lFYGTIWivqD/nx4Kb4MfCd69ML4+Pflj0vSiWIa7zR1cs/fwp5IlA6FxUqdmIKyBhIpDJEaacE
pdfzzBMIAsiFGtCw5vfxh258HemWIQ7XYUgGyLY9hpfKf04nHs9y4avkCHBYYSXOxpagYYzQTlfb
c1kXUwmRA3W1dUHJfPBdPZB4FknY2VZ+wvLW5kY35g4zxyLkYC2WH92hlAjeKXDEnidQAx0rdT2m
12NDsPHdPItiHrkYpf3UadFbvjCbkc6KZp980aZWhuB8nxdY11Av1bKvItmtBSWPGZT0sgg+TQr5
VFbH9/LGQuFwnU8SNQdpPBYf/Sy9Ta3HaM9mc5Vzw0JG7PotBRfHP26Px32xTdLLRiIxJ5ilE/iG
NE1DqktN98nngqp5saVqSTjsE77UpTjcvSNe+Xt9XNviwyPRTdEp4YxzjNdtzP3GEbeaqPYG2z9x
aaWI17iwzebLfwT761boJJrnbnTVZFY0P9GVivLnIVt//20dPiWxqyBV100rqC/kTPA/jR89aGQI
QETqOcaPHLdodWJv/FquKOOQqn/UJvKfK1jD6Z8tjGXALZ8UmBbNvlWpoinxx+G2/Obj1/TBYemS
fPjYl93rUath9hl8v8POcWBeHqvqBMuq+MK24o1RLkvWBEPQ7KwqMo0FYPLIHAaAj76vabvjLfi8
UblDB7/8XcFUFcu/cKUe0tQR+okwVWaUicRMI1jIGl4BfETf3C4dYbXR+UUhePvUxZ0YoxWbdQlZ
Yz5T3UrkNJaZ7oZPsB0VKnRo/hyGl8iTbCho9keO7Rwd9AXf5RBdz31QLzoBJ1m4a+TyDvGU43jr
6uZzrzUDugJLD3qWWdOfiK6SeZg/Y06cA3pbNRexf9nIGdqzrSRUh4ml3f9coFrmfj8UrlkUKZhi
gQq3aW/IVTUexLWEE1aD6ZHMMnkiPvHKWHORyjB4xztelNdkYxTs2N+zoM33LB2Mm5abz6b2yxjq
63U+iJ7APk6AglnyovjOJT452Zu3Wjy8Rc1MI9PBnPZPZWEKqQed99IdV/jNAX73tZ0OvdQk/Jo+
LeUPeI2+2MlNGP5VgE3DoNLL+/z1eO/YZ+phSwzzLFAOc10yCEbvRhf+OEFxTloc+SeDMUJz+7op
nmHmT/3snHzE5tmEV5VJ33IlnS4q/l0siDDQ13FUFcVYkAt6ibe7Pn+dYR+RDlcJJmJjMo4BMZon
sCM5Fc4/Up9ql4CXnjSwbyJNm4h6rlZhRBLEhtkeXlcaWkePUyd5CzKVS4ByyehGQyInLYChb7H7
fm9P+9L3zf/t5hs/m3s1pibbC+1l9GuCczKAUpG+O+fluWoy5q5NDF5yTMZaGloh8qrrUGRdBSff
CMnvLw1siFepErtI0Q6+A0zuvlrUc2ARUKfkjmOH/t2XF6rhc72LvtvGzD4uly0M5w4rG/GCsQB7
SB3NibbacMAx9GBubZVMfkJz5cb3zyr8YpWW76qh8eVpQ7h4ern1/Mi3v0RecnVbs3BFfQgG2X1n
aR97F8INSXgpmpAVD9R5cjNTvKCzNsRTlZVl9cDCXk0B1GjybHFgwQ3nSO1S9wq12pU39aTFp4Bs
9uCmvrntzDgtBYbHDI0jP0LHQjZZsMNh/QYhyNITVK4fKxoNGZCPN7mGI084/jtL4EYLrKRyTI8e
MqyJzegHvw7Incr4ydafPt5SM05HCumdI5MPX2iWXLul6WkNWdCQeUWYuxkTIgOuTI9oEpPdi7e4
ndi9efoCo/rIf5Fo/M+dZIzarzVvp6NGOsPe1NMueNXI5Z0H9bHOtD0q+KNVnpPYRWJ1byQJB2Iv
hyUXoOfrFhzJfWRlgV7cE21d8YsG5BSDxqK7wR9y/w6DkdHJfxukd4iF8dp63W6l7uP152Q/rQbg
FR6wK/rvZ5UfIYf9S5dCCtwBYPCFgui+8cJLwVC25VTlh24e0HwNIAhIFEckNcsZ/QLjLppHginn
P+60a98UAs/IedY4Eolw8zwVED5VaHp2SQjpvrJ/pd7V17FNkeHFV/0btohWgqVjapilPOM5HnXH
r1i4St11aOp+4BT+YHfu601Ln67lvigwKcOHgrfdFgyKc1OqT+/ozENjkOMMyVE1S3SDDjYCdaQi
yeFmHM6Yk7CISyvz88fK3aOgGaLPj4iGoKcwunxwZHQHtE4i3njh8YiDx74gqtA7qkowEsx1pzoc
j5G0ERkswF1SeDm5Uh+bV9nZO5vrfYfViAaI5ar2pkiN4/DfiR0x2Qbk2yD7OXf+5CyeVyTwAYjZ
+D4aE1JgLvkLEd9VkjhHE16EV7yfBiX2KV2aCIPasUpkDPu2IM/zWZbt3j7c0dgxUkT0pXz65f3u
yFIXmJyfnDgvns6RrI7IP+nz3vA0/4WSKeuNJM+0yxuEJlguyBnUb3EPv7EMEaLVItb5/jLMu5B9
zX0E+NuzgqbcX50U12qBAtxlmBNoosUgnd8nuR9PDZf+ZBmWrizV98YQXQHmtAcl7uBaDgG4drAQ
Cl29/Hmg7rITTgtwb+77sVEMZ4lh4vVCBPi74R+Q1d/Iy9E5VFLVhzIei7aMuXcPagHsnfBCt/2z
JpFbUvX9gYI10VlMrALQGXChFai+Bre1xBOOBLjZNG1C9C9GBxYYHzL5tkWif5IAxC7kWw4f90ZJ
0u3Mm5Dvo+/RaNjO0JISqZKMDYCbVkC9EQHO3Wwqgzh/OfurwcfqpxumE7vaLifObxI+oybwnQCn
3IqodgXccrnCImlNLlgLvDEb75WD1TATuslg8YMf0CWHQWJXnn1/RZgftwoFb+MhdEy8jQIbc1Yl
TmpDFBMBWIfnNb6EFEFHH3BvtgggSVTjMy/4d7AsMZwbONq4u3G30OzYbgoizLQvQcl1upFZHTsB
+RJch6jw1IMtp80HF8pb+wtaf9PZpHpldBbUwHp3JFkNgAgKwavDWqpmYZWgs6wBLDJSHZ7xlb3Q
ZtAckN3eb+nfwtva+32ZY7DOCvvjYQWAApgE3qYnbXDuCNrmU1yYGeFLpYx2RDhO0HLFajCCqs8E
x3vWaBUr0nbvrDCUMiMa5lDdndk04VkavfrwQGca+hIpDwYc1cGTP50+df5Cfx/+ohOmrCur9wa1
GCNB5Kf7IYvXNBnehAK1vWN3+e0EPkekKownnyH8hAqXbic4cjeSIZ1trCOmPaiKvwc5EEJ/hQp1
28EazZUZkfNg35yrHPePVElkCqp5nWk7pKMHsYOr2fi7j5CEn+YkXPdSzyK1dKQfZ3qZR/82WsNF
rEFQcwWb67wq96b+xPLhfjaPpwJzOTr4Upc70zplRyNqYCjdsQW6dqFdr2u/a62pLEGKoPf0D3Yp
EkCAw+ZrN5JnahWBcpMQhzu0EXRkA+15AGT5Xcqg2twj+Ezz3Eo0WW/vk3Ra7m4Y6lsPO5NmhtRF
6aOV1Io7aK5ajR4h55MdWBc/a06+iIgEghaHJy+Mb9V09RfatDvgDsRYEBsxSOd/RtDW+/prxZYR
FuYVHqgwQzH5SjAXUzJvwDd9XbSbQCwpMATBm7tbwLxGO4UVf9SHFYB9ROBxO7VvcJP0NOEGrtaB
R9SMOsOtnayNvc9oMDHklBLt5UWVtmTqD4qLZ5LGuBwKEgwUgKaquGcT8eylnsnWFpLLp9hKBRHA
hj1oQ/j5E6QOdaE9foxD6S+zUFmuOwiABUCl355gld5CcwkdmC9Vy6l50/zSQj8SSlFUCHuCIjfd
/XEoHE2sWCPFmFh1f+jDIb6QP5bd9Gym3VNXDkyBrRfAV+ujyR/1iFxNNAShUStwER66A3SY4ghH
e1pugcl4luLFKnRwgEGsS2vTLLTT8GRmDStEndj1CeDJmL0kvKcII1R0aP8O329HuS6SSEXlyKso
kKNI2/+RMWWG0dSBq8fwrYQQtD9y6AlpHcWm3eYqSOBEcpSV7lOLw+t89Kr4oXts6hvNGFHk9g+a
rsp+tSLipsqPvaaW/mAMFmtm7oqVXwB9Fuo2hw8HHLvaNvJzayHmMty1sqMxzLYs93ngHXx+ShGr
EiKW7qpQp1RGJpXfzg06Hxd6owMopyniuoZT33Dtp8DDrPUFcTpOItlQ/k5mPq+atV9QiFq4lP0G
pr/uFKh9tMpIc5miiDKaoROD8l0Pn3p0F9wEzOe8VFMWdE8B1oHSruOCswIr3iByxlSddfI7PIVd
aMqAQ3xX/4/+VQhIYFWBJQVIIZUwaoH0KiGyF+H8ExW9v+VG2qD48f28+RqbGAoQONZr6aTu7v4Q
qcSnscIkXgic1U7fSpKUSXsanogMZVy8dHK7fCMSvT6ip724DCklbG8Gu/KoonZMILhxBpM4Jqvu
5TRIbR1OAuDUFUGH3mE+f2ca951A08tMGCbUgk1vrdLItCq9AmlqMevhcIZg1FH0DrAsDYmwwD1W
6tHtbDnT2IBh8UHXM5r0XZUaK3kfsWleiu45hOV3H6G/vzsWz0AecOtUWf/6qLPk7bnZufXC0xGN
0VKXaMOTQAODdbGYvc15geDvhI6xRuc/+NecV/IqAWaNtefVT7e9wgWj1MxIv8+lId9jf4LNbZvp
hubYMMxH7uCMj3jQUo2wBPw+DQrI+NU3VV/i4dHYVdVV98ePxu26ZLJMsUxHqtiWMNbymj2nuLXS
0nHXqTbmRsHh7NGejUtRQqqeG+kiTP28uwJGtTwmO9D/CwQzT0emd79cfov0z+TtrJ+kysIxF73h
7YLbqfns+m71tLspb0JcOuqfkgJk6K/nmYi8s2NAU9epkGennjDvdHGgOE2oirUpR/2OeJr8A4+I
5sStcjHGkeUVcTxcmfxuXQC8anAUoHGojgErTfsO0fCmpWUcqNpr7mTwqeYJU2APwwvVZn9qYwpY
MjfFCMLh9I+D5HXnvc1uz5OyvmejdReY9cxLiU5YvyOlJDY1lVcR1s43VdVtvbd9YHasySZ+FvBD
ew/kzMFhVNYr1m73KA8enn4NspuiZO1VICgIizlTq7HDEnzqvH12JlpPRmUUVwIcx82SBCZHLhv7
Gk44RrtwGfvsOECLOctHCY2ZKZnXSfMRnNaaSzGOiiIy4V3AJoFd9s+SO+/0KOUE0PYm6/jiWRQO
OTRXxRCsPrQb63Una3EC3cUhLdfEgaupIqEvAeXEjP9fwhCwU4j68aI//OJn66xdDFW3KUkaxllV
oeESuzbFr63SAxtQBBq+1Zxhizj2H8L/iigo/2kRAi9NdHzQ70ewTZYh/fq2QPwNTa0/ppSvtMd2
YvPH2WtgzR3oblSaHyev4EFlEdSUbTApBfwzc4uFRpHQZ3t+vH8fFkJ3vOOEMUfDAr1/eIAZdK9F
E9KwlbmrhglcTxBoX0UoLxReIrSHK/rA31jgKmB916Uc+WmRDCZL9U1hP+BTPjuZnbvgP6zOzsXE
bm2mwHZVibrrhMaMfNf0h8VEGL0wCKsTwTreAqzAYEyg4rjecTzw7Sg/hFtU9xonPvTAQV5kfjEd
CSimkKStcVvvzPIwSPkMryz6xUMY3y9aR6TKHBlWr9Ptr0gXdaZ47fXpS4MTkqyQw0egqghQ5pNz
PFaenv8t1+ZHzmY6UEdpOp3yL1QQqABEDMYhPUgj5u6OoSwupTr+IexJ8hf8MeyBzc8TaswHqWdR
AHf+yBGc9yYCVLhRRYj0E5cmNxLgaaFbXGegnDrTZL0LNkW3HHLYe33ZyzJ8PplMUwcybaq+xWNT
T1UHS83EKSLfyaVQi23amvRpW4HDl/fwftWwW4h53m9nKcB838OtjRAyfNRTBNYHKtY+Lhc8swV2
oSE8yphi/HhSVu97P7K0HT2s+KHG7YYWmTCgvOCtvRTndby0KB3EcUGdlnEDoSxtG2EKiXYAJZbL
uGraP+tQc4pT+9WELziw53tmlv71nn4CxZBtbn2XXVOgyOh1jSFJU5occCDm/seHMAiV8yp16wMj
CbcW1piJ5MhHKxn2r3tIIQlv4fHbWQmNR9Cb7GRQoMRTk4iWsePcH7qfdIwFybSzMa8NY19T9NIZ
rQ+1mV2wrtTBsly3LWieghLUT/EcvLnYRNEA75vvug9TIeBiYuOIz+rxTWBXL8iMTa4mmSGQy4WD
oPFmsBOowrheuJ4jODKSObajSGEfk3v+J28+x4XmHFIoV9N0q/dwyt8RO36B0v9TdwxE1OhWNC2y
acMPdzdHstXhupqk7K4Nk7IeDN+4H5Zv6BtR+8uUpvawqNxqXhUvp8F89VjlBp6sAG5HGaAjlaLN
lsNJH02OAcq62DrxLY2CQRd7bNuJSGZRdpZEhgwQ7lW00xTd1P+t9BngmelHFS8IWzg0dSI6PXci
bO5tKet/TTWD7zepEyiDp7Z9Hs3OHDNKYWNFMaSh2qTCqz0AjdMl8b2BsTwHAjiT3BoBYvfWaFnl
6+nevy5BcRDifzgchS/tjBLuu0qZJRk+MTIusHGLAbxdN3ueUYvdAqRM3BfvKFhwt81qbmixE0BR
ss221tE2+earLBUQz5aY+fTPE8lJu1YY7NnAZ+z676t7n1B9ktNtB8nAS08g89UBfAnHd2KRjfow
nrdxRB6NR4Z/xHTRhYlxXnxmTpVmNT3usjyVlDLCkbkyHw8nXBgsVoYXl+kkUEwJK6Z02stuxUEK
6o0M2dVm+ihGBuKJpgz51GAT3Sh7/8lOciZMG9XuhbiNu9Oc3fVurcryos8Ug5pjOTPKEtFgQN+U
mkWFRJqPG5k7mNu3BxrjApJrDdPTpNZhd9bLin5iQbNxsf2lAqTPleSV8qGGRYupabI23OlFoIZs
KsEG8IMLFAq00MrA2Y1mfjviEjBL9ft5CFmDP1Gc8SM9+oh4QPd4FlNP+JmImpMwVq/gXcZ4WJ8c
cKHkPy+O5ArUoOz5w00c3r6VC1ZN5tb460CW9MFqg9brh3CBblUqXF8xMdjASt/0vNtrKUsnLJf2
8ONcIesS79MtqpeKxDSGsAZd+SEEiHcicd8qrILgmq0kRPyrXDxMUl0Bo4j7TBmBjiPEUcdNA2aC
Q2DO5kIWVpBMT0utu+MPFblmAsX64jiRihvU+EotjMP85N8Rc/AUBkEefkLOhequ1afNBxbmqZ12
yr3mWaXuUYF6CeXo25pwuEJKtRd3fx60V9UDV5Kr3EZjQl+HEPxH4QtQzarzxeWhy9Ha2etC0aqY
xMpEIzrT2jrBuKzEUdfjQ/5c6kaG9P1Hd+3R360nNgthoQwFoWxa1Z8nMLGZvuH558spdkGnIOQz
a8w9cSTny9bIKlzwXJdzxGeyXvF2fR20iygOawGhFmYc081+sBOPW/2XpVxanqRFbzjdsC4nf5kt
daIt1aAxxeO1wBcSf5Si2o6di/9W0v6F0Z0EL6ny2zDE1mUrvdVEdtfm8sT82Oi0nw3xskaB+lx0
HDv8PvyMxhQDYFflPYrfG5yCbHTRibHvbJypmQ8tprtqBvLRceRyN/zl3Nq+5zOAV8fthOCMpZRr
Sf9jq5APE2BluHfzAeTWR+1e227xQRettrPdjgh4IhYei3B2O7vnXSuUQD/zYmTwbK0/SeOmBWnH
axdHHUj4B3Jpb9C/yS16/YAOGOmQveupqMT66Otz/vOnyFeRs8kIn5fRfxHB+Cxi+m9GDON+xH//
j00IqjhE1ATa0ECTfm+b4CpoYmOfbNXJ40DiNz8wouqY22NogmOSetgvWUHsXrLKANKA1Hmme8Ns
k51PPNnfzGMNQQc2HpJrqdvb3AG/aoyfGDIKKiN6FZnVrTL5+s6el9epbz600XXCJ3EfgF0A2WOt
b3JwYXEc4xS4kcvTFmQMgIY1ZsrkvVoGAk/hmAVqRCHyb16N/7vZfGXDwND6gADYSCB0FIYM1c2X
cuUDovsJuDkiaZur19Yyy9d5eyTCxdAsDNVf0IAx3ujBOmn2wxJzO0cbVQHFBepyhRBcOHA1pQmG
GUxiaYY8alj3ZKBsL7LlLd9yexpmDHqlvJz0tLEFn5hWCDS5LXWj3ZUxAD48xbsckpGA705yLgWN
/ayV/A2ma/Q/Q6Xk1t9S/bYJtWOhYqvsVzyVL2E+iYV3sC3s3+ENtb9zHdpB5wydHHEObqveaA5s
qulwkNkxcO8hAs9RsPDu9Yy43cEcmmTwdK91MZe8xIz44N53L+gLdlipxOJcIQ6VDbZof0vzmeI6
78DfruWjDjODVi9UaqV+yn2frHCuNxyKFhScV8iDQ+JtbTTnzg0GcfKx0LjrSfzKo2UMjvVyF98A
u5xDofGef5FWZqCV64k+hbts3l7A12QpGp+O5ic+owgAaR4ur/sn/Bh/4CRQYA/b2LIaZKoWEkmG
Y7QILSAFxwKDUhQJ3JnK0SvtIctdL7jZyg0xCsASmHBxRy3HoTnaXLovzpIsCXkdSllmNrNpTTUr
d/Vq+FYHVdl9BZWj1M7VNLYEaF7IQEWPjJH//RLOWqR52c6nE9D/5zsitag3Tac3GU0aJ7UKS57F
ZiPLAQSdUTxdaxcPNT0Z19OVF+vlh9Z5QyYyfITP8ICQ6ZCsuKDkOJyQ1PdxtC3ix9H0u2yIJdW6
/GNpJws40aDk84ccviI5atsLVnUvnmmpnEh8Qnew/SxJE2/suphRAI8L+J/wYd7Jbz45jA9bVo77
3INmIZAYB4BD8tuEJICjsdubG1wMZzELwhzBgufrW1aeDayhEXHwRxP8mVLjZPI0L4VIK1yviHZj
h/sRDynSQaS8vesEvwRGdZH5p0o2QGl1RyUgYjWAhFkMs2f73+Uo6+9iT0uQTghgZiDQGIW7iPL7
Gm4MSsdqT6HArSgG/5QHadcaTj0qnieOiUMuA1++PP7fa+4WPknj/V6XJj61foFYnWLSE7/CrJNX
tRI99IGyW3W5eq9eEUPf6NXYkHpC4cuABO5S/2YQKL76PuhKL0lhYyZtkJZinPMpZtT/tF88hoQk
N+AKBu0Qie1wQQw1ltiOuqn9zDXNz4lfSQZcH7848yJpu3zq+p6J8K573iwYNJXAkWjwyfXcLI/j
85moUUc1jTgecuc0Z81a0vU4FVD4nsraHx8H91bNjSN6nVPhc/RPbr4x0m9c5RtCH4I0kQo45ggp
P2SdA0WP8o4YyuD5YUxxuKiuSb7Twf501e6CUzF/ox+2l466PEvhDvLMYl/a2jI/ZOmuIeedBvqY
FJVEI/HQBrFR98QBzA2szsTPgdUu1BFypv0fR2vdPdPJec4VRhZLpTd3+JwlXap/E6Wy7I3S/l7w
fWCHJ28nhI7p8TMOdm7qnKIgm1P0yJvX5mWNCFzgvemtB3LFut2G4aO0aY4d0o2pcnixe822Es1S
7tajFYt7xwdW1JH0zlLsYOe9W5vrUOeN/7txa6opGd8Y55rRw8lX9tbOxn0qyj44MVTwiL8Dt8ah
Aplg2ngMtJbgseu8GTWps5kBCfwtao4Hz4hHcdrh0FbgdxLSxF3/T8e646b18s6xEvliz+vc7qO8
FmDpNpNU27Pwmb5XiUoqT3R/BLThTNVxy62SD2AC6ufTfV/YxlFs+BDgot7ibrFKzZWCSqjs6R/7
IMeAvcqHumqS6lHMKyLuvC4aux++PmAYnEkUO+bZqvMBcAJixRQkOaQX06hMoW/802VtpoI1U9LU
EGd9AuYD/9xGGlh20s/ozlVlO/84bEJWwDEmKOw6847nZ5DDTFwOsjxooSJks0HoF7i6OmgZbGW6
Xo2zIrkQPKb49ibobmebl7B/fsllgVixKS2vpRw+9CmTfSBRKViJJFVj+Tz/pK+Gd2qNsbLPwws/
MDaWxiq61cPAFw0T2CEhPVzjlLQT8jXdVfP7Xrv5WJ9BnGIgJIihqAexPUGPb6QRczgU1BbdDXep
8xBb3ZrrHxDRwNgyhIZP5QEEfpaWvNxKgvdcgLjgUPBCxhrtisopSAsGiILF0dtzn2qUa+zApIvz
O2BuBWgZUCg7DukB9aoCf6rnCr7hUHqiJBD8w9LONj5bOvUCVUWYUF7mwxtyvIQNaKpkybxPUYSC
vOaXxQ7oXQCUKgRted0a6dWL9A4RKNfghqV5BECeq6RodcLKJpBztTnPuWxE2RtRBU7BnSv9WQdI
LzdsTjKz1wQ90aGNauE18aYsaBRLQ+P/e5VNmHaZhS0zPl6rSXL6XT4jf0Upi4yOcUfRZrY1ACD3
HbGMjXA5zEYwmdocdEGzvh8PGNrjHC9LtQAIAGkjNRpUgnv4jz6S8NYoVYOow9X3yxSYCajpAicx
URL3FFUalxe/zY40QkkyWHRWX0iR908VjOYBIZh4vTGEjXlt0Xku0JwbSRHBaIAKnggEUkcKItzD
uAAkqFj678jazX3pMJuZzxh1NpVU7YepsSXoO93EUQykwE+Wv/JTd1o8fYcd0+TrGjMhGxi1dNQR
Y0KoruDIZnlWJkxvq/gbj5XlrREUlUE5z6CEWKK/udGwj6futY9oWijzOtGHRrobbU9VH6sQ4BMU
5WDKSlq/jW1bSVb06dZKKGiQdifUFJTaypLTVoUdl3RP29CvxAYgrqeaRb4PGjO+7RI54rMkwnC2
/GLJdUvN9bFqPb7J7Lgd7/gXLF5qoH9F8Xt9jNoWPlqxo/WE/Vs5QnU+8N5YgbEWTjtQpkZuVmR/
ZKYYP8L43SGUDd7M1ZCdrmbZM7FGVcS2xE/m2pTQPVeofmpGRjLrrklMNHxfyAndqJOymV8LIAiX
8rKObrogjBZpcmux14YQXaa3+BG9HJl0qRIZyty9L0l4sYl3IXC1v+aZaFmDKgnWXfOyOe6pJ7Wb
WeLu7kY6QB/LHj89EH7++GuFpDS+yx0pyArqnLjTcbgao5UOJTtA2aBH7VwJYdPNfeSSCcsQLtYl
mBpEdwWeOKcjiKppvdbN6eRNzYQK9Hq+K3xhKeKbnDmOHocS86XPh3ThG+CyYpmS/wMdCiHjRDI1
HK5TCnmm4ha5Q+YCj6yUv2fXSnUlsejPCOwHr4+7I+m/Wn0052o/NOMAZ9YQozuf8P4SGaFABmjD
37s6j4kKUJbm8EBjUPPPKAmnIb8DKaQPuYjwkQGm10WiaaG0A3Uw8YW0hPtdXX+gqAk0MyILkmxE
1iE7j8F0TuDZFAvPuFMJ9d3/xpkD9hHKlrTyG8crx8BRoxSy3YA9ebipRMi9Bf5B0ShYO7PqYLai
p9vyJQhaiT0UyuOuDW5nKWGtoIpkOpU+UG6t3noQy7QdCb/oPFi9GNPSDmOj+tdaB0S/LKc+kfJV
88g//Ub87mdYp8n4u3kPgSRf13wixhDUty/1PihDuU8TYy17xobkbE8rLnRtpwMncneFMXUay+Yx
z2aqhdhJXOsyclREGfcRqLddJ4Sekfft38snQmZYNtkfZLHBwsbaLI9HFCULPfl6IJeuB1d0WiCP
HUtv9lRNgcQlQueayvsTq7NtdJWajbH4WeK3wkExZhuLsiBSek+FF/oCyrTk9F9wDYGiuQ2OwX9l
rrixqZvz+eosNiKFpLzb8olSjyowuqqru9BI8kCeKBhPRsNE60dFygOVKtiq56HVf68tvxRXZ9jJ
GSFA2Zh3q8p4iIgI8m7L/P8NI3IykqgipUm6gdewBM022qrAtvxwR52++MO/43PqQxF6CKwwnjBZ
g8LS/oTIF6Ve4ER8YGq4clc+5y9d2XL08NdSMGt9Ah2VNjOsrxR6PwjStlGlOb7sS4/0NXzmWNxj
J6cZKQCvyvSu/zRR5zUdH1aTrLCSboDNxAS9PjDmKWGx6u3t57BbNqjjlsUzFgsVvjRgf9Wp8IEi
SBUfBCeaOTPrUbEgpImy21A8FVryt0FBdo/mXhMSRhk52UIC+nc2MnG39QV5hGwtIB54tNC8f+tL
vH4hr5V/bh3zXiZMc5hn95OI7v1H0gbrxvX4dOreqQjNwsrTRKI3LKad/hG6o2eK79wXfaD2WhOc
IyOmHFDIGwc9StfM/mTJ3rXH5zFPF1Bm9NzpOkb676Qu+rXFdU+8zSip1FtrA9AwcGTQCx1N4yTV
rl4VQ0S5aIvmklr8gOwsj6O0oca7ALQuIWePAb/69+Tp0dus2RLzMcEdBNl4ordFfzn6kl9oL7W9
czpxlBuSFf31mO5D/iIOD7jtu8O6AbUE+aBmslQdapNvSRnMw2ZCaYGgAR8zZ+x42MCGYRSSYV/F
rQ26R/DcsgY+v6/yZDS07xCF2Nufn5hHu1U8i1mTP69Ps5bMFog3r7fJtPbTfHNLo8/VCGaF/JAA
Y1s4cVeqs09XvJ7SXX5zgZlusvZP0aSlCIEpFZPhEYgU50A8COyQ62AWBRrM3eDgYQHl7ndC9fQm
5F+7aAvh4rdS8G4aHuMgMazxynMvsrHt/f4cBoDuHxaA9D6hDzvqntlPuvNJ24gAyb7sNc/KHwec
aRz/gwWcUNrCrel2swnt8HaysPYTiO6BmOPmaZvzs1HY77+qwDlEOPpCXmItzjZlpx3+l2g9cTU0
1IRdtWLqhU60sXYrnPG3FxykYLq3wM0RBQWkVzaCBHqN8jr2n/lnBS9ij2hLMOUOiTsnKNCF6U9y
TvzkCSmqkP0LDDg66Tq+DbBzhXiMqDoImbCCW31FApXzsdo9K9VDwUljg6ZSQXdte1ARaReXkuJy
x8OEFdZmsLwbDw8I/WtbHrISz1+6+81z8LaOtXCnRQk4ygiacETr8yolla0CU4stVnWMVTARcWEu
cnleaHm+WIuCv7Y9WKLWxXvjyrSEmvFrDcFC2i58XZj6zBIOYfeLY/m4wabdTkmp903mu4OK5G2L
oFh81GDneVUI0qDfCsqGB3hib0CTpxvxCVr0AObKnQzDt9T92892c+HVQTcHWVu8mK335mij1Jn0
ByxuODD9Hz04HM1LKMQsljmtOagfhQ7OMB2hutvRGoAGomLNceQMw4eb/stEklEe5CTSbbih34qL
6arpQObRft1cQ0Do3l8McUppO1T6v3it5oR/ot2VYVe39aFWOrMLvZSUYgKliAj51wCOhkZ4Rrm0
guJ/Akd8r9qK3VH0QGnv6kY/9v2U2YAhxiE/MMi8gxd+oSFRW5YRUFMkAHAHWrA93yCPWcM4m3PF
bRIOp/lJFutCnIJxNNap6LcmCOxyGdimiNdbHL9v6+bSOcfA2cTrqq6tSBo10wewMIHU/3rX7/XW
6TbGR+Ol7LS5oGCozrF117PWiK1mbQnBGjZAo6GspEhoTFofFOrznSuiM1SYjGLSwBLhw4LmG75b
ZGv13p/wbPcoPmhfpiHhFDhNNJyXx5ydTd2vB0UoQ3J4/0+dLBfGgkCGvVLEZBiwvmjcUwmKW3Pm
XM4Yd/C/sPKGXoPWQELgw+rkkfa8ZcCnmpJU14/6dLfnmYqx1Z53dD8dlVE0QmgKZQyQGeQI/Gis
vHpk1En6hYb9Dp8Qj9GMTdhFFZlPRCI0Y2PP50HpPHiNSSUCNhZBrFu6FrjGBqf3EyISYUgoA/SG
yzIPL/kgqhPknsK0KtbSt46i+EX5hpqRljEowlwqo3GBqoNqCl0w7BnnqCkiZHTgKJDPoo2KErgt
mO0IEsTapAllS3yOBQhT8YLdHgmNrbfL6sL8RuAFh6Ek4oRJzbxqfhUTTIkj0nov7psgEOXG7Edr
6nATrd+nFMteh4zApOLgs4uLKy/5bZhESpj1J+Nr5l2049AEwXSeQld6vBMyOOMioqY/Ge3ZjW+e
KmmkukB73LkhpvBirXsAMGvkTtt+h9x+dn4T8DuemgEKFekq8QyMZg1NoZD+/izv0WTWXMq2uaCh
RGPZ1sJDEYVMz3djYT9TSLu7jVbBIErFi6KdwAuHW7S69CsLP6/Tb8Ea3f1Gl0XW5sZsDUP67+av
IjtZ+pp9y6XCZguF3kpaF5QyU+WZ3RqOtco7iDvAToUqg46f2pFu1n2xQzjjnkhPO7eWGd3PdTXu
rIXohi8hb+FFjw0WZIcQWl5kW1bVhvOFsvhPZExu3So3uXnUD2biniH4critooPKGUHDpDB7GO9d
6vTzw1JRf463OkDKxNu0e+7+ZBjDhfAmHKk0OzALUuHgcydk4htVNb5wHuHp0WEnBHvWudos62vy
11XF6Vxw676UfXi6VgGkkgSiNkD5jeuFumgNrUwhnd4LgSXdqyDPU5f7ark/t7WNhe0n7GqESI+S
9m8bmvaRpA0jSxyfepnfpjFxoGHl2frVod2H+eT4pgTB/3aFTyruGORryZHCZxI1L57psht4wQpK
U4GZ0FUMX65koYd7XlwQWZyWO/qtu/8woz8fFn+OqKq3Ej2E45WHT3TATIa2miP+wy40/LhZjbWZ
ghIvVZPPWG2FE+VglS0Vg7i51pqHBHSQAsjR0DFrPhsCNTJshOoZTmtD4i6dmgkP3HRpY5jPiIhN
kIEnNaYJweAK0YsrfUvIjcmhg5BCNipK6pcxYmE6tZl9983KHXhKBSB2/iGiE/r0IOdtPeIp+fKG
vQEc9erc9dDJwcKHruHajO+MNJ1iaDBTON0FyJIrr2uNRdaRa2+7IWc0zPN74xsuT4ohXv0WuvT/
EQhdlY1aaAhfPmi7MhU+NhmH0o/7jd3YpwkAyVWyWGkuoiEf1pafj8e057ZmdBffgem5HpKg9fnn
Xh6Qd+Plfh3OUY1TqJVms6gAan/M5DQAdaH3W37UylzgsY/il0gx50KFwuV4/EZMBXeFrT9zYQg8
niqVVz23pK6nzOetXKtWtuwyojViL74uvLP3sM/oNiWYOlHTJ5xGeQzX2G5WlwsFIIGzs5Cy5Du3
gH+48fPXlInQyhMPmigNgWO2oHWy/C9w3I3dhsT6t5gBaMhZbTUc39bxKBftl1dVKQgIq9tglfGM
PJesqBb8y7UEhPcj5xnKqQjfxea+4rV0lYDOvKLJ+578UX4l3uDELaKizdwFrqQ7TV61CIb2tgUD
HTVA5GTJOP2OcCdV5C3eh7sq6w1VvXijOQsE7dPooCyjdoOS7Ycwf75xEl9v15U69G37l6pYS9QL
a359VWDQELBE8Yv8XzJmcUa/w1n0z6YKlH8yI1pzhsZEaH4t0YDbayEvY18mhZccb0EpUvpWpUxP
NlNtSNaxaw9cfbIx/1X8UySeWcDdEFcnwIxZBY0InJO47TbpRabovZCnx70Aml2SrhmPsN9nHP/R
lvO7cIdbh6jN1NEPfl4bj9ha8iTmnHOac5MTGqIAQfAfci8eF7sTaMkopq29PXOcf0PjFZzAuH1N
t6bm6H0fxO22XJNZsG9uOXN56HyFZG1/bLP1KgH8awr04rGo8KzFsGBY9uqOFvQ1yXFj/vvPw2ee
oDbDDIM+jKlhxRB+iIv0guWJvCQ2O8aipRhCiydCKCdVNi0smfu6CPm6IiIzjSZjY3kDPjnOu6W5
BX9wJH2jUTWN9mLbNcYi+FMd/6kaBIkXc9whrOfKtmqsXXKI8JO57i5zin2rhbjUAEq+9IBTLUjw
HnWemVxCa2mTbLWMzygtnOeqgKA1a8aR1LJcgopS1jP8/3OWDD2k+EZfiPqIbMbaZtrX3VzN1Lk+
dGnpksux65Sm9qvMU6ikcr9Jb7XqikmlN/0mE3x5f/7onEHWex54olc+2yMUgLI4mRFSegZ/qNjK
GRcNdlEU/KMP3XIxfJ+exu/3A8yKTuquB2SLtFpVwXri0y9hcDC3JjU6LASV5SXNTTttNU40Xxc5
nEbECGROCu1n8nIGpleVC+CaFMgDkz+7IF/LLEjJaYzpSX1lVYklwQL/nQ3QdHogiD+JAidW6Ijr
NYVe4rknR8lmramGKAICm+t/yUZ/yy/Krfb33zHG8J7810S01G+RZh9ftGLggM6lKrX9HEYNVMwd
APwWfX9+VZ466nOds9N6rQ8DSVc6fhIEUj+C0PbMLqWsjIVdOfcmyZx4e4HHxozm9YVAAIEZni2k
hYeCIdbPkammcS2YvlpVYihno2IRtsUOkwj9vpmBIzhxPiAXl62SGuJjJvkPMToAVfsxy9W0DU40
RXrR24yULvB3W3FYvqSgRKQffz3tJkTbbQxzXkXq+fAQluKpw5CMXQCCIsxEZtEL66RZF3ZxsGLB
El3psw/I2otvzpuwTnHEgqeUxbQrodmRY1puToGd1s8Ea6YfO2zwpCLvlwHFj5NJDZdX4iA1fDFw
iP8ok+ACVKo1eUTytlugO0h6D4v44MrgEXlaGStl3PdZdJo8UBuqPIGzAJMdLGgOtGOgFW3nXjgp
q0G8CFrjq4bEXwfNF43eKkGrcpIMvaY4eTl8t+91VfAVo61NAHC6jt7kpcu4GDXcQp6R+g2U2zL+
gH41Xj4QM1yP/3ckThayhXGrby4wHd3EveN8fgvtJcxxh2EKxVaN68I6JU3R7G4M6a6zU7VXwK6F
/ycTzIYXAp74WrPecpDoK8jUqCciQha5TgGI+s48ptw6LrLKPUurBPWHt+x8kmq6rTCL0wBfEsJB
Bqa0nIEDg7b0wxO6GVumSUdscVxfKK3dGP5XOOp9m4R+2EjeRyPIBcbO7bWvIQMa3/3r39yFtJOr
lkLKnaXfrDO71IeA4oAyjU5nIlGh7K3US8xRczf+XLEmYOGcbsXxFNeqL7odympiotuxLjibLLcE
NqHtHhEvo1NNVaiN1rzpvJw+XpZQ4lOb628thJBVKSZo3lcdbObRZzFeZDGZ5LszuuVvecBgCa5V
/tRuxf2/J/OH5YMYdMFGOWMphNccTkk2S/cHdG+PeCZO1XaJxZhjf7A4h6aAxoD+aygOdJFlO0nJ
HriHdgODa5e34klWuaDi20tsEq3pO0CbZ/jvlASMRXj2/vFTsWoB+i7QF5A60CTrjx5h3O5dw1Ce
4V76IH0jvtHdHSwvXBVvau2JDdq6FvmKaUa6ZmAheWEweVo/HGSufOoEYH7fQkNsnpEVv3Sug3VL
pb1w/1E6p+jr8tRxutGGfZrxPA7+p4bHmdL1WdkRS0EjmM+n/l7xpaNHh9W+wqx1HxRJCrC/ZwY5
baCFgXSBVS5ygq/i0seONfHtk/XQVoLfkY8CJEogOuFH/v7CelJwYtZfGrSztNoREP8DOy27Q+Ri
26+Mk36sa+toNb2S7OAoxDProC2oO0Dvo6xxGBgTXjhwljDy320SnsQDRHQzw9VurDp7fy/Gc0K3
c1raAXUHKfbWRNZ2JIeLxONU3+YGAONdVhNEASD1vvPcSvu8FlS4/k4MYLgVpeZQ9nzASkCHKdMf
ZnYdgpEALyQO4BrJf9NOeUyL+GH5Ku6S0J7+LisyFhFISMnEOGc0iyF83YeRfyIfmW4PeckYABz3
+WnxiqX3rShVeD2nRBUtvjfrUnq2E5a83g8phgWG6a8YgnzuKCkunXRBemQXFcMWjAT41n4K48Ce
WBPfQzu6g2wASKZneN+TSx0IoluBj8bMn9XC5SdVE8DQdSKIA9606h/bmArQIxGZO1fXgEAoFbT+
gss8eLee6DW9g7Y9R1C6etN6ziFuVDZK5aAmBrHQDlI5tLfvJuRibieikjEw5z+27PIvpE9GtG0Q
oTcZ3jkp/uiLREil/B4DVvJteWYgGB3xVOOS/ab5DuQ8kUS+Kd7tDdYB/7ItYC4NIT3UTzoLd2Wl
XV+3lA3AJB2gUyKGWaHaWzf+fh+zHypU6tdkOTr7mCN7UPmvZd5xduD6B12odQplAoSrjv1X4Iz2
oBHiVRRlSZjC6+NV6wZ/rztqtJn8tArCEyQDwLOsAZObcHJ53oIwsS3pBNJv+IURYEznQVq67hY/
7XpiYQNvvpAk2Jp1IBpUZ3RgfjrGiAffeuGT+yr8Yyjy+eLORaxX7iwC5W3rNbuivti9/Ih3fM1k
yc31qeV5WHaiXx5XyOxXXRRcu15HiBh8fd9lbHoCDbBs1qYxGfzwCEajtwE0/Z5ZcHl5NP1mRnvU
skUjxnFXXGnQVz7YO64eR+gxUf0xGe24H8Anv+XfKNGXLgelS95VKWeflIbiC5Tbi/8Srx3LRtPG
RxH11fpU0irqa9iFSI1GnCN9w31ukJiTJg/P5tDOjUDbyVdp0mT3dGDWFfUZKZSjNC69nWkqmKgg
td86cvHaNyrHAyj3m3vgQHr6VS5zh/hXSR6Sp2Io5qeWkEcSe+BoSwMz9Phmp4KB6zc0STBkKBZT
+19v+ltWyCUlT6oFhuqy+zLdjDELHwDWvsGA5Tpz9fJK0CeLtFajHwRkO6kFUGFj9Cxb4p1QwIz3
kQAZj6YhwALv7aZMyOZ5rVZhX0TdyE2cm4hZ3etE9cPrwBhNn1Zl3rInkeg3gD1dtWic7oGN9jwD
5IUmbpB9VAQZg+YX2Sn40ah33vOyPLsYpe2+8fR+vjQKXtFg8qfEHJV8WCNPEWSE3gLlK6CvqAQQ
rczVdqCXwpayfzwAGB1428ByptMsgARj92Jhy61VZQjkZUiIoXiw7sucWOnqOe7chWrrpNtZkvEm
E8QpPCluaEidghABMTdU4XtLRqBHX4eZ91qnez7Gbm4kIw++vj1B5rDxSBawcwHQ3QXt11V13UcE
WAeIoSYRSTxHoVCvFB6Dp1DYGJ7AlHYH6fNemZmqwKbYvO0LbeimgTMxzNy0Aedi+bXZ6ikraPGZ
yU2ZyU3JfthCucY0efKvnlIwwtjuSD+yyrcnGp5qbhwPrAdZu9ZGZRzvg84NbHen849toNRvBh9L
5g4AK8nHdrG4wD6DGS/xp6uMONPUp3WlpdqQP2m+y/a2krxjsXx0xt/NvS8n3Uav/fHsAtZZ0MLP
0EdWRDzORiq2oXjxDNKD6VxWQjiFY8JNneC7nRV3CzWFcSoo8VE1Wl9VunzMVXaUg99RmvfkO4Wv
R4uPnSk6g2QMLr8n/+8vYkKFeZNDzbFn4iwGHNNk8mGFaPSIcHJe90bFG6FcPYEI+jArBhLnGd1n
BppyGagBKFrGHxdXWOyp1nRFhYyS8X4avYTNaObfFXwrhBTmcIXpicL8eF1YfYWjIpVZegFi/zaE
CNIMq61FRP5wVs78UR4/HdZAQk0WdMX93I18jWnLDvFRANPW+1sWyyAXLCCgVCacs6iXfsIOb7EE
eEwLngengQ0CWs8YdIBXFIPSNm5T/ix7Fg9Qkf35gHCb8VwDJhYOYMkBOKwi0/EyAaqPbI0pcvk6
NUFtGGYjCcC1H0w5PfQIIB9XezZVSTErmn/1nrhqzx+dN2ev1YRoUzWPQyhlNjw564JG+j4LJScV
RCe6sklPhJlc0zA5pWqvx2VG7E9cah+uimQ0cu2os24qHNP7UcCs3R5h3DyYYxOXufDp65BtGFY2
y86k8Ry5x+2VYSMhUsX27CBOS2FhxCFwdEG0ErjAAoOVNqxIOLzSuY0XfHVzGT9bYqkQzynEgCfI
Kqpoek5rrzMy7RHd0cRMPRXwDGZa1L5FBqQwvEQ5WsLHmJe1RjI7gtTMZXOvc6sVO7VAjfhNBPx3
6O3XncGG6EdzbK7/cOf6L79uocOTBvSSC1WxMBptspOqj4ryU0T2dw+yGEGl2QgYpeuTsYeb3eKl
9dVqHTDoyEsd85xZMwQmbZ8M8FdkRJ/ZHDTMVJXYc1KUm4ExT1rW+Chm6RyjKGa5xp9m47zO1saT
QDiY9l+d6j0xKlicOkv0qllX09ZG75jrdKksxaxUIfv80GOzsqge2Kc4w4SA/dCd6hkh4Ya0h0cy
2H6oDryRn6dRcl6aplzlKf4DViP4c8Tgo/e9MpLQtucdyROu3B3DNbIEoLulEFpb5VqifIH0iPT9
ioPKDQDeKO/J9VW+3x6Wv0nvx1o18zZiXTxnCfGiJCbBGVafK87OMYASPK/esTqPusiQBojdVUHx
p5R5wngFc1sODq/6pPcZLT4eaeGw8cxJFpp1hNYuDYAjG0C5B1VfLKI4zi0y/6/FGe3dplxB6bSP
HvN5O7nP7sFadYmtYIU2MfVlFQz3IhhlH7G8oD21hhf45O4PCRrd454s9MZhM2y7E4bvyhf2mKGQ
f5d3DxtRQ/wuWvIeNyNcl+Ss0kI6dxI/uu+B5bizNWGMgvWKVHAzNCdNLlEph+vGRY44n+dDlfXc
0WZl2wvYwaT9CnnxQ58ekQg24qmte+9YlD7YUZ7++IZDi+CSw88xh6VGzLpYXGVSZa+/FOcC/YSo
sh90Rqve5zPqhvxrreS3z7wD5ACkfWifZpWv7RNkaMWh8/sbpTZL4+dD2w6Nbwq0A3oxXSajCcjG
o9XgTQxYxjY9eiEgMi40oEekRPaPgzjHxfNoIoJ2UlADthkLnTLVSbikuGEFwt/O9A+wXQdJOkQA
9ncq/r6O1vri7UYQTNPXDlynuPD3zixat/MyObYBa+iyxx6NioIdiRynMW8NKNQKR6dMXoxd77oK
W640uvZ4al4gZkdw9f3MHhKvUCyfptPcO6EYdrSHFwXd+yIbwnDHifftZ/6bPjA17n82u9NkquIf
9VmYx6G6M6vpQ0t8KP6pB38iMI/u3cZmeLEeDjXCYF6h8ly3rx+4Ki/wfttfFS0CD6GI0V9aYTWd
+Q4EvmozqvS615V5QWfvhWyUfVqXRpUsReMJGRodbl2C+dYdUvyvFbDO/M4KSMdpckKFooDulBil
ZN9oBF2BPPPHbtlnbJetnjTJTcqi38Pes/anD6vk7sgZHZL7Y5gyRxPGXpUin7NB5VV4F0zxyrkm
V3c4A+tEc7oSFLDzMmfJAOJMmRztr81sWjr2An6l8xUWiMnIH1c6P2+/vFn7aTaq61joz9DiReiQ
E+yrhrOdJtuRVLw1pEqnG5noumT2c3tUT5s/Atn1Gqc4qwCpLWp62y+T3+4jbmOwtj+RD424onkG
SiPS7nnLhUqmZmWE4Eplb6DfbDHNmhJiuvVU7P3mgoeUwOOF6x6Lc0DjGIPdHVZxP7YZBPeGoSJk
0mrkpNGkujevl4H+fsptBSx0JywNY9v+xcytYpWLaBBpJBJc9KrS1yQs3xZ96C5EisAN2MdnyFD1
PgJkRJT/c9VlNBt2cZM50EXUZA2edawfGhfFS1X8MjNBTFd9P/00wOITmCBORGvlpSXpp57P3nyj
yyNhg33fpg36Bttlm1xm1n4w6oG5KSmCGJ2PljTun4tpzBdsG0TA7XmBQS5PKSHyjO6q+4jGPvCy
azGiY/CNSGDNzkgROawFJ5qR5Jez/TSnjsAonuO8gziPUx4dkI7gxEC33PftqVzldlNyq4oAZ0EG
oXcq5vuO5znXK/z/Y42SFb1cPO9xWEAB+z5dDNULyQRF3X4EJM07ezyrxa4g2vMxgwHLe5huFq/G
5cKqYCGxq3dHlTpm51IDp28YlEIw88EH8ppC20kYIgsA1tCuGhDUGIDzgsgJZneEftPCF1/+U14M
a1+ZJTTlHifpXO7iGJbkhA08wnx7FCNudXNuEV+kODMs8qWB4ga+BPal+JOVCBDuLoZe//yYHPs4
xiM90JqAucUYHogpeemQXjUrn3wLud2LPsgQ0UKvORLKlIE/FJYIc7XikQ5mTlaXQ23sC5AkXIhr
sXvOIB0zLz0WPTDDQlmOu7Uee6qbRVwECSl7N/2UAOJA7a6cvTBHP8ZdVhKf/DcW7GOUfyQ3jV66
1sifvVTP3+15hBS8cjGGcHJCYtgn8BF/UzuPH+nYC2gIkt8MDQWkA5d6A9bN3jFy4pCKHmxEdW5u
wcUZx5HzojQFAi+d4szfo+3TIMqIng3hspAr+nY/SzwCc8T0yaQdNSFfVPHtUeYb/E9Bzph07uhj
QGy1/lmLa7UjGqkhOU9PoDP6BVnVLkWW6B6g4vyx6ROaCRKDKN4L2Tcaovv5//f6qkDbp8CfXuZf
hYUmJACg14DPDrjq0nDSBMkeevxr/6ejrRSpZB42pDGvf+ZgDRA5MUl4kyIDXjIjtFaGpNVk0bXK
bdNUSMY0TT2Lk/P0/GXpGCPt47mjRZIKuBJEwYOu6Q3Z4Js71NFu5JDeAek7MvQbytqt0FNFDZ5i
fQnDMQUhkwR+QaCYzcA8chYBnlB/fq7O9q8wi5zmpxUU/5kGw4YkNxDhAoIC380K03f8mznTiF7N
tnhLDfjXZZ+yPpHWCIKA/6BdFstpWGf6f5KjwAg7bW80OAaGSZWnZuzFk8YBIijzay1HEwD2bz7+
KAXgOrXsSzHorCabXKCpyNbyMhNUX3iH3TEvtlCuI94bnIMEtIZqtjjdOTfRxsAMQ98S0jbshk73
FUzPV3KTmS7zZqcTu3evqmGFwTKs9RqXe0ObRkm5aVatzYtCqN2lNjnxkZ8yb4j+sGZinTIBlxeE
oezeWSwWjIy1zeNJgBQCpiv0IahEAe3AkHd0VGGuj6XXrzgcyQCnGtW44VqmTtO2KHAHL41SukxR
QKYXGLCyLIfNjcMOTlVk3sTW0nyvqtWNGEsXxajoDsX7ksclWMVe2ZTP6PLmr7guHrjSS+EAgtiL
OD36MLL3K4BNZvV2pkmVcTHuz+eVQyZ0dP4IVKu/E6AW0UchUJY3DVwZWBfQmmGTg7vQwtPwpD+M
nD0mdGwPr/gJbA4jr8+HaK7mo061lW99sB9D0NVYQAZmpW30izbGEyzBRPQVY4BzhblydNEcYQQI
sQmVUIE8ZdMgk8cAWW2gVsyww4pgsAw6KMlecGs6mFq3yf+kxu44OGcNIglFxIidbWIbg2+ox6jn
THHQ5FfyunjqSYvBxlEd66R12hqJPja++Iv4KI2lXlBHj9Xig43fD97xu25oe+ptZATKmGhST2Wb
25wDpWLnhy1TnGy/HQhArjlQImBPArtKbrdjSvwgsc5AtiXO/oB1tIm3acS38cFLQ1Kw+Sn6+ay5
4cCzcOLj6nhfGIdV+1UTeVrOmUpKW5i4/wcanfgqSDjsC8TsXzrevdOykg7Ma/+ikT7yhiTJmCpQ
7QFKrlSdWlsyiWNnuaSrV45GdQkaBeEgKhxmHOHy3/IHccC2gBh5GCRy4ZXKW4/TzSYTNPwwlsGY
zk4aphn7fV4jRX1ccefExRMe8eUCRnSMiV6dr1BbnmR97OmU6LCmDIxlP/BG3nTG3IR2GYOKi8vO
HO6aJdOuo2vGol1Qc34v9vTcj1BDl20A1F3+yAUW208R6cnFx3dP1xtCJC1O4vD+Rw98H+g5DlU3
zMEsqDlgM96Vvu6ySNLepDaqOT9V3LQc7uULRkLz+vgPq9clEg2i4LFKKbN+ZXLtB+xsfPVQyTgz
9CxK0lMFc8zBC4cgS+zLge08rDP5AoSmHR04OiVW3iN29Lxh9nKMSx0yvLAfgxU3dYmh2gmo8iJL
cJXG8Js5F6enszCO33BV3cHaJXxo0Vkni9aeLDwvSkiNdSkzFxHHyw/v+5nJD69jCbddWn5Xzfhv
JR/A0pPp8rEdh/zb58j5OV7PfipnNZ6wK5gXZfF5HWNM1rYpgsczLzgmbPn+2gRIQKDKCIliHfE4
7nW9b05dIsK6WYGsBldNIgqWGsCYb3unROmOL6gP6yoFKROSizEp2dmh8YBJ2np7+P5JCN2/sQcf
jJc5+t6n3YEp7OyaruWlw85StDuTcYjaI8pHvcMT8wWUqw49qd2yXNUsg5Kamx8+Rai5BKus6aR9
NR2RzLftpdexMPzMiWYxaa6w7oeh0YkZMkF61h1C3UYpks79Siez8klaKwctZDJgZRtioTS+X+G0
PRfS3rJHDNpUNWeyQx4MdTOuGHK3iZZbMbmKwSJtBmzRvYj2dKJDFfGrS1ffF8eA8Sq/2hRLJ48G
bmDvXfGCC7IV/rfYzNBswjgJyYUeJrMw3E5kSuLdV1oM4d8QEBX3oqx0kgvHw8dVm42ZH3i3SSHP
92cC4wt17NdzilD9FPDzfTQy0U5UR/c/ResF3PO2LIwB101aYnNKctxGswz3lrx/PcwqqwCKwIKL
/MpQWLQNIRfxEGkviZXvqo/w01JzNlRKy2KX//vtC73fG86O9hvtUVjXS+xKSdanfnnYMKM7NCJq
Nf6WZJyWPz52y9tc8DlcwIlgzCy2mbwDRc7DJVrhm/0/0CKZGKbmgNjcdJT9VvDFooP6jji1E8Rz
h+6xFxr8AxoKzx9oEboKC8KzcqjHDzJEqcWmP7YPoJU86My8elxeBenqZrWu+LNXVSNyugKKzWtA
+DbaLVWexMVs4xGAi0NNYwd7AzxrS3MlWe6Jhr661/BqXtHH1dGKZiwyDywXofEy1MxHI68sekFu
PkW5hjotOIUSI/5GkecqaOLsuvppY/HzOOGlDkb89d1b/3SSEBjnQ32EW+RP22EZjrtf2Gq1QBbr
eKlHRneKpkQBMHi6SzVJtLYVBpsIszRugfgwIJ2fJN+0Xpjlt9JDNDleZRjXMB8+G+N3C3R/m4Ub
q8Pqo3mE0na7BqVGLa9xsHI5o9FieYkqxBkXjRTkHE0q2E9Wbi9weyr/QIP5NqTgQqg/tcHicEVD
FDHqypmoqSiEt/gEWeXqFfLF/W+qPASuZJbYUgXUHIvSlGcCDrEyA7cEt2kOnmqrn6C7fZVoO/fS
6SGcBVmOJPvc3MQYiJzTFYPwAII/XrJDXW/iRVnG5Ywb0hgYDybaUfqgHMKHB4NyHphgBQ0elGLj
uTRpjJZ8CpVjYLmwY0i70FaiTDYVZonX4bd5IMUDtAf+mClLNaB5qmrqXMor86mglCLuhQgPErUG
JWMfeU18qmSL0QB7ImyL70HvU37jrP0GsppAcZklydeXVPXL8u/ARcZPf0JOjmv+kEVcerOrlWRY
E4hMKuyrf7+3pYHCXUZioQITQWt3cY52+2vkFadTxn9SMVJbEqE4nb4uIoUcuCn1iD93ZxTfUjKA
I7pBdwMvbxXo2STRZn8JbqL6iUJl7vzXdch/rMfEAIrRJPBLxrSaaxlhmDBgtD1D6LNF6WcuW9It
Gyi1IUuo27yLe+K+l2nr/yRAjrlhRqsmHawfWVGudkkncJ0HlDaYAhMjgWatcdysYemvpu5r5Clx
p006SSRiKa3ptz/sQ40MunsbPg/hO3RHLyYM8zneuz++HlD72v5I94+xUxYTmOHSNt5rd42Pic/J
zTXN+UgPvq7CaON7NSeq6gKj7MhEfeuGWJtsbJtz1BjhBgQ/PBsYWWr1LXmeY88UVHAc3ztR5Jka
VGoUmpBTxncqcOALXkWj+TDZ1ZwwAWIlzvPDlqbjj4JvEg8V617C51kMOsyW9MUqTi7B910TRQEp
Np0/JLiz/dbwVhQB5N7nsndP0gah4HIw98buKOOUR1H6Bq6FKvW6B9jGHxF5mHbMBkGWhs/tK9n8
3uGEIOUdHjI+UvbH4qwPvLWS5MkL2dar0lH2JWONC2zLK4TkstHRIE8X9j220IJQ5cmAFqhFDb+i
ZQNehbjh11LmGLjuaw9BYNw20IHVmW4IvxO4JzA2kVwlcEF/d7Hc79GJ4t631PxvNFlPkIlxt0BF
GkZ6Tg385RilIB681EmRJpZ91l+axBOJwKMln7To4cVjHdoJPb+KfZrTuLwgN02tvXLczRIEqFUx
/aj9jpRUFGJYrKabWlOwwdrPtPkzjdZAdPJqr0VegoyXgUlkqDubigc/aiaO6jpLcqBKqgeL0rk6
zOm6uTCNuBME1mtg8AES7MwEP0H97Ju5eph+cJfXlp3XRq21NQm1vcWYeMBYjCTlDNJWAZ1smSI8
fL1gMMCMNEVyoSqHfBihjqES+Ud6YeZPx3VkKoCM6XmlskPn2HedsNZr9dp5do8XBnKV8atVSRcZ
9aDaLOsP8AfctqD1OinOehbQK8vMqSJbwKhh3WASF99y0aKVJ+uVWWCOF0fXOCgtuvETss0OsNkL
bR72RKDZKCECfaDmsJp+hP2aLsVgn0lXOWGM5yijdetmRWDI04l6P+dDP4tHXpjr3CKXGG8rSWjP
5THz2xscQoPuU7pFH7vKEvzDT7Whm56Fh4uGttJ08R7wSRS2YAYvO2/mVxWHsxRtPDoULxTDGdp4
R3ADNB791ti2jdkXDumvQNyGsEWffcTqwu7caslvXHOG/pdCIKOtktQjp3hyDfsWbZgfF2btb/1w
Uy2b1ifggbZjD0ggUC5SAIct4NPj/sb4sFmomr5WoDOse9fIV2BQvlLMsSeNoy85vJB3PvycfGOt
w5Pw4INsb+SQqJCJBQiaJYz80fUq9mP/YgVO9BZxs7Dnm9W/yDrdt7yvGFS3H2ey1yCFX7mFZNnN
Iqo6kvaf6Z7fp904/ilkupU6NyxCMp/XF7cXzT6GVJsInDC4vsaH2O49HY8ORGsQcOBMe43kuWoy
mCv8Ax/ZQMBmKFMhPcFqm0Aa78mkUtwNXl5UC4PQhRL5eCnfsh9CLcaGGKa/P2KbJvSTH2xut39o
OeMv5VVAM0vLCASYEfPehKT4KdswK7B0TFG+/D6eggnj0Wb5AE9vXNxx+i90DmgfHClYxRbP08fH
lW9+nJs02LLahnkGP5x560VpRGQATPthJbSFcYeull2gQSWaBEgNga14FgM/yx708gi2waYmiW/a
bGZoTSv9+JEsTYBNqsf7qgYyKDm0BbI6reF5O9a9nkgU1c9YIdXQXSxGSIxzdoXrZf//EXHu2P+K
69kX4TPfMw8PcaEqD0svQzBSSNIJBPf8STa3oN6ZwuKYGkYv73zTJNXBBdM2ZBlXABRsOE1eawwE
Ia1UmytjaDinDBy5ipnYtrWrVteYne47v6mqgWXRGacMG4t7oKPLoNoT3Ba29n3u/eKeJZlfOhzg
R5RD7JZV7MHqvMbnW2psri3Bp3wbhPT0NsLLQmFu6nLUK9Lvyygf0dWbA/0Wfz0yQGVhl5QF3JNN
UQC649uiursZr+dz95pwq7i6jIE/xIcJih8A3+m5/r6k5RiArosB1IhP4U/EjvENk7M62zYMVt0l
glGl94UFVvdvlpF/VrrtnvX/dN+mstoumRF3/zp26fDBqChF24zn9yhLGeq6BoXiuIAGn+ZspIAp
OmlNj6q7A1aictmsurmTprqQiBz4YgMj11LINe3QFw/rige++9X7EETUgUWV1s5rksMEzurw0u1r
tIymxaVafVZ4MuXWQTB86HrOXwYKcUfDP8E8/HGF1Ds/fmq2ZOWyU5El0ocNFh0Y+1dpEe2oMv3c
IBvxhW9fCA4aYsDbBVV0tax3Du51B0m3E+p8tEsuFZAO5OUMnV7Qf401ix/fsV4jNNb8MrDXXS5A
9MGvTs5FVKAfm2Uwas/sTSISOXVlEsXGNWI6H+qBUrkmdYjuM1ztd/tqt7mS23evOHN3GcOcjZgP
QPwZ+po+Osj/XGxnZkfPQ46DuPaZWj82fda8lvJCVP01jzb1AlvUxfEwf5ucALEZbmDJDIy0CdSq
t6+WBOwSSk2TY0yl4YnOpucfzPlqRd9UkoQWInpcuaqqfFIWI4Qkn6P6O49lXPu4GqUfrp81MbXH
077ywom33arnb/cf0lDM/DmWu55RSpswA90gMj7DaV375ca0W1hS+2TW0kbQDY8BTUyQwXV5ooYi
cHBXXjhZMDkzTDTZZlAHY5Fd745kozA1fXemnzsnZJeIqPXrqjAY3wnxufVMH3acp15h8HC7WrIE
zxERidWkVwLJDqI8+1Yvtu99vOuvSIbzRBdAtTlZL7TzDoACbkMMV4E2b0p8bZSVvbL8n1TO0sY5
YsSe408p7dGYY9H36V+oUNqL/77L8vm+Jr99WX0T+ajKQWs2bzAEtifnRq83/jh2d2A5l784WC07
Sqoc1NO9BF9+h0IiRo+4JeGsR3JbfTVP+wefLwHxwLQTZklWO2J3MXVIMQEOz3mgMUytQmAEx14Q
m0nAGJEShovRZEnA+dcEC26+yICfrd7O7g1tRKvBWa2MwGaRIRnPHh7Baz/M/9RR38D5VTtsX5v8
jofLZt2K9rgb+EfEJKq3V6WvjEaNxXXa5HtlSIqkBfnP1+1eornBsqeX1gQWmF+tJxPLQ3cdJILY
yyRdh5lYRkXbX5Fy0E2cwskJlW6/m5YviBWSO2vHTIvHYOL1cD+lJzvpuEhMx94AfQ11RLVdFh+6
22agdrdLTNWJhtTuQkPIp1QhKSppq5WD99AFUD78XKNP2uRZytNWbAUdGzVeegJ1Wkdi27E8CAKi
iIJwPHvZ0tPDbFNJe8ic1AhdcWQviSInnhL+0jbjDIyNrgIP47sM+C6f5q/xwIM42rCXjrvdDhsr
wOCbtQgJVtuAYu7qND4Jhd4y4LCTZCQKkbN45ZWl6UClr+3NTeRCTJf4PaeFyyCaMlAkgOGnAuzl
SOooNLU3a7CTtJUWme8SaT40JaIr67XNrcDtr+7W5Hr2bofUS+U6SLiV7C/oZsNta7sfeYzasvDA
avh0uQRc2Ui+IjcbILZxoN1hKM4VQKNXkMntvCqIE8/SDAXHelRQPFLEDs/2fn6rdU8FXXXkG7oF
vU5ql29WoS8XRvkXR58o9iPWujNFnyoB8dzHH1R3lo8sd/aLbfOnsGcIqz664ZjEjqcajytaitru
GZher2PMV2LNCcYJC0fJa/52EKwyzzaPP9hQW/HZ2t5IQJSwsuqwE6M7+j4GSGqiTjarlR2dlABq
Eq6a4zGxaIqjuXmnGIYoiW7bzyXwtNxi7udoUL7MUqIReg/r2txY3TUK0JglZH2Qfg3tGPnoMfdy
4JajnGtzJO4u6a0um+2efMDbPI+qTpKmIJfeX2WY9JT+RHlA1irGssILqdh86JOY0QP5+fDmAY6R
CHdcjQqfxIJojRQZ+5ra1Ug0voeOZJtDAD5M1STabdUj8MxIo5kD3Oks84bghkogZLbDJMlCP5Ij
ab1RlqgdPfDIdWwrVjIT+z5z6pRnJhANLdB0WnXN5WXnZuvwR1ZEf4lr+mtiUzr7MzRvzuk6UMM0
D+q/5lK58BrgpQnAz7bA0D8CvlaQCUZhGUgNWZ5AkZI81xPZAkYEhO1Yekkp1WU/YMvSUCJspj8o
KkibLE2yATqNWw0s0A0si5SGn+5BKZmAddp7mU7NoeRg/+Ff4FzGQC/YAb8NkCDhgfCEfMLKe8EV
Xuur9Rw3URJt8OYE62ssmzEiLuWi9hoYhzs/hgvTw97C66W67qM/cUfCO5BTvCUySzxNYNPAlyLT
V2J1/CfgoPqyuaN+3nR1uw/llNHRzjW8jxvS1eJCp0Ywu4IvnWNtXznFxGfMH+E8bE2W2zr0Bvk2
hq2cfoM7rgNezSiRcK77S3dfx9J+3x7MK9HxZ6zwPxIyelsHCwkQIwk/NpnvuEda79x1LjRCgdQ2
DPTQtdyIrAq75Ro+SeE2oEu4SaQMZKhnF2nw7tgdRTfeW5xfp/FkKUxYXyp1P7CgySg7SvV78n/n
ukN5gvzk+ckT1p9JwpgajyKsBDsDMexReQEnS/rK2wqp11s/zJQR1PHBvH+ox1tuDksh7CiAurL6
eEstumYtVqbRlVago91QChs03vMGmgVfquc3zYnHKK05sIYCFrFnNK/8JWOYQJVYZ8qyCB2rDweO
hjTmJeJgW2zSjvVq0wFHW81cYtCRZhqqdLYbsOB+02ujFrGfO6McoL0LCBJEdVhhYoLZzBdFUZGX
u+wFVZtK709Cg0jvifzlXIULuif1OfgH9/hy1ixwnmrHev0ehla2kNHpKad1ngq8BSPU5qFzB0nL
IuZQycseb+tR41pTmJL27w+9x40yCi9aHCEVRGYuKLDTo8J7AulNHJpsZDxWaTZkWGoYhut4Jvu3
27tXPKhHFbACgOiPOQAf3McCvRS+3msDAyOCCSqyOKlyWE62TZWVY+GxAKTUAuBgX4vfwCj8Zv+h
vqKfZ1y4/87MbmjFdd4chRR1LRC5cvC26MMtNKilx2UdAJaWVPTtBAeTAZ56cgfeibXHI35axwUc
4SbkLXqG+x8EYYA4Ro10pUciNZKXdnCOxbfm4QA9mgnrV77ZHIjRQ4CzZyCfNDuMLefxGWFi7gXe
9Gy8lWL201n3seWqJQv4UYchxfSW84xNLxoo2plDVttpb4l43PEWnAGlsLLLciJy6vJB5+nwutzR
vV3yaOQogz+g9WM80W3d2or6t6EL1xqyQRXQ5cTACRzmKcfg74ywb7R01ienTDDa6h5uPq7LloGB
hUBzG3mr+j4jebhrug/oX5xj2cnWA/m4u4qDribMpSYIw/UgxttBu+OHqxxqJeHXzyHYsWervQ2G
UnxRydTYuZmHYmTRDryvacDXs267U04JGw1YZsRYweoe6DbWOdRCxSwanU3rmzVorP27sX6iY1qO
Ms2vIN9+jn2dp3z05bBHok9X/YZgMFRE/D/LZYP1mz2qcZRXBVt2KY22yl7EIi2ullbsqrXtp25r
ioVdZlgPxS/B83q8hQK3hn7Cmj4gJFI+NPzoiHoTDqkTDSfwPuGRv4Q8ihWB7hqdP6P8/g3IF60n
NEs73cDJQ0RmhKybP648SN/uCmWGkZ219hcAFf7CMCW+jcQeg4kzuSahMSSe7j35y6q1LS57otU8
7Cqr2FZbVyuoU/hvWEvY5LHxdTJ5CZFtzLxazO1Qiew3jyh0DBvYB3o58K+0UekY0BvLeUm6xRNc
ZLC3kay10m8HnNsW4GRH0LofF3U5bhPm2okgHDC27uAJw829LkB3fI5YCo8xIC96AcJ61LAIl9P4
0NtRlegLAUV1UtRCc8gzhdoKEORPPnhHrxnWeW6Q4iyW0AlVq2RlT+lPF3XfDXF5KwYPa7ODyuk5
dbVsENJ9n9joWZnqfTzepcsv89/t7v6vvhXEhiqbjYsB6QbzsKgfUYIAVysp4bD8HpF1JTeublky
nBr90KNm48wX83pY2iQ2gi3roAJgXupvcXIR08+8sjyseA5xqwBlS+rI6Rmps3i/D6ibtq41WB+6
yHY7q24gv1Hv2Ps64799k3gj2K4lhldsP1oc43Zieigm2LqmnX/kUESI482CYZb7TuVSxTRG/ykh
cthAqjYt/eKzzUVEIiRecnPkyQ+RAbMObmupBKRkgpseK3dJbWg79Zi7+yrlxGvdAWqYNyKcDEnI
r/hZrSHy7Ck9zEz8+UWptWa1B3WHEhkYkmCODRrj9gj8RMOoM5f/Xxxy1bVqT2jkxIt1B2MsECn+
1hXxJjeX8kAHBuUMPC7qZBaa3kT/jnnOO/rWAxeUJvVvg3QPcoKO7+Dfct8PdO8ReCC5JOBBJ0Gt
5+sPuJdrZmvBuybaRLHqwMJIS50tU0fo9GQYCd1kOtPtWODhkrKap67mQXEjttT5AtH2FsYupZnA
Ijr9yFLLJjBo88qPtz5wkCJAgJKpkmtVN1mVv8+XPEIySh/zhYMON2H9w6+sdRRmt/zyRF4a1187
ePobvtXsiicbRNRZQmLii5SkGI4NBlvRQOEIIb2PTrXUi6y7k2C6WQowYFXdcs208QD0YfjQbKpv
SJyIN3e6Zx69Qk5n5awFnGN4flJi6S+wx9Z/N1PiutFcAQ5C5DHBTqGzWMiibJvK/LZOY2sVhjPU
X8xlhX3fkt+pAU787p06b6vXUf0uH23nrgsfi4+LgPjtfr1FQ6jvG8OQxtnix1ObKP+LwCzuY35m
S6pEyWxT9idrKFT/x1b/cu9AMmhzBlwoE1/YskjSNvoHiZrPIsQHO7jruzatFasnvaHhoqAcU7HG
HK6NyZxbXadgbJTIbD9PdU/SpHNKUIDYSPfgA6JKMjaTmY3KbPQr82x0Kaap1KSxkptmF5xe9hQr
iUtqY+R1z1DJ5B89XnXQuHxX4N6fQh9w8T/KUZFTisHFFAW2ReO+UKyNbjbVIMx9VCfVfb5p6e/z
QPVx0l7L3/JC5xhNSWCxdjsniEMwHmc0++e/m91EWpFGBHeomzFLQf6CVXADBSjx2ZM54wX68XXE
/WwhUOGkvvlPMeaW9uubn7n+dHbpOofDAyJ+2NqY0XKYyAx1bJKMsM6HfzAbxl5mS4cCa1VlntGn
KyB50QnVJEqfDTj4mL0TWIE7N/OCmdSoH3hhm8k2ODKV6H71PPfABEufvMAAGX65eeMTBdN8XzAH
SbaA9SwMLDBTfkYd9B34cyQ6Jgt6+W4eHvjN9wLEXtxpVweG7cl2z87sIJKoH/2p6GsY8MvRkxTH
/k8MAw0vn6rd2qNVSZwHrU8HFwssCGLeud6H79tkHxVYqxBX6zmZvCtYCkPu8AtQeAgorsGPX1UP
/Zbz5p6G0fJbls3Fi4OGkIUKVxYYo2LuWqRtOAOJRiSZOoikQQDbuLUCM038HEG/IlpdzksQlJNc
9At9F6I8ZZQcndwUR6ZDzFBwfcHeHHPyABfylBXa3m6FyMOrwIJt7fEatPLPhcic2y1W17VfMsuX
VoLp6VYyaZXF7+lZazE7Ut5r/h1r1zV0t5PgqiyVXWizpn1vXJhQKQ+Td5i3oPH7ZSwro7c6BMKM
Yu8VqEixQIVJ5heYn0xPnVaRaUhkEj5aJ9KlUwagdM7FAmr3gSpp7IiWszGyVOZ/imjpx1R9fo3h
+vjLLoc52L5iUaxnAnXlkoXHJBgEozMCjSHqW4Vss1HnlPcQf9eJnJTisjU0moOUoURlS15+zDwz
7MGRc4DUcRAZprErW4AnmpHRRgUWyUN/Gpm7jj1lQkc5GGb41sncuxX1bjGW+tWHs4vyHRXGD9Z/
Rm6xq2BmIA6WeZ8Sncc+8vOoBNddBu8S1Y9/1rQYOWvQv6IUerBHYi3Q2anlQ7L5qkBrYnnkwamV
0WXbO9kA40C0bRuUI240p023wplPzmMhX950J49+zz6ETdv99k/V71RRHF3FhCYhusN8jERcGgZh
pPRAWX9DyD29IeX8a64qUfH+GdXCf5nfe0coSwlHAkSxv4DK//KPx2P/mcwX60NDFIJuzEBm2LvJ
Cw3JXAP9MNdG64nj91hTS/xCYuX+6RiRSCBxfY/7BCsiVYiBvau3A8MHnnlgjGgu1XhRhAZ6tObE
cVMQQ6xzAhtQnBEAvz5Bo7sp+jjmJM7JNWR2Sa19CkEkhDu2RKE+khF4n4pM8nDca2PJEXwX0qgk
x4sTggO1Hr1Ra/9Z5P9WaJcskdFJ1NW81AoFSBx9VPIJr+SzFSDNVAPYg7iXDO6vZ2gddfeBrmv+
tkQi3nBn3z36/uiJwgkceaTpWKtMICIZ60o44CYwJbhVYZwaKf6wA2m2OCpRAZosoZB0tWU5YpeZ
OHRk0uLm96PWwU6LgACasenWfTyg0vLwSU3avYZxGQvZ5W51MyDZ4rMLy3+4imcA7gVZJxshd/3W
sjf+4xZloDkzam4RiM2ezdI/HzNSg/Q98WQ0y9WFBHL7TnQwF5evLKigm9163yy7upryucztEj+x
cVPZfxsCOxpRHM57E+X60lWlPRzLTx2FPfHndtfEM7GiQoKFxqmvun5bq/xM2QAljwZM7iYH1Ryo
jFD5UzZcP4tSsIAMepbcC5aBinMQ4a+ZR2BYqTNLhg0L+pig4iEnciaw+ybJ0ItC/bke5NTo0yXu
rxtK5RuyO4WWbIn4R6e+/4Ey2FlE0QiLjlQzKDeydMumx1C6D4IQWezZ9VzbnTYpM4wMtBoTWyTA
HAYDWe+wD3hmVFXasEjjGpwbiKicumJ7jVBYi2To4Ka8Yv9xFy2eT7/+iuw4mtK7Mz23TFkf1vky
aN5ZfUJKJWw/9JRF5BsWJnmbDHo6zXAjrPGwaeXsmOUcGf04PG0izRCY3SEAPlT9JSjvMRJCQoOH
BBw0eikAuB3FnAAwKZ6smoMq9UMUpmG/FAg7paEui/3xbVfRBGfJKg322rFul/OCeVPPJWWazk1B
vxkhWGS0CBT0H8ZOIrlUFwmwroiuJWhDXnmcz+znb9kNMciypJ1f0Qg+A0ZikrPKMCJMC3583PyK
Bwzkm6M+bZBfKZJAm3zqvBSU+aLz9YEseA6+flncTjMzX7nNHmMqT8ctu614vKmuJqMGj2UT4Y6d
BvTslwca9sPdKVjmR8oNl+TBPj91MKV6vYKRseB2l0wylyvgN+kVb5pLz+1WL9L6EVVSIlL9SA6o
7oIGNnW9n0lLNoSalVIbngV8hcnf1zrWMj7Ft03YKxxUo1Coom/Pc4JvotW/RTSTf4bl9sWKHxM7
H340WVtAXVbq3iswm2DhrtLR6i9fo05sThbHTJUsWlOH0riUSverG2DwFhzrGoncZbUEwfb80Lr4
FzyTdodJXZbOMMtIlJHLw05aei8G2Q1BG1lpjvfFg3tJ0/oFumnrbdTmx1JNP4sJpm11S/pVXUoU
iXl1VQd5VIFuDWsGXKs7jX/xHFOZyhjs70OphLe+HUTWFZMHS9eDDwsMpxDJ+409OGFYmdeBHdce
0VRK/1+9p7hN7WencYMtM6W8yL1I+o18Yg85cQfQYOfJxAylG6Lr6evn+d96SQaJKJJyvScshswp
Wevja2l+5N1PllMKE8zL12GiGW+JgHXm+5vPOp3VxshG0PBX3CX0g0eYl3hjEh6ME68+SZstRqSY
Ubuu5TZi4FNbxj9T+eNhZ2/KOrxaleXqdswlrOl2KH7MgPilKZQeYnPFwMIA8XpzQ+DNMSN2EFlF
oFVrnZc29A0saG4iSgcDgJ13fY/IvzxjCfyViEdYUVmJi0ZioM/DcV1ffuAfZhFsjWlrxgD9/GcK
fKoFIRi6N9O5saWsq9rFLjy64DBpdwwa8SN+5LS/lA5A5ly13YMGosn6wibNj64QOyvP9oxPUsSL
TMaE9LYUEytTmS0HSmGCIT6XiMNeclzVcii1dj0OjJRrQL3d+aTTHa9KhpPdypnrXnJf1t/trr9w
zKA9G3pzWLxj7RpSh5yP9Gzdduxi/jNNg2SOy+bYnZLvwMQA0AaCo4znXjlDh59ZybAPB1X1oMue
Ul5LVVzn1xB/cDVbEQsJ0YiAlJcSRYS5MCe6mRxTSB8txOuBE8zxqVlDRZ5DtBtaDjbp86mMoULT
3F2HY27s4dIg8v/ZJoCi+MC2y5QsRTlzkuRj+kbMbQF6PI8w7Lxg94ZC3oGk9WmOz/RVzK5FEIOp
EZH0bapH8Ci4IHnmFrzPNMEd5nZMqadIxCFwh7GZdyEGHp4L+Jb/ShuoGCxH9AOc+CmBkPj5U7BW
3zQuiZrhv63k8AuQpMw+Bk/zP6zdYZxRyw83y0xfU22c8YdfKgGLFyM7Rb+2O0bRZtaIiET3kmGw
kfqM+0dcf+2dB02d3IstPObStmjWf5nxNqjtbywHCYCk3RgNCZR/UEGO4faOtMDM137/a8cjbS0h
Vb5U56ToqbyTlwsn+shG6qxcjYezyPPeKUs3eymhRHhX1GvLgNCoxmT1F4BC4M9wklcXzilmGIKJ
GcwmP34oVhDumvWx2k/HW77wqtVKoKjb/aiKs68Xy4G/UFP2IvMQBRX08s7mIExxoT0yz2ALu1T9
eEu5xF35OhEh++MFEY2L9QS+ICSr0jtDK8eo+3z1QKiTwBUREkFrnK81Q+/0e6vaLLquDVkYjlJX
0hgBPq5Ge8RZtAeGzWLBSuIcZY034fQH2NazrqR/prru/zVcyydr1qeNcdbZltCOsoneD2cyiBHO
hZaZqtK/To7T+5G9OlM4CwsuzqXbEH4dm8Cyjlx6pkFJar7Xvn2jvRBslNJ8s0nNsispYGASLPsl
FcE94rbpe0GY5Sm9SwqArohvs+CjfW3UOyqicbligMYHKLn3fGnSVhp0+IiWCuwhB38D7E0CnD6+
UQMPOdttEMVuKlI0/DRN3Vkm5iPtNKlY7wV4AWZPAoEiTl/OzDbMEfB92tEq/88FIwIvj9eTaQtR
7mqzqCdlmZiVZCw7ebqOalomUMaewYpjkLqqfRs0cBhcNbn7LgL8MDLOhj6dzYMn4LFLulqkdfX4
EjcGmcZeb+M9X/MgAJVLimp/6X3bvBlDPu3pxc6u+wcEfnQY3po7zQ+eOB1irwhqM//yi+9+g4y+
FGn8/weZcaJofsa1gZ17efZsRWSfsFJSzSPTt8Sc8DCtcVc0GWwGbMFQmG+VYZ//BezToSDAHrdv
kvRFq7/vVhK/0FFQ2vnjurdG3hAELlCcrpc1JXAli0vj9SrhObq6bBbb7Lhw5/MzzcGsKn9Gi9u3
QSyyBtLOorAYEdxdvoCwkJnh41gnhmyDMGpLtQJPXWwg3+BLV4son9n39IID2mKn+B1x11/0tfS5
YOI1xfl9PjwTWQhvgvTsAx9CSFHAliiIXo49sxB3GhS7Nubvbtb8raHfpIP7cWBH22XqFv3zVrxW
kPU6XEU70yMl1mSqWnD1FrO6Bb3WS9O4fSFqSUoz9SNGVK+ciDwHKTww1SSFuGhGXPfKozfpSM0Q
/jS1gyQ0iDahj549PJbZQrHclq9pJmeFJQFbzsCvsXVLDxMlTGP7yMozFgkPlskuswfIh6DWPfgy
MNz5y10G1Ywm2k/pMh0SedrfoSVrjUb/PWuX3T1C+O4crxvsZiOB6rNyLhY3jHNBfkcdx1tIDVDx
yEBwU37mdAl1V3RbU6NZzRO2tuUWflGM9p1VxkBkA0cW6zRHlPXHnp0yU1n4hpWF5LL5yWkNZ4Ch
3U0f/F+9Pd0oc5eUOc/2esCW/mXosgTlTW34s+DbLXSE7y2AQzYlZJSOuNzNgUogT1ox3uHGupsc
HKaWbw6vDxhMw4NcxHCd6Manu7Dj5v83Xk9iO8vJ3ef8FSysd7/pPtlecHg2QloNIYMYd3AbG/ta
mxkenlVRCEfXJJYJRI47PNQOVGoihg3xiWEayQ08CDdkyMH5V5eTdAZfeLTEqNtCBbXU5ic5w9Si
l/mvf+iTSYqNOvrWRoliv/Q3aWs71hWAoz0lBWkFUFzlxf0b/ZHQGij7lUW+tDhYE0lndIP0IRuX
Joxw8Iah89U+W2egzjC/TE1rEKHxjs/kcMQJn0lhbq0VA2XUWAGSsEOHLmmfrV2j6oCejw1n0Ibn
WYBY+gf2n5RGUZ7hntJnuwL4nZ222OYv/zuzscYAYN6gBrEZpGVVqWfKm03G3jNMIthoiQ95dDDN
Lty2JBJlbT687t/iBf1e9sj5y3mkjf6ozkXliO5Pa8HXwrHfUYwQ6KD81JnPIztmhFGAwP9I9j9m
sElUY+FvYfcVED6aX6v2zECKH4q2+aS0pKaAYYmtJ2NUiDcJ7RYrbcvqkLXHJUd+Cm/td5yyXN55
5QmPviBKKmi1p5q0qH4YxrrmqsR0ZW0EYDPhMvEHdQdpX4HIKCEgHYqV7yshj9ahQrWjOy0xOTum
IR0l1QqSqwho99vxat/odSRzg75WHZ/7YA96puGoB/kVPHTwJpL7ggASnmmg/1lEq7UhZkhb/DWZ
mHTciEfz9xjlEeJqX4dovRDsRdtZ+j0HCEOd75sc6VCT7f6FsbN8Zwshb31lakUUr9sLMv8RrIsS
BZ841gNwzp5j13ZoxgFnUu/bNI5jwOaH/MKmElCdd6+SoiprwEAUHZfUL9HkSjcBhDL34+MuApB0
iLEYY0FoCcPtqMYPrbiaEAnKTweM0e6/brUTcHGa4B0j7ODV79P2jvhw+9E9eyeeQz1dLXUNDR9I
odV8et6aCQOhqmJ9SaVnq6oMnUORA7yb6TEZwL2Uer7+V7oGUulgCd8mSJd9d67N9sXol7kmiiWe
hoFG4pLbCSd1SAaBJNboEpxq3G1UkO2j16czDwzFJa/BQZ/NkDH+ibpowTWjQdrpI6vDMy1xVAaG
IKk4eVPaUPNE5GQLxm2V+A7gXM3Cb7567RXkBEiM2hbicRuYxxokdubqbCttPFXMNvsTV498DzjF
g5j32WL9V+5dDhSOJAAb8cSY7JK0AKI2TWx3pFlwmJF4a0C2NXS43lGBXRdlxCuKqCntUa461IJM
+NDV1rWKCuX85v4a42Fb6l4HJ4hInfqv1ump9LNhI4IglmS56NRRvALGy97RaMBOYqIJeAQdo8vi
5MJ6Tt9qOWURIpGpRzGqKI9n2bfT786FLv5SS0PHolGC5ZdeO/VC0RVo9qbDNX6Q85NJtYip5gdP
zELPGH0yBdWkwM99efepmZtY+QEGTm3Mnklpprw1GNIdfEy9wsw8nc6G0Tap9Kdt8Mmz8I+7ri4P
W5Ey6ArsIRRQHVYKrAoiTAF6yCG1IBwmA+967Wsbu3K2rXOEt0Ua+k6tv/NAGNdlGcuLDqdikzkx
lfTEWTZGWp5S8cdhbNKLMkveU+lWo9BgGeJPmJFOz6iKuWSrFTT9GlNYD+ouw1FPMbPRtW3GO/Kq
kVsF+gwF+9GyUp7Pd57jxV58L37JMUKmOt1Dqoe/AYF1GoovuXTtCg4fDUuIZ/v/BBDnlDrwg0xE
IejhOCgSQuxBieFAG8urAn5DwWbAME5vk8etP415O9NfBLg0HFh0ZSKnZeGQ2nVfMZfPFb2ZSAv5
q09PdTvpvKh6pNJ7X4gaL503uVUc156Kncs2X/X5ABAfCKbXZkjfLht+73JfCPYqv/qNhJ7nWI2c
iglMYbSGeRPhhi8+V4h0AHQ9GyrI4oy3B1/CTqDJ1vvM8h7mm/Dl7gWi1zLKEnem8aWu15m4aYkm
KjtIlMuLsYOXi0S7Jk3jHYMMqs5AkHPZu63E2xnCocAxWwxe5i2dSnPe+u15+aaVV8+7x0u+MIWF
Tm9ajQYbXSPAtI3cIZSlRq/FOdXJCNszLoToDlNJmvhxa5rHY4RuKFVUmWadW0doxeE0Mh2Jy8tR
EaHhguuvYNx77QB28mGr6MmJ4qSFMKBFPDD3rAnrFUlLMnai4gSUtpCuw06I8Yfqq0BVlPYNx3yM
tWPWihwwBBzv/8HNN/QpQbKuAb/YQ+EzSwKWr7HAzPNJLErgf16hHhnjGRPpvFXQceFYUy17d0c1
E4YXj2Axdnih6+VhO4gQB/8tnlXOxiXBIqpEu9DHqDp3Ev/f3tCZZs2cjN7tBQD5OdacvgQxH47o
b1iFMi7QnY/vD/ezXW5Z91IYixAJXTY7OADeVjhRyTLy+xVYy19ZbGZRoAn2eiLVLd+4zS7RfCRZ
cx4ANinqEoPjDErxec3mjV4ZJA0j4zDhrT9qdgOs/aaqxaiN4ZgkREa9DR7QeXzBJLKBMrHr2Z7Y
jQhOd6KX93j2f/Th60twwkcY4rnle5GrgCLuF0SDj60LkxBgG4nGbvrH05dtnOz2BBouZ65HnP8e
8TL06FXRzO6EPRCAAiavkI1iRgiudPFwwkbn4vN8Q6i88UGiIz9M/yQypQdMcRO3OBTjQJC/PfjV
v1ApaLSC89ewAJPRePd6hqOxv5rCtPqguUevpvhLRdtwD5sO3Eu656ZQF8tTO2YNEWkS7T3I3KXo
tkKcBNrGrvL1pY66NwAc6R/4pKl15QyKUuyrb8JTnrCO4Bpi8tX1Wg1kZwFBFpNYN8qHBVoA0Z+E
VZCN2aY1+rj1cQRvLdz/4TW3rFwIYwBgGdglXpTmOBLOtdgNEFPi53R5I0v6mI5+1WgbAXbZU2Uu
QStjwjW1mqyyaMIME0mQkTzSA2k8GjN3vSARTpZSbivXnlzBA4biWw5jNOF004T7dxRHVsdA4lgh
kR/CD01p/HjiFUiBKU7OXj+7rO0ctQrLvq1QRQZGTjJzM5Tyj/pjmq/Ps4DJvgn3NW95B3tP8cwG
6hgK9slohgApeZ9ABkbSgIhFLlDXv74PobxDRwgL5k6PQMOqcRmyDhdgU+HY3Pey51AsvB96RTdI
qEGk64+Ohve9CYcBYS+cNhT3f5K/kAxaCYjAoYh2+T6BRO3QA/y4E1NU47Z/uPXbR8KVwnWhUf5P
/SAzfxdKaYllTj2sm0+BbhF/csednKomlyGtIEUYhaMq8q2mWXJJ7iUZItzdA0Jpx8luroN7SgyO
UVO5Fy5BZxGzYNhFLtTTcxJW9X5eh9gVeg0Q2e45gsFALgpCEV5M8PyHaMufVIm7FB3h+/F2QUeS
2TbYW1YzrAK3gDIkqO/WSYcLsfHbjwW6Uf4fJayUSLseKWAxCvysjqJYZyoo7y1yr21xqID48rUT
qGzUNQBHlxJlE2HwAjFwlG6Am9zgQOGMP+2fgPBxBmPYwCKT04LUDK323pZUkKvLsG06BZ8rKvH9
0MxCX20dqpQ/m6DdEE9/0yOixjymBFwW6YPGt7ByyNxv/a50/n5GyKcp1Adzcq97uwRRDW+w33vK
CpKRT0qjpZVCKEXGB9PEdqvtuZsI8mD4+SsZs6DkQKQF57Hb2oMymkzGzSnfxpthQAvU7iXTxfiF
8JcpyjWN5EGITvbH0CopO5rJBd12uk3IkK6CzYW33DdKEF2DPRVDH3t/YCi6NnN1JUTgfjLa22oN
AQZyiq4SLpORdvHUW6UYwfhemiSl2Efa3I8HCWELv7jy7sN7cSGbWA+azPgNPWTiz6uiXre18lNv
9KR9YdmqwW7Rpr3hDVY2FCvdLtfnDzOOvnd2Ov8oOJosmtaGR5OYvkHqQgGQI1/uCXFAhnVmeEr2
0i1UwWhQ6QXPGexI/Rdc9SiDX7hPlGqEBbMRtOkvhsRF3ryrCO9+OiAFHdwqDuNafUwtOiHzHldY
6NuCvRWRH9HxV50urRrpVuz5/FO0uiqA7pLoZsfS4MMWezPJVcFbYmVxxodNgFLlywytV6Cnxz7E
FDUqx22cJgjMavOUSKAZbYDtMHbX6xOrScmKOu6TpvEVemva8lfDbxNsGnXMa6UdlMi9kzEPSeeo
QzvG60+S1GIUkCQ1yWgZCgBgglOTVLlhzAR2UKC9dDusELJsIe4CYByCYrT1bsksPf/zZgO6usNG
qetZm/MKpErFH5m+omVCWCeTxZVYkTIx0cNaD2Jh6wP9+MK1CJGckU338SpG71B3y+d9N89oyBnD
zN1T6CzjsE0uxtluCocBdB+yrWIo6i73+fYJE5tKEPXu7UIQd1mXIixzlnRfKiujnqagDAGV0CxN
seRmalnHEYVcVFwkK4KA70bv6Rb2MOpauJIUY2wAXdMk8x895FbjHaegrC2isT+Mi5sB5NdgdiLH
WU0rGRuE3zp/7sl82pcLZSRZ3x0DrC+tRPUwncL2x6MBSeJU5KfcujP353G2SDCNvJaS+DuQuXlv
p3QI7qLusjgkAQETOuT8PUJhozHXHejoA481MS5uYuaAqQse9ILIbn1HCSC3RvdQgz9WuJehOFc9
1ae7hMJJp3+9WQ1TIATP9R6UagZLE/t7GgnzHEF+d8HiXRlkH0gF/SKcfxDDM8vZwq6C9XfqCVYJ
v6pqqvC0CPMAUr1SUuTHS4nu5keMF+ZDTr9C8Q2tcC4Qh361ssAZNXLHrjbPzYl6QmPe1jX7MQUs
xKvPF0oXBD0GPVnPqv45MQ59cs172zYdSlNJJufujwtfXxHoa/kDBlnq8i0RQWnYw1+dqhogowOP
bV5FnCZZjwgRQCQihvEpAD4GQxZTrX5b+FnmzNgl7vXtdUSmLcB8avxLYaJALjt6x5zPDbLQdwUl
gY3xKb/pQE1iNpmMU6R0qd+CTE1/OiktL41rgFsfYf1qtme72iQ2pEcph8jYNsglmnHVQpmmUQe4
S7iYcJlG2s1ISz9jQf7jkL4grDSDbcRscyWBVEcHJSh96vTSEOp9L4Sw7Ij8XoQgtFZpynW2RIOM
DsZKfoQBNZZvdmIPhTfVjKRNS9kzbm93HYA3/+hhoTdTBM15s50ZiJs7xAh4E1PvbDtv3gqVdDI5
yavvbhj6vSDN2TOnmYdpG2wE6sUuSyD0qVW4g3aIQPnXWfLGFaHHyM3F2U9pxOt9wOQMmk/WeDCH
19SohU+vBbyOWe6wkKUWMDWXpUaMsabGQP8B3lwQkCnpPNnmZUc4CVmV5txxquwa02pI9japbYrs
5tMnpwXcA7OMiz1oC0bMwvjpUEPdV79M9M82JW86qQ4AJryHYyIC+0ci2fKS132Pc9yP+Nn9lsxt
lb1RvEdP5y+pOPEfOdfhujMt81Bbmj/CKVVgx9nFQv2L7DqO4sS4rBb5piuzZDT6+h47Ri7BqxDb
W1B2qdjoJPrDvMXHJj6IV+o0IFA6QHA4EJsXnwNA2522XvrmVrL6Q8fwKenVrfrGtFnk2t/H2zaX
/KrRlckL0A2NhWSx9GqXOyYx0TEXSP6xptl+MBEfThSZuSvMPL14yyBYPHKNjLzMbXo9OvUJNAFd
GxAD2QXudAy2fHaWrD2x2bOyyPbswIZPSs6uSm8+XP5GtzLPweCUFR3onGSAGVB13860BUpnY3Ip
od9jZ6You2AMc0QEenelda++P3jAsEHUBDqWbIsvaGyBKM5zY9i8vM2rh9+LjCxfsYwliRu9GfDq
sV05ckBYryCUashx1yaI09MzRYClUekFaLg2qZPsAQ7jcYKaBfXEOqi9ZvP4Wkcbp53Jf9GiO34E
c/KKfFWsQxT1eJa5nv8gpgTd8+6bwwvIK6E6C0qs2MkbC7zHUXcRJVJzXBMuUYUibiOyc97fKYYZ
IXCAD4BdBdETQE8itqfK6zW5R7p81G4ogxny1WihCHTQNdyCTo1TmaLFsu9+4mX6l+Dp1OW+rESE
c4lf4QnAjJoG6Y8kwBaIbsDFBX4/2w/P2GK9denMtT7Q3d5Q0KCMq15xa0Bki38+v77OZrwln+j1
Xzxd5AG5gA5OYukMNiaupkHCySVCARFgVj5t9sAfLmBNuVHVhtkaI18WBnZRYvlr1iRboq0wnKp4
tCuART6nKd5vkGG7Hsxk7VFOPFis1UUtCjjpZPanHqOdFqLc/EgOoXcPZh5NfrKjVxTKXCnxG2Xj
iS1kyPdKFXMRdzm64+XoJSPLdpj1mDhUKsWfWrR+o8wCotLkyHjKGQI2oHynm4P8H3SCFUWStVt/
0XYMq+zqMz1PFhPw3Dx9i4lLhCKk4kGuWA39BWqdId55jMhHjawCLb4iMAKtkHyAx8XEXrYdabAR
2hde66pA9BdnFvsDVGZ3e1rN2LJsq7iKALsbsp7mY3HeOQuBUgQft7somKhOg77RYYYe8Vf9nVcj
Wqvd0aji/w9DjfwE5PMNASCRJimCURc/5pvMjiEUqRl/WNSyFMAVff7sjYngZt5zLgVPLbUuaV4W
k/8HPoA7qzVTztxPlFU04yJ/iPLgmpMQtoDthBkgd6u4sVUuqRjXtpBrATNNogFHIcZsGc9a0wPM
o8NLr/DFHTKSkr4++4c4kd43PP6i4J2yQ7GAGXUOv/hw4m1qsgZiUvEsds0mtCL3B6Byg0sHkr88
Es0TLWnN41pLY7uUd4BDS3fATeLtOpFyKRSDlCP0jz3q0cgN6ifkT+mVlfhbcbnI2iE4j9Q7LCPL
MsmUHzp07g07mZFWJ5v52BIuPrOSq1bIbkC0SRhfGPz0WkNbCYKrBp7kjDxUxk4UC/26AAFGTQ49
4L9KKISXNE12bto1VWxLAL7gK8FJIHhfj2XAKBiwpGIlu9trLyKTDScpDUu4x9dJjLsNzkk3a/9y
O30SIyVpFzAe0jCqsq8bsKJWOAmoeuNlcj+SaKCSTYa6F2Hpl8n8+sKIy14i11Pk8gbHEdYHbY3o
ph5coPkL3RnMOF4TrsusHFA/8ZaFPXCLRuKe8ikPR5aL+MNAJmxec0pP1BdGHmm0EuO9JX4B02ca
Nhgtpr0QIVGPl/tgmDWmSVi4+PyalO/fPL2RW+CSGn11usTnirTOfMwYtrAdte9mESvXxgQNegnR
SSUVjJhWrMTHvzoqB0ZN5pl2kBlrutuYMlA1X4OOU1SEMabDxec8I3YoR/zcANNMVX7zQWxokuS9
1FbtOI77UY1n5uW4TaRh+z20UUGzvzilomyEphG9qiNDK9ps58WjSOgMeRrXnLqYGYoDuIuMEyxF
4i0O48ky2hDbxKpn7iSnW1Cx3aUAEnBpHMd/zzHGxslcaHLtVEvdE0AsWMVntGBbZsHdo/zlW/VV
u6PT2JkVMEMPKMDXObfn7UnSTDtnkedm2FUwyU2mvUDghm5ETBdRYyx5RQSW61sZN203ycoaqm3O
Q/PMyMC2At4Irr940IwSf+1Hqe5QJM/Xh/XtZnAZv58qdRGXGHF1xPNT+4JpPxXteATT0BSWZssh
BS+pWy6wgyUdNM+2zhVd2H7N22KVEODWUy4iHYKN3CSxeQVKwFAWSkyTQnwGQ6ZcPwegknuMISRc
bxxlR9eV/LT5rHSfR3sCecxnsjwgeoh6csdYpvdlWbfuqh9uCWFUBGuU4MsL+XFtPCdyQHJ3PNvE
Rkv27cnq+5Sab/ko8zrcWvjmKBtHEHdEErXEmwTGgcG23+ai+C5l7g7kRqVrusfUtwc8YN0xQ71e
dUiw2eMzdQN12GTtL8L26veWLSO1dmSUN2S8B8N9TYUCiyWgCb/0EGZq+le8Bg9YyI0tVFrEkyO6
rkGgFMQI43t+qbJ3eZ2kMEHdqKP0QTvOtSpSxipJJBoX/a2hUtgx7cqnG95DYBBsYGdEytOJmokW
dXjTQi7VoE8O98bu6t9WY+XOZc7fl+m5lD7xbz0Q+dBW6pvXS6nzXYETJmkLl4ZfWVO2UrFWXDaN
E7X59mkjHixmnkCm5JxYxY5DvaTF7SfurR/iDBzTasROvbRa6gkDzbbToZebNl6Bw4K7nnYoVJYa
XiFWtLelD+OAQANcAvSyEiuiv/RctQnXMeYVmm1mFe+dbLy8qQLVEpRjP5zSbl8O6PmOJnExpqvu
RI5BTxxuoRa6L/JpJrprUL8whaRc504yrKJfCpIrc1atttwLGz+JpJ6eH/cLFFPOxHLx7VKOieNH
vpsJMI3y5Dw69t37oOsXUizE+Yw7cJMek9MF4BuX2Irqju/HI0yZTFGvvX30zh/tLofYTvW/sTGQ
26zPNMMnDH0bOdo3KZt+66y9/MA+EfoPofVWL9HwEh752ZgTfmtfBgBKH41BjHKT5afPzxKkrCFU
TMHaOde3PqMKwFlcBi3P2WwlYT6DFre3V0qL9pQSMaT+hJdBEkgevjtdw41WTUvdTNlVkx0zrKK1
C8m8je8sWL0u8aULeLnzMQAk4355FYI49RkIomwmK8C94y6HGANGEEajbJxPBL6vJtyR500Wdj4z
qGbsq6q3Nrb4ZiDkcXIPpHBrmzsAHZZzNmHuXRcTaakSTseupa/n+Y9K0jLJ866SORnYjQAU2R5h
feoaTed4ohYxXiCGAdgoYf4rDqORbJadQcuzjUoDYqEeUo5AS/tPlPDXlHqQtKExemDYskuP/wId
6XP79YkgNseA0RoAjzdDGdyjBnioFwJLJuLCbqmKJe44zo12Q/65HRQj2xfNlH5PaiAlqSSqOHUU
R7B2A2vwiiZD74OwWoNC7xv3FW3wnqh4R+051Trj9KYvUsnd3n/zwKm2bOfWTLZ2GP5xJgEWtK9Y
TbFOc66fcLEnUnM6HsRpJfxCqSNPUFtqINcz3cWviFEBLjb1qrTJSjhpDt50QcuRmZg356mhgIMj
1z+u2MsiqA+t/r1metzeUvlnu/F1H+shKh7o9rIT5k4Mk1PFciIoWKq6PInMU0W2NhCBwJWfDRpG
JibM2AykUYIyc4NAykhJp+8haLGzzTcKFZ/SCPRybNeaqLxgCVLU+Lk+rGITPamGVaHKfXoWusZ/
a7M7rt5g/I3ijG4WYRxEsz8w/OSeRuKvZGH+YtPbW5OvlLNDrnWkvhmJGut9jNHU5JcCVoyQdMJz
H9cPdZKx0g2zZA4070RgsuOnpL5RvYRG5W1c21stbdPk89KYUEV7dhM13QMKTgux/xRf5EzUEV7M
BHO20lkRqteLTdTQcdYzspj13rsHr3KJpR7ubfObArXfIsuhMSlHIN7+iBAevrINoEMGncJMlXCG
UL1Duladk8HKHzUFRAwMigDNeLqQTLGpJsq33NWq1IdnwMe9OgFOPWu3RRzNrp8+2fYQ930IgYmg
TX+itxKXfh1oahnEF2OcJ2QFlDQBC5023PAHIAR33Ea8HasYG+cidupMcwlyrpOeKZj6bxjEN3db
Brctpm0scJis+XYwhf6PK81qj4Fm6zCrEsxkxu7mGJu9rh42TAaHQVNGrUa57iLoqlXZfu3/jn6E
MBZNcqUfUSIOoM/Z0XF8OnGykdQIA4qGBZnwWXXuPvMiotMb1Z69gHNx3iU3jV9zJsb3610W9c9Y
Dvyrg0OLwwy9fUXodPum2NvZuhlh26jS+T4ZmQx7djCeUsSnANUPHKVKhmvL8Riuig4+zmuef50/
TVq3GH6KS1hD11JwFxLv/706OQAtj2087MNzmisGMrqn6CXIBlzFABgiMxOLOyOHbaOvPZlSKFDt
VpBNaWZUQ/XJao7sqxEUOjjpWOGfKcd6lyZBpngI0J+gIL+ovIHX8ouh3uqs7icLQDiCZhNOto0L
aLP0SmNz+IjtG3ucySZiDf2THMYgFjn6qjmr4rkAGn8N1NiYucP776koRUoEat71YY8sdoqms4M5
8qLzDjN64LWgPR2pC9Uul5bO9QCXJ071pVe1vrPWz74A8NdO70PekG7/WpaBFxivuJb/79grctxW
nuDQ1nsp9fssung7XKRa9hM4LH2COv9T8jj1at/xN5GLXDjuFhTdA742OB2FFAg5QUVVob9jxwXj
Ol7vaVHxGVWBqqic4vET1tk+uPAjHgDKfNt+t/cRGqd+l/hFzGfFxYpJUSTTaHDx2Pq+5vK75co2
yVQI1iT2SzhjrAS9YP7PgIkFR2Rx+o8pxvTZxx+wLrwLQA1IftXJF7mrU9Iuw4gj/H1CEGPCBInF
i75JjL4S4XqKqgplOUoyH78KXekO55bjdXzmTfluAWpMzHecQg6pDQnqC/Pw7/GUKpKAKBl0JdLc
sIcOrJSYISKuBC0nYXSccpYm15As5u2Qpj484x9XHX/ZLkmlnTdl00x8ocohJeQOhe20oOOOOuI9
JVa2IC9bU/PEXK3LzRmE+BnMvhHqk2CoC3jHkXFbOiPdRzgHzvL6iBumeFguDSlVbvj+V9m5QpWZ
wd7541ucSDnSZwBinw6JV16f9oW2FxKoqOeBPSak4EH1o2xsQc+yMteIhBuWAPEICLjv9QBIlPip
xnnAMvH0Hp099ym1MRqHd3TlXS2WVzzsgkO61cSENJJiVFCUfBvv4MUoFEQuCpuV56PxeiyPdb9B
0PsiOjBDNA/7i39s9CPZjU7tut9dcGu5p7rkUkwpRIO8x8aCuwO+x8Bx9M5jClX0i2zrIv5FaZAH
S1h0hXO7+u0Lu+/M8ZU9dztJmcWiubVvBDTGu9vO+6rzQi2VuqxI9eaRaLirKQ2Pam4aqZhYxkqh
y8pvkmF3pdQMfg0ZAvpxHkkGMzkMVBizroNfyScuPaRzVGsO99Px4tzxMTMIEaS7tvdFmXzG/Ydc
L1MOCFyoAJGIL8p9P6PKdeZkhn0LfYv1gm3PHg2nRYNSIXUPpYbeX4JzimXAqYupcNl/pgOFOqur
kGNJ9M/Z2jmB0XWK47eh4o6HmgfmCW8+6dBCtXBhLYNZstAtR6yquHXzv7gl1XdyorbiMDNVtdU9
XxMaRGIlbBhJ4LP0lMY6qzXRk9jLcDykFDqA80cahLAHi1OgtPAjYMLuXrq/R39SYi7ON54cR/84
wqSQ7U9Q0v9fa4BMe7Zh2vpy0U1nbjoSYUhxacSUuGnZ2aFAfEhJVqJQlP14G0jiwItLlBy0fFaI
YayZqOse2EtT7VVTj4D04n2/XfEwNOdy1qEURxAJjSDYEb71OTAjYw7/nFkLtND0RBVJTyvT5w+l
dgH90Ncur91tHJihuQowpMHRJTW7bQgXjuFP4QMzAaNQL3yK5J/BSbBfGdcMjlI7NVh8uYs9gKgr
HrB2Kr69uiBqCsVEH05c3ox2cMSaZ8km0VhvU5SdPxki7OWPnlAfo2/qwQrvb0MyllWHYN/2NTRp
ELB/jo9jEPJ6Yvsy4AwyjK8i2vx5Hs3fa51KRH0xcLHff/INhbSPh7vCWn1mNJwkxFxtRBrG/Z6z
Hm+QmQ43idyRemKfU7LMTtCQJFwn+UJJvYvpf3MlDQ8P3D4fQa11acgBYRJ120Qxi4YII62wEd6K
7aDSKrk70JOC8SsEwJig+I/Sp/9rAh2dbI1okiPNDU2ITObtjvzt0uytmkjc1HYE+j8iYZfpsicE
B/zzm7NZED/oU2oldPHiU9/9ZtWM9btyTz0Yw/XyBajdY1IluBDm8wVKgNSG3DxgKLzyGJXKZZPM
umOCram03f1toz1mCTCsftaJeZHVM+OpjbD0fc/ovIQ0uumnrem5+sLRfw6jMsAu0uDfrXTDhwbW
xL8JhX2MxFkLXS/C36ZRmkkgURkFGtKzElvoT8gihbQJwYbpm47wDdyMADBtuDIXD4SpOuWNYjwb
q66lSqhILf+k9TExEsmJuPQnzO9NPY/cilYjY4qn1YRxQZrEP2aiHx3PP91ceePJlqJBoFboibId
o9+vFhC4Yn9l9Q6Yztp3Vk3Avmsa9sB7pbC9MBilyqpCbIx7IC7sr+huWZtb6wwXvyFgt2e6pfE/
ZjlIDCjhVdKb9qVvgjzA2/el3MPhN/0zhxgKgno+P+OnNNkLAq6STylWp8ZcOQfJb28PtjFTq1Z0
YytU0qWXplYuciEDN3AaL/PubwHIvGAQ/RGYKHu0kNbXgk68huX7kDAJuJYA9bJebUW3QvkUMOBk
iT6QLMR/Ist6gPH7FXegK+DEX3MSbqJRbi8ri21CYHvBOLe6/Q8RzHRB7PyQNruz7ZrKt4TC8KUB
vueoFrLcN0KRyNudRhUKDZzNDwQuHW3YY26cjyMw0eczFxG2undrt7+QMKonqwCEH/7q11vzrMy+
CjbAIGXJPwImQlThHLISKENf1bLOL9Q4cM3WZZ5xWiOHZLunSM+A9NVqXnm+fgHiVL59Jpsnfkq/
VwnZ+k8eencm9q26Q9ikV2MJvaxCpA+khokl6EyuGwbhTlLqhBC3h87LsRxdZ7iIKCfdXsz2MBGU
hbez1H1KQFj8pwzNGFqNkToWnim8Lt5F1qtRdWa6MCOmlheb88Ia/+UvBate8h2h8qPVzgBQZkJj
wPzqSznhxdS5ykuXGzlNzde8qgyoe2YrX7FS5QiGNmf4LeX3n0FOe4Ei0TKNWPMr8bo3g+VtHtCP
+JngQjgaiTGUejaQ4YERR6iph3PWzi0xvkW8BX5/UzcarF6yfAJAvrtQsjeh+wP0SitxSJL2pMh2
wKSRcQMWBCKSffyni+dpa0KtNIGj8LeeEXLDxQOSfr/ZIVkS3fKAsk5vX/D7C/k+CceQ3PiEYHbu
D5V5UfM0oW5ilJU+ZOkocPEqyuU6tOax5W55LE1QtWAVQBUiK0I+Py65SPw94GMTgzN/pJlu6DqS
1arZhx0ztHg0KfEd7HPS4kVCYRtQoaeeaPJb1tzy87OnnbcTLp21qU5orYkhGo3aVldrF+BePZ2b
CpMFaJ1qY4Wv7bqks6z5/KlfKfQ95Woq3EzNfD+WNtJK+vZmXtLSWggyeqXPU7bSEO/Lh5lVUKCf
nnqrhG4OevfYM7KMPd9sRHB0/DYyOphlMWEtZxOg+8/PVsjzK1hPazOYUtkWPdgpCbSZxR4ldqTC
IA2DEGran2Qat9cJH5bGtu0xHHCCiZbhxLeAJdCXPIcy9H2NdwcR/tQBW8KP5PTGAkkoODzqaIc3
zGXA9hANP9OMIl3O12HqMdirmI1+SBgm6s4FfkvoFUpkJD/lT8H0wYMNJOwsOrm8nNx86kbUEyD5
AXs6xnurebDELRsT2X+hkNEVmCqEPk88BXy6RCgEUHh2PrpKkKBvMl4kCE/MEdhyCYtzGz37ZJYS
nAsV0N/H50qFx9/MPBuWlUoAADGBfq41BwBc0CysvH1deUeMIgWMDQq6bMCN+e/R8pkkk9k+6Cbm
p2asAX9xicx4GcbAI/ZUH/8a1BNaaLIIGV7IKuRec/BKFEfx6U253sErlkY1LoXF8oLKgyRmKPA/
1PpjLRreR7TpT4/2L1eIbTqTvbNdHQNjI71I9tyTTGcP96TNga0jSlx1jItbuKwQfbuEdjzCFrjv
lXF+PF8Qo4YXHGvrq8oipMeBdfUELPHFJG7KYd1Vc6Cg6PGcR57ZLH55gN4T+OQ/P0JTy5w9cnpC
pF//V9e806DVCxE71Iy+e6yA5ON0RQLwBLJUrC3+rptX1tPg72o2IGrX78iC3KhJynoLlnGep01M
wkui0oAR3m6n3eOKmbEAIOa9pAt+/ixlDa1VMQXM8Lh4KZP5ikUg13mO3CjEpa9V82pJClC5ygL2
vOkt44DIlmPtgS2+etjQ7BnaeoGwD+GMqB5EIS1+YJ4ihWkek+12SZjGEr+RYOhF6s+SCca8N8fs
b3IwnnNXOGID9KecJ34Ghv2YbPD/3lSHDKj8JSN/H6aC32z/20yncouqRnZ8PvvFY+zlCHm53Vdx
IPbU2gVqYnUbgczKFDkjyMsQNw+VvPvBzPR6HMpw8e0T4jkabHSxTHpcmg0FGSKVw6milTT+Fr3v
grNT/YA99/MBQhv53CpAXPTA34r131OIuAPxKQA+xnew8AN+UXlGkihp6lqDRx5Irlvc4wM8cs0I
/uu/Br7kEzBaXSo+2K6JErqALD4xhuYZNhOczf6AmnXIwpDejKDUZtCntolg+j8XJz+OgB/+l1yR
TyHoeFu6hEIVmjqv8JZkfyXOTprjsDlQ6EVvh4IPyNaUyLe396KjXb+b0nh8S2FvVSF7Gmimc6f9
yTCQKUwiLLMD+2j5JIlfIbr5X4Yfu31GKRmHeADBR1Fm7F0f4ZHId6e2R/sG6cyV+zRkZvaAjLST
3UO/Kd85B+8YKGSivMglYqkeInjzA4W3XOnhbZgHgIpLQ2e79grWmxtwtnDcgbyMYI9Bm994J85c
I3P/fv7irWnN8QXC02JVXkmf/BRsdFXp8gSYc0+WjLQglc+/4ylMNC67XgLnuDNsgQpepFr2MnIx
F4sgp+4kkIblAb26MVFWcPIHdli4iE6cVl30iOV9tGBNkk5LbvA49sKsqhwHESAMgGKVbSx/XHAr
0nadexTel2aL6HJXwGm0l3Ob7MqdX8PHOZEdMs+rmQDbHsF33pDjINpJvZg97gz70F0vrxXoAAb9
RH/J+fewNi3NmkHct6kki+gWPwqiKNESfSg852bgcluqSFBs/G8iKEuju6v8lgkig2yyWmQKyGly
+Cawo5HZ2vvU3nuypSFeuvuwM2AJmqeegl2UbNk+0lHjaMFdCMvvd8LTwScItjyqtvBmKUpE1UUo
rHj/aadAjqbxH7/68NLpMGJsEcKs0wkpN7NJBaG4Xy0H5eVvs/GFjxyoy4MHV0SD4jFaaOoxUfKV
U1zW/M/izyc5gvF9HzE762FHZC0kjc4Ni8uA23CUKbMW2wRK5fvqfEdahhGl+A09wUxpmG3uGd0N
czVSDwWvlv9yxqhhPsD2ruDDL71CWzwmIvl43vA4NHD4qrfUyRiQkliWee04buRTCvwJYDP2ZJHP
rX8AcxWAvxFG3kM1RARzVEsRb1RE7llJ5J1/JlLj6profCeucRZvjghfaYpVfHslPtH6ALpfzuzR
WfM/sKaAdj2yMNT9ohncp4KVyKIkoZ46CZuH4EwcCWdiGYdXElHSakaaBBI/RlSNrzPh0kp/I+Fk
VoJoWHyML8W6E5CJDuYQsVvD0kEon3IwCiBUExtUi6pPGY0yVljAZLqb0JN9QIw/3fse6ebWyZrc
6vcL9pKeegis5TXSeGFrpGa2mo0+q5T7PIjI4YPYeDJM0GaOLkP3NcuLtEdR8teOSNb9TWe9BdC2
8dvHEFzoHeGYrPMg1uwNGNKtLz9cq5kLKiIyYx7cvNi6dwYuTCgd2AapIx9EzkgtGHrSVhSs42LI
zwAb4CSzA61j+nbbYouPoNImVxgtRh8rIDzohluSdeA0gHFL4HLZ/MH+UGdNorzEpUFcIAj402fI
mrlOErMqhoHH/iqBdGH/PJplQ4UjAWxms9PT63JAqp06xHddfT9htys7zg9VElL0lDKjNyL6YqPq
xAYXgGPjy8LpvGxQKi1qGiJvZcZLaDuTuhnDBJJ4PCnB/re+rs1pPr8T0B+LP+0D3CEkjdpSIXz6
EM4Qq2yo435+STlMQ5Ag2hyr35xHX61dswj9JuBC6MFdVlkCMEsAr8ykMjYSql4+1pOTIxi9XvjR
IVqEXINq81AT7vww71h5pGW44BAEA7chNXt1id6jhtWTxkBQLIyyZwNMUZ+j/wr3OYrF5ClKphOU
mJA90URTEHH/NdyIfTvV+H9WQRniN7QTK4bfFKvxPeBa/3+/4KlweR5BuRfUSe3PAd32iPm/5cPL
22/AeijucQDzXFl8rjtXdBym8Jf+0zgvHBvowolfQgRtGGOh6B1czYwTVktSw1rEMH0x+gMj6C5L
oISi6zAUSUj36k4SP5CL9PdZOviWRzamZzozvK7Swb2aFr0QHAxEzjW1FI757Bc87/xzZt2oSsCl
HhydoMsfCa8bHsr0eN40TgWear07CxKQwEgewrZ0+bSp29GQlsEBhzWRSK0zHKiVTruxtoLLrfC4
rRyqhXUJ/58qrdWKAIVgdVP6q7fMmv/ah4mv+Xgsglp4ZSsLhNM1RytBhxzn1fQj7XspJuo+chYm
/db5SVY+/h2jdqgK5H7ZFqoR+8q7+i2qyt24eJ5F9QNlD7QTl/Hw7soX6Etrv8I2NgdNdIrj9SHr
rcbM6nS8SbHyMjQpclODDs9Os06635iPa7OoteqykmkRlHcvzPiUT6cWmsnteCFCMkdTybC55ymO
2uIf35aJVbyW5tQXnwXHPxhP8lPbY3ceONkinE32y3mGs7n3/PeFtVBdmGLu7Uuj3gQILxjGmBh4
v7EVOtO4lYIx3IAD0lvARogmnuVcFKS9rolg1+kyXt4TSM1UCxhIsJYZO2XFD2eLQLXzS1c5+fpr
5vjOtbR2FCTB2YJARDgOUSyTcuGYc/GH8+Yckc0uh3xYBh5fX0P0gbdFVjCEgT/nxFhnR4eHWBdB
gIFZ202qhaCNUg4E4rsH6QEleFyRwgZoWHvHvqXSxxyleEyWdvxNyIvryUF9Txuj7LJGY9MfrnVK
7wmOOH6YIp11z+1u7WEaWNlOtHNUW4B/eOL8n2k3KMR6X8W+CfiqDi+DSYQI0ut4D3AakBsL9rSc
h2Non6QGhV3iHEWlaG2YT9gC+z9AFPwMqK6W3oqGlCC3PVmyhe3+u0zYRoffADSyEOEH46+ku5Ho
VUW4eM2HROAAQGglYoP0rpc5+7myNbicsj76UQJjFj3XIoyQzU8EIWjCVywVB5Vt/TYhUxkkCN2P
VkdEiews24/sm+9ziNr58nfXnbEM9dBlTRkZecQV8UvLGdKXJAtKTEFOKYlHSuGku/5lt5ne2XJZ
tjtfItFLup8b0xrr5b+1Yrieqne0VGZOyZvMk0/UiuKBl+k8quNDRe0eKM0IzNIGrq21DaJx8BsC
3WvTmuXAgh2H5hkdqi1AlBLuGC4wvDgWcIPt6mhOZzgazuEm9Br/j7hUxXgfvlOS+Y0nJL4H9V+0
2mgJ702jrVjSvHZsdjEozaeLG5RSSPr3Q0QyqHOiE8BeouNRhSi+5WKqk/34mxcXuvkl4LQZ8scF
NuEH4R4dzWdxi9XQxerjhrLXm0S64RG5gO9sgGKfEZxiswZ8DwQZiLSDOXc0INU05x47n9B3Ujw7
kDHpazOM7eIAmTxecxBwiSJoRoXzPZQX+9b3nsyW9Hcokf++fJ54KtE6zZ9IX0jjDYRPIssquDEL
AVEk84sMQxj31jmFQ8xLjlUc5Bpv0faN+ubGbaGmP/8cp//1aE0wjehiEQTgX10vbxcz/TUd9QNc
GQRR70p1MStjxAWNTxHyuMq2sjUMLxluedXxCqoILdyAygPtDPF7ysSxqxcreqeVeTaI9YOYhN19
WMqsv5/FdB6r6NVxrvVsV4aHL1xEIHwuB//nwQ3pdmV9H/Dm0X2s1e4hgSOcFeSEzkIS386EHJbj
7L9L9eeFEdQrNCz43vaI2DMtaaa/JnDa+IT70L3UFQwUxLrEWbpq8PG1Vw2qFfTzkx1UiBMyMLAU
5ZERrFUrqPfC3DwnQPiAU9CXoItsYqWvRGfTRdtOGgFj+Xe+OVN6ZD2ScUIWFT9Yu9MvTsGJUjhw
vUj7HOy0JoAdkPRjmlMqE1tj/TXS6dx56DyGZvEf7PhpM+rsUKRmyfLlGPQGqZE9K7sYjGzxpF7s
b7IF1KSVGlyo8lanHQ6VJqgOvzZenOxQ1qn6BOzTjIEJkiLxlF8eg6Ku4nvnxFQhTVa7Oj58We0Y
lg3rir5x5QXw61KwJglmUja+NOYe03nCrgA0w/cv0UyB4ImEW5IEFWqHa727QruLuI0SvQETIMcq
/ipp3nd674nVpkmuzOT0TrsQNf2DtviUOsARujmxa/qBTaIILwDON2EZRD5m6ZOcg/tqooce+bGl
YqDyxf9XOgv9XHXSyp2E2CcTSNuoT6ogmrDS+k682ea+05GVC1dFgLC+aXHnE089tjux5qVVJIVz
UOvJ+ptgNm8132dUspSZ3ve46/J87E3i3y8TFiyJaFCHIdB9MACcxHM5tdVoHxtNEvWmlQopmQ15
lEl9Q0gar9UpHB3fP8cGnbCbWGjI1i50NdqxHtQw7vLTFgZE0cXI4hqA9MK3TARcVavcHN3IGdNn
VKrQX5oaNT0JobMbFtgOZd+B3HIvH+Z1NzefcBh01acbtPIy1p5hRfkejuJo9PdTsAEeDv4CJV4G
Y/EZpj2gFT/Saxd3fqcinAtaUlDpDCD8WbhqHmefgdHFmh3IzU/FTimgEf47sJ/PfLUm6kVOlHhq
mQ0iZOwo2iv7xEgdT0/EO7ZSHPSi9lE6d+Uyc019UfzTxN+Vre7Ui9UON0CU6MAq/rVZ00V+h8+k
B4thGzVKJz+iz34/pk1ySctyYVuot/fS1v8ZXR1RCt3lVJzdzHCfZWCjhQfE7fkUUkatXgmVAD5i
oFM7b7DgCzBAHO1wcSLjsGvZt2Edveo37bJok2tG3rzhEPZjtpEsidGulMgQDUsP6ridF0nk+neU
Ia2TrifVofH+uMVf+MWIMBvA0PE1HQw/VAYe65DOgpK9fkUVV1UayCvydobFx+El1n9UnsqAvZGv
taHCmdtYhpxNYNITt/GoOlUM4mSAP411LVQHpH/DpvXey3cB/oNZAXohIghPAJ3DuqP1cSouOAmz
SENXQN+UwXN94aPQW9iddn9Jgt5mnRLs6n/OcHBqyz28OdN8C5p3cHSrFgz2TOXIqxsP1pYOnxD3
4bIiYSK9eogmmm6NQOombKZ/f7xAxj4zJwkco27rhzwknO9vRQoqYEQTKjwuwsU9fm7Dctql8i4S
sRMz2mpfPICqAOqoriJ3sLhFkXWD1aplPTuiRe1WaLfRRM1Aetid/ZeHV0LRHBh5s4yFZ4qjdEEE
u9KbJepHArJMWpzFPcelFaQxPG2TkH6/zKDjNvMEgGRKD0Z34xdwSKVGG9ZDhWLWCQy+aC2+jAme
7bw2knNqQCjEvaiKqiGJhluiOKvVEmx2ckdNMxsD/hzRqNUGPr0CsFr0Koe9IMup9qxP7OUeoNx4
zqFKBOXs30zJxdXpiI2rKxCp78sbI6M08D5SgVps5TVKaRAoxr9GDGpl628LuhvvF5tKCCK/Aouz
LsgfWse1zr+ehEPefMYiVp8lqcLP97RAoHK+HSp4BiQ7XwnVNUd5ZBY1C39hp7G0FROCx3jGYI9h
WZLVkm/2zEDHnW0W1RuipL5AjXr7whLK8fO+5Y2283ih7Cw5uPROb8nh6awQlRc2guL8/t8UD++q
zS7/IB1f5x4GhNF1HWxfb1ViBqk71UBStDgJ8KNEZNCyxG5oajAFUxCTBXkOKFzuqXr40RPIjN4U
II0xyeHolsN2TIQWTOIosq9n9emm29ul5s7FD5NpC2fVHeKFnD4/AaKdDGLqt9UYVOLpZtsB4Wp8
R39mpZ0lXDuQ0fApetjLEN0+NK6oIamf4wRfLFUluL+GvvwMMZa/zPbzRk1F6XB+jtPsBHxzjSPM
tFEkj7PcN59j6vi5v9pjdRKUDeVvnXir19f+A8kJZlY5bejkt5ifz2+xGA5uhwUBVaQKlPFWVuyN
HEL7sZS5C7nGC8j6JcWm2FfUy7L1wMlTEPfoG3NHciVxIzuwKeHc0+Djw93IOrDlRUDvZdqe0Yxg
cuWIhEUFveXo+DcJ7EgOU2nlUHn3C36695LTHBeTZ9uCKV6nTW1fqPIf+De6o1Pz/K/W+YcMK66x
DwzFeQgMfKVCCxqCHTx8Sic+IucnONVfbFsqU4O+Zu/rLV6/RNWKADsa+oqow4vNINGOnNdIxwP9
B6eDb566PBb8V6BHvDMkGFqk9MyyOym5RhVuLPEa1RbJ6OK67jxlnCjDe2QfVDJdcS0F3wSdDvdq
TAUoBfUMS/M+t++dzwQRtEDER8wvTxi60DqVcGKeeeLUq+aa5TaHIbcoJPMmlFrHloX4j+OyApHL
IhnyCIBiBVUJgGXcTPsHlxHYosYSnPlKvYs3YvZa2YKKsD3r6CTrd0kNq+yaVSn0HXT+PUlNRtiO
zbqGcwQ50ZkqUP0RpZ6HodsQXlDi5FDYPU4qnFaRumYFV4hdFz4hEhlCXXKv9EdfnAtB0v9BaQcd
Abi4kMzPBgo7OFG94hgpqqLaqnWVrOHoWarBnxIMNKO0B1Ct7BPK6ftiij7S0hcQr/j/QOxzYbB0
mFxSJEI6NXVfiCB3OvHTcss3ufuK3wCcvxmUsyDxht9TNwhdJePHAY182zLU5d/9mT2R4RfYY+v8
MNU73AxImC4rKhc25m+KZPJqN0EieY/bkLcCeNJQ83OaLPbCLMa21YRBoIXMwYZkGUekCXFj6GVJ
snt3aDOOAZDiEdYJ5gYom/MrZJbyactTclT56rgwvxU1PFYaSNsW1Smkau9FXLmQZEFSlGMKANTq
uFryRcU+c7gPevKC0rU3OPn7V+zKYKozQbCvnYaPgoImaGVGuYB0WMhhyeo/XIAu4EVEY1oeitwY
Su0yG+ct8YEuDqX4NTJeDG7bZ1niGngZRus7QlV48y04nKBqZXZpxE+uZ9TxcLPiHWJ66WCkUWzD
YcalNCjErVG9B53hwPajYoEPJLMS96jhm9bF0CO5Kwdm6lojdKIo97UFHVnFTSMKYHWCcLJySrfM
21ZUckDaiU1EEq5SjstGEtyuj4rf90PB4qTt5g3zCfStyh181uxxY1vQsWk7N751ii1tFEYRBbD9
48VSh7eocLBjOwJOAr3x5yHEvR3Du//k5EtgRvnaIHbACucwJwxtxMogAbh/cbnV4zG9RITFi9c1
bhg+CD5np+GW+8kTP91er7BKzp2NSIL7kcxTo/9u3EgKH51xeuoZZLHgcoQRDVZWOwKy7c3xZKst
WkpsWbjydLIVWfgGOCnVP5sD/ePAr8xVRI0Ar+j3mTj39TLC8/yHOLE/ypgmvJcbdgdELsA0Aj4j
S221/S8kzTtLGOcvpPai7OJnOlKJaKKTJNik3qiVoCIys4DYzzQoNCq+TKwxs6864qguwbnqBCbK
al4b5c05zv7QCIInOjKdRt8zQKErg2PB9rCTDSdm62dkSxU0E2YoTVuf2ySznsyrG862n11Y+OGQ
YTGZmbZQgWrvL+TZX2cUNZ2EeJZtMBmyJK67e/MhJPFRxlBeB7AaaNa188FMPtauyLb2v2SMVvJe
yvcdAECo25AKJ93BwJzGOrxmDwKAokUaJTMqYS79dW+ZvTbzYcEoxh9/HoPz+4OdLSFYBm6GrvpX
E9rqxVNBia/hSnAtAnIcDwDcvSTfgO6q59RQ1ENmCSxOEJMDhy9EsDLh/ERvbuX5KrxtUL64aIP9
nnLNCfM45mjj+Z2jOjvwsrro89oa2VjFvBDA/cZ/oJrwm8dPbSFReYfDpuK2nL7mOVD3yfNE4/c4
88d7g3FcCLv/or+7giCh6O9RatLhob9lr8FiHk4wXvFRFnIK8yAD1w1Nora8HDh1qMt+IEYtRsAc
HOAZK9PDXrklaXIZQ1DpTAj215Q8vFBQbeRoUGiHHrUI/4TqUZXn2+Pvsk/0k+IsG4ih33cTul+f
roF7KDmzV1HPk6yDZdTNWj16ue9HWyG4cZSZxZUOoTIkdYiWWF4iU1p8pA39lgM64Y3GpLJL8/xQ
/eOjLMpw0gGzNia6h1dDQSJuYG7h1NwB1e4T/z0QEjtHLOxCqikt7lkn8YKOQUOrPCjoX9lnelYr
uuWinCSCVqS+ZmSrNdVfUG9CQqtQnCI2ucaJdU2WyylF2qKfHrzkKt2yQgTpTg84Cew3yIPbiAMC
9nslr3NXecUSj/ty/WXoSCL5CULKEfwOsyTaVKDB9UncyS3RYfX4kkrBtR6qh4Rwd9eAcAQ3izcT
GnOTvgZ4HuZw94DelrmpfxG/JzyxS3pKPAeoTdE7WVraMUif9QDwxo55jTLi0znkX1YU33c2+iXy
sn3/Zunp+sZLdUL+Ytqo1c9/tOV1QMRtkRuNxB9K/tgdntQ21T5InWj9kQG5Jf4KsfmcchfEMJCu
bZGllDYpmS5fJ2SHtX1nuNJ120Nif/SJCkl8VXzBGhV3I8YMMjhTkmA6y/rQpNjZTVq0FRiuSsXW
ku4sLlZzRVBj8ucF1UjHXYYxmWqdNF+2f5RAqvfoJuTep61NKYME9LqGWP1EgF4zvq4TDEl8tABN
4cQlEk0n8nDaGf88XQYcHLif7oMf/mlRsnCsNVnYx7YhZbIpGhFCP8OofHzpYkcQkIY5qb1wmDgQ
d+ZUz6M9u4sRzRR7klNq/xiNvCrN7dnrCln//AAcHC+o3fv9M2zBOib6EKJ/JkVraQmax4cfwfhW
Lw6UXHVA8HOYMiUvydAagwwRuJO5gTLgcHBbg4cmpgzy9TDHlXVgH9inFXVHdBqYfrjX7Vv9uD7N
1WYS05n6Q+LfvoFw8ZfJfEursjsqf6X6jw6kDMvDDC4A4JdcAf3IaLfMgbyXq4BauzCP9RaZAOwc
c+a0R5tK+CCWjY/bvzfF9rLaWpVUz4wj8oG+ya8uDVew+5VyvSx0Mtn7Px7m60O1EUgeD5MNq1lL
Xkgsj+gp/8jaE6cNjR/kgSRk4HW0IlSP+6sUjqWhoOIJHrYFcF3DSQS/3AjfvokycStcdEb+cm83
BAoPeotoPVSoHPKufqVzkubQxYphGw4OA7+Ssyl3/fKAs8EqQRu2KICt/row19IYby4s9682sOJp
fa2QVOaI9yAxeskWGT9L1mp9BHLJkQWuPe99lLq6CGB194LQSbVE0sDvvBCyiut3EYLrmUm31Zsg
RuBEoZ2XOUJ0H87toIx3ErpvocgebEQdA4tYD2AJREsOurJTk5/02glXzOVPRZk0QgNzVgIrcWjG
/ftMzfHjNNfYlmTkNO4tYGWdsR0r1jcA2qt2my+uGagv9FtrvoQW4d80yKHzCy8eEdV0LOJfWnqj
u303WJZZi9USOiS/5Xjp93GOQM2MP3WDDbLXccDdQi3cFkyigl26xBJelqdnkscYUg4TK0cnVfoa
xewBHo/neKdZJ7sknkMdL59ICb2exWD+Qeu9DA5GMN8WYe6Vnqv5mq+O7RW3bYJDFzOFwjSqUFJn
ZYFk85cOjV9W3wE3bd1D/ysqpNe6iCXCFnq/d6XUKhqpRvQVcYIJgoY2pvhvy5U/ti1SnRNg5lu/
B3PprXtcfqv2JnJtlz3ybNVDb9uQUNuSOmqPIXytNeRwLZS8K9ESARbzxmUC9mSY+UVH1ly57suP
rCZxk1ngGDhCDcV5UkxLRMvhe9XOgYlNnqIUyOe9pMEGW6n3mHGxr6pGGLHXs6fcaGacRawrY7aO
3rKPIEsu51lp8jZ3PUz0DVCTmL3uhmDY0TPEX13eT+1a4fpE54sF5JSus0FAHI8WxoLw5xjC/yaE
yF/OfnRM7WSR/4sIkAVorUQ3Ju2f4D6gYy0HPTkR2v4RT+/cpXJgFyCRB6NWomqCYkInnAEcl8gC
LH9fNK0vFOu2plU+017jXDr5ajG9YAFY3ss+G4rjTOYEwxEVrD/SZ4pDZfoRXJl/2qjT3+nrQaqJ
mBhp0js325taaib5e1E5ZvE8d19u0Ald/zRyljXRTqu3nubhfiYAw3gbj4GNcN5WbZc+JUGSZKzW
02BKGEw6KRmEKUsyaMV0cNYdFf+3H2mKJFQI6CdFeGcyP+g2LeQwXW0A1l6IVTNKpjBCAhbIrDDI
Yq+mOodtPaBFmCgworYSLaUo3UJbiMx7xcrexQjy3EEXUIA3kDlYTVpXi3qT4+79aY3czfN0edlT
ijRNXcLX0YAb747y8ioIttfT4qx6U8AoSBdukhAa3fzxMcu05FJV//O2BtCMMoj4RHNp6Ye1Zleo
hmnClEk7RNy0QaeTiOt18yMLG+TYvgwDgIBK5WUNPB4iFMryb3nNpje9DXNmhY5IWi3Wdqn1CgU2
LTm6MX6en5TGVP/Pt863nD+yJkxGC7zg24mpLZ+YnvSa0qS34hzEO/NpXikIbl22XW3xSrK+FD1H
s62DBTekMxCVfUnTNFAKDB0lbwlcdo5Sp9qDCIXbpf0TBnD4Edp7l4c8Ce2CHPnhhOzrLRkVq7Uh
NhRgg7bi1QBtLT/kGDPo0mR7aPaUWhmmE1a+s6F5bNGWrQzMgjHeW0qimQVgdgPH6y83B8sWrvBZ
uVitThOyNas4HdYXuaXx/ZU8YQJmtJg+gGYmV1jLCvBspBxs9310oXfw9KJF1gA346j++pOs5fdG
wubOowIoMP146jtUAhwpMd8VgIwnhmqa4GAn1v5OWwwYQ41g3ACzy24tv9mSGJhDsFiyxTJZKorS
YdPbENgP9r0QVPpJbaDpz/Fy1t3ooGVUczN167ZZyT/D1UIbpS3qP9D9vo6v8Aiy/MxV1Mjm9PZ6
rqYwNZxk60mEg4Elu2Ew1EiH59XZhEsMI234pYFepvVdxCkI3eG5Pl+jzcirkgfUyAhioO1egnOq
/xUB2ze8HW4PmAP9NC6WjQ6OJS01Igin6nwXJrHz0tbV9jl9DhEDFbD1u9LdlYcaZaNYlnv8qYVs
Y/vh4CQOFohjl1x26rHKGkWruYoYHfc5uyER7KTX8dr2p6Wlo35MdPuQdBdGwlFhpLOkf5C4FbYV
9l5O2WP43E3OdFBBoSMkm9Ou83OwoKscD9RBzMjD6w5Nfm0zpQqywYpwPK39No4AKgOXDD5qX8Y3
TH/T5jBkU0OVCDu8mZ4fShpC2GkU577A/h7suS8pRVj1igFYGblSsvPli9fGh3AowMfVpEdGf1TY
VQTk5vceFmVf79aKHJaT39KW0K1FgF3CTby5NRmNO2LpBYZnOY5NcJF0jUhNXr2vKJHJw/qom5rC
cNmsG7IWfbka9vdrZAaZrGBv53qUkUpPyKhuuY5YgXngag+lhm+yxiB58xolLn6CjFVX9b5zAxmP
w0ktT2dMU601e9yeGnVB8aLOMMW2neXjXsgpcuENiuvcb+rTq0prh9ihTcdCMo+pQJiQBf6IN0AT
5sR+AYn5bExt2lHfg5c5KcBJc56EVlZFEVmR+ugAlWYa4iYY1Abrjif47eSusfh/eCKFyO13l6Gk
OeZuOtSO692RaWUDiv4eZQHm1jx79zTfc4ZJeVk2aX8fVXYjWpTS70SDXZmMjXBxfhUljR9h03pj
pgbNLGtbkOyll+gQ94YuvFeZHufWPcvMxqencezrb7JGHdERyOHSHCNpImDPBzcIk6Xh1fzYdbey
ANKypsQ68CwRpQC8uI/4+NcGvkZPh3yUM3n78mpwdMal6LBWANhgvx/u0dc/f3NcvOlcOx8BOgsw
SWvBZeL4QJLrRVzLDGBL2Swr26zPV7EgqTTe1x2kcQaS/PZfe9xu6Z5fY7q3v66EJz1EPtzOu4ev
OTR2zGEMbn6NoLofAKgrjdhBZDlaeq3GowjATg7/jSFCuL6rAd17FudcW1wXrvOxPGdagrpjoWKf
4vlZFQvJK5bkhGIHYBZM8VLm4mUzGVTR+QorT5XK0Eh/85UH99RRzBTSjiX+N7oqGtZIR8o79wdb
Q6ZMcPm70PlDZIeqxvJKesRscwq7Jj/kRmhkde3BNbGtNggl3F/kLGJtjnEuPPp0B7CTHLWFy4wd
THMxgNk16AdvulwjElFfZCMmVzEW4DyrgGvzI+WOgW0OV+3SAG9RP5l/yhiZC7RTYtg8jNKEXbdC
XKPJrBK6uMhIW0TC5MOukXY7go+EVuieJRrbakR+xy8K1he7ssBzXmfG0oPn5vpMhWWNXhT+o2cO
rEpuMUd1mBifq1vVrcqHKTHVVjxWAQ3B/y/sE6bkRY3+Bvz3AM9gfAcHeLEqmA3CV5AyWRqhxQHE
UmUPnich9IWRxvDsvN4i3JfPkQL7HXibQvjL7B4Et00LXHxTYQ2p+VgAIDYu54gOW0bEkkwA6jDa
QtWhc9juJcCOGfGG/ZQR3KhQeXc+hrco3rw2aR1KoX0Mf5l7lAsOL4HLNwYhOCpff1JE3x5aA8Gr
9EuBpHadp2uowlgZ2eGRiig0edRkrreJNOVu6SXUlUECPTH16EqOX6QvEf+GfqrzWTpady3D1Nns
Ak0CBNvnrB3kRB50lLOOieqDQT4hQSHYQrnY0A1DoWpbV90mnfYs80FdzS1KACc7bMnZvpAW++W8
GUbwGKEDJ86fk5x3f9AaiaQaG6k6M528aBax40xp9TosO0sFnnPrkHD74lf9M5T+HR5ho16g7ryJ
WNnmdFRkAOQMBQpJQ+xlzuq5YiLOaa/JveMuqT0/hrjc4pzCIWclgvtvjTjr2QqRrGKaMxbdsuKG
zLsQYyg7zeKgWtHPpwyz1f0ujQ49ay7jxKxOntit/rXyrCKZ5BbnfBGSFlOlBlEDhI4a1Nfc75jo
ceyZ0VnkcBbzPfi4eza/g6/wwYNKfZJzQO2ODnjCAIpKSovekpgnMt/5Q73DgcnAFTtPniVuXXsu
mG7BTOjxYj2woKmEZ5A2cCR1Y2k1JjoqhTPNIKBZIgtiy9a6xPCdOtmbjN1tN+NQUx6IMBtjpUGB
WxBwhduY2IKwy2tWXgxX222hNfHsNHBrry4jC32SjsISJSvnGW4vHjj5bk9+jRD9CNv1tYwNAlIp
zv89OgVjAwoh3fsTCJaQJFyIoqpb/5yEzxgO9pHW1tpRmm+h+aWdjhwVQ4DlukerRtjdYN58q6J1
5Iojkl2ZDGaZkW1hlFmad0HqjSuMEtpxKUUe8GsAxVftt1gY2sH8oc+/lj9NZ/NAibt83g2lKlBt
s+jj/SvP0hBXKzCzhMuUK0J007FlW4AkQKySaB4+BIcihP02iegQS11LKtAZCIFZ+1TipaifICrN
rpijczBGXPHjGCIWtx1vlKU+DCIMzvc+6jRUUjuWpzNS00vIgfVhKnYQJQZuTun6pIPeH6rn2700
cFqc8MsRQhLeyfjFtnvqqGXg1UFq8N0O/tbTxH8r0Ir+pT03BAQFjzfKBpSdzKdhCv94v9Yyy/s0
t0TwzM/wmHxM0LRGs+4ztNJV8KgBi6/xWTo7IUtbe87CozEmqvel0JLk3FQz9sZT6nzD7p5RfdvE
0xerHG11sJxrqHGmr3SdiQHj/R9D4tPn8MTdFr6sMt0tKC8XVGy0ulFqa1PD+74Lj/9BFpLzPRv6
s2qq217eCZbyrERgNlrOJ8l5hPtbIux3Jh0YCLx93LpclFHdM1/yJQ438BP4GxEiamvFrPaxDepe
7sI3AosMaTjk6ntB/jv0ZeOfOzqeW3qHxBXRfwV1A93zYqJkahN+gjQtBXeqRTXV7ctGrDSMpHcO
jGDz355shmpShwaViy5KdmiBtFwdOahReuiVLqKPktga0hh7rtQ9QavuiSxeOq+3Dxhm+SRkbzJ9
oQyEVQtknkvY2ZG05kyuP/Nh+tttRjcbDrFruIzJenqmD00AjWgYxsGoPrL6r3N3ayhxvEKS/2d7
BZfgB99xrHrjrYP2hi8FLcn2MvqX7rlo5pQTnpxTgMpKuGFQg4HRqksQUdKT/5/AN9GKeJUJ4BqT
1bJ3Q1KeyoiXnxrXRNDyPR6fQX18ENQ6ZFUP4O1Fu8hpZkvwOiVzB3NZoS/PU/YqLnNaP04ewpt2
/ghtVzVDeAfoDw3fcTyHdN1gI+qM6txaQVTjpELHewd/2Ny1YvgjBpmGWDsEnthGeA8mnoD26c2b
H/S+03y+6talk76BzxLRQju9lHssNzB2oVCU0gcS4RjX8YCS2LDktaU1RhbIEYa87SNWw06aZYrs
aiyjFbthsJtX7tzGCFzw/mlD3V5Iyb7SppIz26I/YQQ903zcRex21tgGYfUrD0zrtkTjGQv3oQks
gfWnTaTcW91DINFqEaO5T/4EI3TigbbS8ZXPydUGNszq/hQReXZ5mNpGjth95nrodYF/ksmq9BMr
kmYBU88D78SQXoCUtKRxYBf3v9vmvGnp1EQpBHY5Omt5U+DyV2VsHL/vOH2WPzP13pNANixinQhz
6IKXAXQIIeWVCAXwTt5nRDHqULqbnaU/L/J1WmqedRfWXDS9I1YtUjYtc0ZI62V/hsmN0t2RGTAh
ZoQSAuH9XVuuWro/QiY6rsclKdBIfiDYLsyONtDrDN0MRKkhBOyj4AgquWTT0h0gno+xiP28p8FS
q27xS5jX8hn76zYEu5yEEu53qNhdZ2SKPYVtFpgBblsuBfiB6q7QJfPXUjcVZXHLIM5viWZR8bYN
1I7pBxlJ3he6cT2rwHp3DWdk4ubuc4x4H1iQizqC+SRMLjHtR9zxijAEpXTbDl8NXB5atJkdXrog
yXC5OQrTd9bsFUgDwqJgXpnk2FamGT8sMbSwQXEen/wWzdLzxCKiLmpRw7i+mAvc+dUXyyPyHjOq
SvqXOD3HLNvPm43egYx0Kjg8KOfuSTbSIKV0WTEOeWTwVKwQhRkZKCKATiTR8eK+3CsKy7gr1Lpk
Z5NXSRsltju8j060/dJiwnJuxshasxxOjDwYoTmadAoAGU0t//BJaqX5fLo3glqR+YyN6Q1pSKBq
0ZDA5tXyCO+ScZZesRPzbNUwxCdNO3+JuIp+8gFjP4/7piYY2nyxsAEfiE3ELEHZIa3rImvTajlc
G6eYZX12WwlNFsp3I7jTVaT8dPMYFB9j2762J12HU2gP2kLwSGfUztSRaz9dXf45m9C73/MEYvsj
BVQNNhSmer2HPppn0KJvYV8SPth5pHndvaULT4aAv8dvMLFbvzQ0ePCb+g8WoFwx0msH3eSrxgCn
lBstNYuyRnkCZx1Zkh5C5U8pHMqBvXexldXxUm1g1hXBMviMVJp9aNdym7sqY5XE0cbiGikew3HT
thIBr3Gw38GoYrvXhFS0Ue4e1NXJbX/5BoW9jlHwNxJeuAx0s6mTU5BcgQsf7dT2RdMP4/phMEff
xc3uLj55JD9JDittILq0ayhUJxPlB99S7mp3tPUcNI5CsP+24JZorcz/G1C1EpVhR1Vsvght/uP3
QKTQOXU/rwvBVHZe3jZn4rYOZzLC3xE8PhKk6lb+WRaV7rrvNLvdgb0DaLKhiu3z8kcZcpdk8wEM
8RpicYOo36AygaGMHcpV1saRV3fVxI5fjWMJ2HGmGU8Ink4MEXt9S9ErQLij3BNSgS0hh+EGVyg2
GMvrC4TXMs9vgAyckWNZ0luwcR0tBy6S0gKOf3XsV8skC//olWiNOpXbTh9hLvM7ELuDNBBzrhf9
ExGZRgb0tuU/THETuAowfhqKFyywl+1nTZfCHK4VzBiz4Pq/M7PtHWZpo2uLbm/6OGpnioK91e0+
yJPcOCWr1fbWAdEVtK7vyegze6FcTccAcndMCOcMieariBh8FcCRs0IsrvbGrdrm4vqs0tuvld65
4JHLECfcyECISOL7MKGrLVXJs8/md1x7xmP+T3zdIiPXc3qTwLJU1Y2AHTADXicz8FajhMYzvxtK
q1i4v7fJ6pD6PuaDF7TpVlz3ZKNblgRbxj1nZxAZUkTWIRm8kUzpwhpXv7xHj1tR7pxKFIW2jJTM
/VDmzv3ZnFYAzHFPMvqQs/PLahBL2M+2+WiOI/8gtB5Xv4erYnSV3Jy1xXi/qYj2karkoUNeoBvx
XRsnJzsMA1UyVC+TsiBcdpj0lZv7o7LKhI79DU+OSXMKm91CZw2eqTgcNWQR+QZb3DbOvMUhSU+m
O69ctIDfhRBmmv56/1awRbs91//MtRHx9SbO4n4Jqlpl24zNn5pd7q+lvi6VFl1TlIzf9uxnriFQ
m2R9ZfEpJrD5IJ/KQbiRlvpiCsfGLIj0KwEio/79Lu9Mo7JnBhU3bPj06Wos5NF6UT8tPBKYBxlV
f/FslQ0umKK5yXIupC+64NeTdoLyfOI76qmX8gmNKiwV6hIsUJzAYD8/lkXmW3rTdoEqhL92MJvq
9jsrI76KJhVGSOhLrj06plZQ9yHNuj21RyihTTKHeyZnsaY6RRjd/BhovuLCgkol522v0vKS5Zvo
4FL1FCzr/dgIMIJagDjaXWR2a/AG9IbIcIzmBskkb+dO3oooWu7W+cAAOUXEsK0iC7raGQrNIqWf
M/fchxh9TipE9g3pskJtD2gFGM3tzNSgHcnoVVwy4LMXIVjE/B+HaBBUA00CMGTlzwoSIrVyoZmN
FCCHIUlw0WiSAvP1dvkopIGkyPByILtBjsi7cS5CIRkdQToZ8tUOd1kuPamBfqgksbVu7oOcffNK
/PjkbPjHoyRI6WnAPKBEfZt5kuRJqfgHVVTSAxnZg2b8A5z17U/wzwd3aR4R/3Q/X7Ltongbn9Dz
THAGYcXTstjCLCOdyZg5AwNRCM02DL95QqpmBsNAQQGbKOCB4eJd9t4qETFXcCuFcRJGXBjq1UR9
96Qq01/5/rclT9csbESYMth5aGDVj72vVz6am0L6YDJCEF1yG272auJ/yFftbsT5mW1f5Jo2cRY5
QeCgkxvkI4sKAfzXLar6VHOxFgT45wl5hz/UOF3a+9r/v5sUY5oT7unvDU3Ne6PMdkEFjlEanP3g
1UCffd2jJKx3yit3OKJc32zkYJltbXiZZ1T16ygyUhfaVg+0t6PW3T5n5JDZKyEFs3927yVtBxR/
+2Vpljcw9OWouI9qfwICvDfTbnEDG7lV0zZ18xmnTcVi3+oRwdCet6ZOXiPMwVjCrV1+kJaxTqAh
4Gy0hMyhYhIJ8MkBhBXw9Vmu1aJpExG5Rq0sckC894ZGd3jXj5HY5Wv5nDMbjX8yxydK0NuUU4Kq
wm3m9SJdx3BE92j7hh6wagszDo0mXiJEGc2cepLIdFgJd+TZ6gxtv2YaL7nVBhvQchhl5voigh2h
c6k2cYpzZiOsYNK73CTUmiG7GiRhUomuK/CMzKY6VKvoduD+yfEjxDJN1sbp10GTYWAzwBzSOwEQ
4RF6WBae0FrJMO1So/5KA7R/MzkSGGgcrRc9n3YWLLuH1xlT9R46UGVAVWDAHIKfdY8xrGFsC7na
7eomzewtWpbUscBl2DoGXoLdfpXa6jO5GZCV/M3kkniUgg4rKlvZGbQPZ/gnlU0JMVs7JKGfeT51
HN/TXRoGgpr2fSUCtvEPikqwRa0HgYS9geYyNb8Zh1kstmplajQ2wHq3+5l8cyB3k9FbBckGnbT6
GRdrlSp27UmCXS/mfPAtAc0rA6L0wFubMlfImxm73FRJDEJfEwdU57MyjQ2hDfg2txhh3Gp2hgy1
v+eqoBMJKe+CRIciYJbUbaZTTlhRFKhtFIvLO0vAvgGHc845G1InM3H3scPCfkyEioEUlMkDiQkn
S/cPKHK/6C0F5br5oadYTfDm5sy2LQaTpVNyOnN2YMBj8A7VkiA6/6JqV3XWCYm59LWMBxuRaeWO
kKScvuANjw6dj1kMevSAOVmqoBY5kzfXIm3Hy+4pe50nhw9Lp31jZKNOomJKAznf7mei3q84jNKp
cYyEBInPJa0JPoyl9u4dEKj81vAWdpbAm0vdkbevY0oXZhSFYHu6VvJzCGSaZWQxMjn6/Uod2Eh5
7C5B+9cxYEfrcWJejdamRYHU4IY34+1eH4Puyw3Hcdk8mOO5PKO6oo35Nku/sn99CfBKZPnkBZjn
WsOhwE490QdYAkZ3cuJwlrp0TOj6PCGU6lC/g0oq/jse5st7LSBhlM60iVMnm+CIzgoVEdBmgWe5
PSMIRtHDQmcOAIN8i6FrOlRqs7PVk4Jpv+YtvwK1WohMQiweAu/8AzwhzqKJrUeLIdwvOSXE4Ytt
gpDSatzkWUX5RhjUlsqLO/nmTzjxpoDh7MgL56EU9VGrRi51FadlDh9ih5TDxefTLEY56ZgFxsPZ
WT5KJod8TdRT7ZxFNnF+Zt/Dc5imUP3mYj+vl8C0qgrUfb66Bc3HRXkoD1kvF6nJl3k7HTzjeYll
6gfELWEhGdcfjPEWQ3cuzspy5wlKkscW1f49wf6UsRQtOQoqHylAiKaHArrF6ti8cMpewfUzwBmY
WfWYc8IXky6VTrLqV3sOp+R343wkrPr/EwVAdRg7TWhuwbLYRn0Fy+Az1/5ucfFLVkHVfy6I0CVF
88NhEr3JeKUKZUKlY7BNkIRChPCObz/GaQWynhZOpMyM/612HmhIe20bYurOQbTlKhs/hk4MYUd8
s7wZk+tjAVhb8bYgWZAXLa9kxYEn94juw7+BK+Xm4zl9enugwDheVzgdG4D4mvCjwEkh13t97/2d
dc/67e74wvvE6C+LtgrsQwX3nOr2CvSLci5umKj0lil36FhnbSDcgHdsj4pOv2lyJZUi163fgz0/
F1iEil8JhCpvlNd1OYtdH2txs5e0vemNEh5HbdmuaqgXf4PIkS98IAeY4chvM+jI4KZKnGU1C7Ne
kVsmmoRR5p8zJcYHn9qamUHiNr/foAYHEmH73iBe4YQ/J5VINdo6iRNIf0Zl7+v/UASrXuUoVKMM
9i94XMGKdshPB4ZXE8opm/hEC9/G4fzPKLvef1FU5alMcaz2lFhnOJhr7dHK6h8CgDaItidOSrIV
5jpgeVzumQQ9zf4UbCCm+5tezIJlslTG6B5LJAvaeLu9SN4b2mXDxkmVmTTeGf7c4fp50gDtJcqr
SwrC+nyeJThL2ozQv7U2hjMhw51zlYf3pAbIOqPntyv5cCKfL1QYe3mD25K6liHZ1+KlEv5ZKdJT
qWlaYXbCU/Y+oL1hvtLS/nShf2a+1c0CTTdVfgoZBmA9H3yTqSdfLFvgMAMxFLKXkRU1UGabgbqE
R4AE/5vEFwVnAxcSXnSSPVgrtFvHkBuu9F5EL2d7iqPiD3KsrQi+F4Dkrv+DMvUGbgGHF1yVn9QQ
kDWozh9kXC+KIEYQTMHCFH9S6sGrFEEagOPs3I82ZkFs94dWBB11qaItlyEsEKL14oMF46resMrf
XBAzFJFBV6Wqr61DVV+rlYCGHPI+F1Aq4W5wqYcr0MjKuy05qXJ+Byfa0SDquaBFaIWg/C3HmYAn
E24F+tM0m1Btvxxx0fy0RAvLzvxm9LOSjsSkRojYp2rD9gOaDfyYDwSftsZbjB4WUPmkiaNOqwSI
CRK9Tfuh3X8Sf0DMyBDL7xHP229N0gCRbrab88WirDTVnLG9N+Tei8Bk0AGd9o1cc4bE1828N28B
wyLbArtrKRolJJauuwmE1C5/4hLu/6PDe1bF1tEmgoeDsBHxL9JuhmK+33lJ/uzkRJjm6XvRucOE
qiGU9Des6Mu9b/T8h/F/h8RA4wkMajeesX4IiWITVH8iaRYuE8lpu1AHmXNLPbK6Po5BXNzE7wgk
xrdJ6AjMdaJgL1fbxwp2L2U1cs6e+FL866CIludQdZ5cDYE1aihCuSihucAkEhZykiec2qVcnOh7
dEfnL8/F5ySh1DCYbPJgkP6heJ/l5c7bMd0SeMbosmCQdvtor3SJUWHRVdwUfpbqwZ02bliP9/ex
tWmW3s4bHqX7VWvNaYmam35ohNIgxuJqNGKfU8WVdAYpb2qRHmEIvFe6y2AgBzbcb4QjsMEUiznZ
rzusXFBj5f1CXiGWqYUqWHj6+PtN11lQEzUveCUArn7OLDOc0HiSJtmMuMXZ4Iv0TCLvcp60kQfL
9V4CHUxuomVbIwAPslfO48JoxoXojQwOGbnIgrBCpNWgatjN8BxQaKhboPaLfSYJzIJbklU5mI1D
RQ89juW/9ze2e5R4C46xqRuVrPBpGHXf1ZCSiAO9JsSK4BSrB5KmSNHhGvqSfcBK/bn0MJEjrg4j
7n9ds/MQGcYa+/HJ5ekPzU4A2/CDOWc4XmMW1zk9Spkl3XpUoQsft4gdOsWRSDF9OAUFlMxY6Q39
n8cuQgRddgAyUApnZgqdAiuSXEj5ZG4Ioz1kQjmOTuDEXt64sMSK7kcRo1LOsRxPUoiCM4POMdQI
JIqmASmCiUqFzYmjUvJ2ju86baKs0q3mViAfkALWabiwCsZO8mz9AafoBV2TZudPsQskw0Y8H47E
KSENsdaNHiPwB017bszJ7rJElg7R0raOqYsmRPNt1iVB8T/MFnSq3pwAnXisar7td458phVcA/Gf
Is2JEJ4JNYZ02aROCZm9gMnHtVEDEkX0aAkM1y9N+n2bCAkn7nY5KkkAU1wBhkl6d6x7pFR1ywKE
nZe048pYWPBvore7/6eewMHxJjikGED1dFisRa4wsSk0sMekO67VTP94p/g39vYy06BYgveen4dX
SHCQp5Ki4hiE9AMYktkpLwISr4bd0x5ID4LaG2Djr8s8hpYDNTi5d8PncgBBRAxi7qIJ+h41/w5l
Tmgv+xBAIURdJ6lKXQpdcl/lVD/cPi76Vke1KbBmy09drAHuttTwexaCTwDT9HX6Z6AN5CioNE9I
xi/fakkswsATk18WHlbgS+qkqA0T1RwmjoLhn4VWjckCq+FZ8kcPtbWRkxshbqPYApHAT6tEmvsB
z246bJMliIB1Ei/9qxLb+JiPiN4CqQceTWk+qOtN3icBuPT9/sj0yCfLkzWgE6gaSa06R/Wity0K
DoET4gaMb8n0OTMSNb8pUztFFzTTMiAuyinb9LJEuJXYXJz1ZAbOZvYMlARB/lRSl2TlaJ5pIuwf
PJbNhaleGQaMNPzsKVSexqwSIaUWeYFATLB4+PQH8PvCo8E2xUnT5Z8SLVDU4ZbkQxxPaXK1ydEN
XYdjFogEotgD79Zl6ZBzcMSZD1OtBXu2uHHdflxyTPRrBLRyOa+qfS5JNJVY62o65rUd5k8bIk0d
p0s4vm18Ra79u1PaAR5J8O3/vAACS1LEViFH/eVGWDzBTHY2ptnAC7nT01AFta1ZygLG8xeCZAs3
0gjExbFZcU2crHpfGnMg5zC+gCVzTlrGJA03y09YqFY7bOXUyRLswOx8uQkmBnW4a3gfPGbBE9Fu
oUBg9u6U+YD5FEeNoTHXM3Q0kR58/TOXnaRRCgkVXEFRSCnsKtQ3UeJmysHGXwjB+3vQS39unuDX
uYWZZTYCo0FvB2wREWcBvAkNNwnMDV4HDhJeNeIxJyxYPX+oX31gUT9NzXMiGLP8APJicJ3f7gET
c9rcnzz/uTt0+EmLhvTrnmFphSqNmNvuiOXiyPBX29xbR2o3MskwmZZ4bHItgKQyO/pvY2V60lj3
PTEM2rsl6nhLuleqRA2IA7KZv9HANCEJA2F2UyToYqlu9XbF91OOHELwAeBz028UWbaCjMTSZpev
pPmg+6GSMPN2jPXxTaCTr6e+Hkk2+bA9X0e8/kSnxE7/ET3HGtYUt03SqIDp8jd3ThgwrRwpFR98
4s/+alpYSLPe0bN0BJpoBBmM+nGJaA2rCQ8QeYQ6JIgua9oHaiYen/GzU742keNOl6+K3lSO2gW0
tQWe+CNDaLfye55EampTsbzms8XARNCLxe5MVeTYzA8Q1JJV5T0Frf4NLjaaowEou1eN/XsLYVbU
Gc+R0a7NJkGTgsD5pChjcGSJZqBhW5WALjHwKAamGJuzWQyctNduYkulllGYO44e057IXdDL08rU
znxnkClTpvtRLdbsqL6gLbbfS2nQ/NnHbI2HMsLbMnF+uqMVAAxJkIj1x3sWe/bLKctVEjj0DqyN
o6abZ/t6nVvxjaruXDZXg2RUAYBd+JVpsc0DH0/Ls9iPPsyakmj0TOLJ0mOnguaMBoUQOE49kH6W
Deau9g3Gq3x6FWfHrq6NtGTAxB+5VKAuqKUcxmVdxKn5ulp0mOvKe4ZYK3eld4RM1inI9K/+xV3K
VIG4ckyJ3YXPex8an0hYuqjGo6NQ3wqDT6pVFEIYyxpMH/okktSlMz/LqqeEBIE2KIYjeQ4ZmaH2
F9oTxrF68mwc5B/hPDj0/FFdxNYXUg7ZX0FiW83k1qdbTCJfVeKYlaYFOhlUvkkEyc/EbYeZa5Br
4DOkwtDKToTNd4rck5VbYKX9g9xZilYho6Uc7/4FuR+XBevSGqmMIpb639IPoyjy0T5qEEobXJYE
3+3BnwPBpzSlkO72hzCfMqG/cL14Fdp2suEggy2wUqaBg+hzm83SeCxNpV92RfCH7xt7VziTVqUt
kcw3gDo7dXBeK3fYsrUXsEQ1QuZYDKpJY3+SXcVNa+hAWPcoXqMhW6lYmWY4HCvw83fv32T9Mkj0
Cv7tfgKMqq0PBCxHRrBrS/yO86lVTrCfa8v9LktR7PUG8JQc3cdgEpgmU8102R0D8aR3t5goJLl3
37m6Dm/G/0VtdBgyJsvIFv4dBOx5iUpBi7p0ReQJshicBwd0SfDflHYKyysYAvsf2n9b6S6BKNoU
IUAZBNRM4ptGLzxjEJaItpzBXIEyrpzxAPwZtHiQ9jLXb3aiWT3bUthBgevhKUZMN6mt9G0jEvg3
sENaWZ4GpwT/oQg8omOZFLsmrhr970KnX3zVqcUTmjiKauCPXOv421z6WvkvI1rwCVVqSPBHrWOy
/VHmNph8LdbVgGmSgEVzrQ7h2HFojvXlpuYkGeyMcpfn0ceQv7t6VwAstnX8NB73+r/xc6McWQLR
VJUgro3B4GBoJepo6SdUCf8CKMKvXxTQWNoeNxE29IQ/3w5bOcCNnHapkWBwEdqcC6y+jEkbmjql
iRm/fBO/c6DgYv9VTOAmXNNl+d85w336YkXAa0E6zB1KjceVnWxb9H3dkmSunCN40EFE6eFNVKob
349hnypwysKWLhxluNPVea0OI/JHPvxGACvOR2Tv9SCcsOkPikyYnNgeipQoCyx/t0/osxmLdHl/
ydlMTc6gc6cvKtAHCNFucV14zikb/UskpPr7/29niAxWH/TJStLT4lVg5eU7B8KRlsjFL4zeAQE9
4azEuYPYlZB3PlMtPP8HPZHZ8JdFjordaL8WrPMleW57/ZULpp/hJXLY6+gfzW9Qvz7TvJ93mr9F
bhOMuL1W2Rere4zPqezwPtYFbZTHCB7I2R/jopdw4pNBL5/pCNUh6lkoIQd3rTLw1SeGuWDVutz5
NcnQ3LcDHgsMUfMVuQG82dNMLB2DGYs5rRsETL9JS8waPdkSTSVKugJLE1ksLmJbBVq7qPZfJoub
GccF1G144g+wkzX+GgNiOdT85Eojq3WQL3HkKwKMKi7Bq7FfR7Uh7hcci1Ogl9vojYt0jGYhyywR
IeJe7VyFHPeT94yC9oOvpjxp96NDt1yRCw3oH+4UF/Is9rp3v3hGwk5JSRgN/2xFMzNewBuSe2ge
yWJcCFVv6H8G3uMU7pfmvWNqDJYTUbymh0PzwRISJf/nbM4dNliBx9T2ewpjULYFcJAQABL2FQqj
iCZ0Dj5g0+5fmb4YzRT4PTYq6C5DJGJ/bqYA+b4NTQ63djiQ/I1xUPr0DrPVnT6Ce7Vt0/X+uF7P
h7sEDt6KxPqTMIjRHYRfZWM4ohScw0HFNbE02f0/Myq32xRKDCnTUTLlj7164dHBt28SDDY6NE58
8IPqw4J5L1VIZFf7nOLQ8nqgtbMxDdLfbMGBTrQ8qiEK+NAi0QNScWrhx/w3gl+nX+Q1W6NXDU1o
QhmzE6kxS/9+EkhlpD/Z17eiuwW5+CpjcxMV23Ia+LKZpwuJZjQi3NdcsTsBHdxlgG/76pmej5HP
BHeAvHaRPXTlgOeE7eLemY1s6xslifk6qkuWi6VPv8vAXWDwr6lcGZNG01IsMd1kJjbp+8JKl8Ot
7Tr3PmGnU4MxPo3fYNXSDosyBoiGYVFTO3udFY8bcFHHAYF3qvMjJgJ/exyWcTgb73dxnlpr1brT
aIpc0O5tiVSEhOVAnN1eo/mbZSnD7die5bWt80/L1AWnRQT4rthG2Xkvo+WwjYI6cq5hpFErgpNR
Wf2NiC1W4MhCxYdo0uftPV3PNLBVyOmcBwUeN3c1h5TxNsnmvIIkoNd2+OE9LUSKvZ6TGhhnoCpo
s5gvSl6R3FWXnzeZQ5ZOm/e9V77jYzN0PAxFqiC4bf9QstYs07moQ2uFSId3WYKGsJJzQB68sXzC
TfPl6XB14ybCpYNYakR46oNENsi75REkLPWMDstN0PleiMY1NmELotxlIyE8j4G5xLgxNN+9UlvG
rtpi6UTtYswgiV9klCNEMptK8V7qFqyp7lWVwCWXuyMEujVYcct6A7rZFc4e9b6iYr46zbMSZhWn
56nntqgHtnnFNEAzxvLf5sK1gsaZ2hV/HtYQD9x1eUqjTvB2+qsEqoiK1p+WV0p19yqRtWRlEsxx
/aHudeuvcBs4hW+sOK0v5KmyyFi3wjFnLe0IaSWkJolan2brSkMcV3vvlDOuMzPHEN386+HGEXOp
BrZPzVIn5T+ibfrQRzEVtCW7E8695h6L+cmRNPc5/JwKh9L5eH96lrwuTHYS9KpwkE9qUIt+MhM6
hEoAG344+3esxsWRR+A+iLIoNwVBVPuY+S1RtVtcvo9NOyTF9T96y/q+hwvTNxltiy0WUmNmYnsF
Gge5tn3XZ3RX3DF/3m2O5PcpjSeYs+ZVBa61f7ZnyAZbuObUSjkftAF4N0yasIJ18Cgsgvn3ravf
uCkdEYFFFDyZe/XOWc5UGIHQ6/ScPss4OQvj6BF7LeFucshPbtmpY2nrqTTS7+MUEodsaW/MXSZU
9nCBOl65Mz+Si66eby3WsMrgR3dIphIIcgDNoV6OnIPVS/7Hu/KQaDCITV7syheuxfjHn64sish3
sFN52ZrEJSwW5cGA5FkrsEIYxezCaKyPrmgLZFhs7qcR9P1akpB/7W9eQAXAeWsWqzd3hCLpcu85
vks3vMKM3UF4gN2E8JL1ihwu7/cxQuNWqIOHs8Hj9b11ulZ5GVT0yatdA24ZlvZvCvrr7wQUJTLd
pxRdRZD06kYyth5NjIZkUWZtv5lnPCoXQ1nlOy6AgSKMkRzeXsj4LVM/jeJw+NhNrpDFUUKnS8v+
lEJRIwZvcBYR21bwuNmu1ITXSDpVimqSkecTUZAipbBBCqChQrrX78JNnyYfw1/y1/Fo5asHUUov
/rC7hYE0zOgDAg7fS7Zek85KoloU6LqZqaYdKlM6qQscQC3CKlD9kzPEzI8M80pqQSzxhXE4kswv
uSgWD2ZqXvcxuQDcHuntL3X63wZLG+PY7+1JGZc6vENzdXma2yTY+zetEtt8IFBpcLPhzvlWP2OL
dte91A2rEGoPnnaXmLH4MuhTposEsHFEYqKOrYMSAouL4qXtVAtTjJRDxEL9gPES9P8iLzlsjrN/
as1aO6vqQctN5uHcdX687GqcnKq4rpzxTX+Rkt9Q3a+4rfRXoySmx3KdV5BT/4oh2jwtZgfzIZHd
/O/pA7PSfKvxn4+UpuS0GOpEqC6AXYPFL5PBwKuLsjXYSUBpKj4uxeXZ+jCg3w0pO7mwffKtOE1y
gDde+p8TmPae8oHaTYZYLA4figwhtIT6CL8WU6Jbyg6JEDW/lxcYnVU6NHqApregVrMOmMF18z8x
jghtt3t91eVFIb7nCOqpBjaQg56EPwn6JZqcgKA/NqnqC2EhsA3W58F2XBNSYtsmkMSHk9L6RSso
880YJOW88wcdfV6uyWdCq5/Qc3DAPYR5Hlw3aKcWzgSY16/eE04o8Ugk9uEHHDUeupUJs+3sq9PP
hkTT8HOXuYnf/oVbSYthUMBXPqZlT5QATvjwG6Q/p5CSaO4eUHtOtCS6AbazkT++7NBuPQ2m8if1
updzlhFeXGO5RJWkBXAuAkUKzNFZoZNPNL2QX41kweVeSh+vcZViQq7C5db+jHNI9/xJ2rpw+OR0
PUR+MF/s95OyeISb/m1ALGPFS6qJw2c0vbDKb73/saoyzHUTdhLraHO/rWoFpsDCPWgd/r2C52ot
W5NJA8DFIlxKP0ZUMquD/8pJ0uIuDZo/AyCBz0eHZijHXygSSJG/z3NT6ruXntfCZ/86eEJ76guF
IocYsRSNPhP9HbORXhzfYbzwNPxcPV0AFnH7/iHP7OQ5bl+8krATqS5vUPdUmVZDK7HREZGBHBIv
W69FH9/fcYE5AEtC8iqybQUIM19G694HrniJ0+ZiGz+wg+wPFqpLQzOzPpRhGPtGA+NbVLwtJMAH
12wtZlg3IQYrBtekbwnHtQ3t8Rrz+DqOiEMOnWV8EbYVUzp/foMyUZM+HXVHi+lzd1hEoEGfM/rM
USTbs/dgUYdS86vRi7iCAFfXOdD7LkERukXHPTTkPHR2sShAz2EGLBEAoXm1HdMhueUZYbQsQH1b
SWaEMWKzhe8Teq12pyzpxW8Psj0kGe+REvDtNa2URWMgW4+F/nB5uaP/VcOEVE4H5UHKqTZZywcz
vSSR3CdpmZ0HjxsHfI3bcuV9lMXWs4NxkucyebEMRhdrtUJZmfD32OYsYqMEA37Rew4GyU5nA4Y/
+0E4x5IpPpzwNtqwGqLVsnDRg36O5Tmke9gWPajrh6Mkm3ZjhQuxqi2B2V9HYB92+IRArdWpYjTl
BHilhZE/H/tnjX/Znqtz6rWMYh7rz4wWv3b+TCgUQWPn4hZcXb5OJ/EAV9hCd0mYbm3q3S5xg2VV
XFru3G75Nd8QtofxfnOgTEisSCHd0XJpexGhxLavBkYmjzpFEUnUQbwpGwSrv5gxYLq9VzE4oteT
XnaDhBJlUVxbl4bQP2lhRN7JfRbUGQpPPX5vNdF2zJTCRxv5Lea0JTHr4GYRZoEtctCVGcv9EcOy
urCKRJF2NDqtBOoiRU3dh09VensT4hqp41i7sjkE/MgOqi9LL99J90DR9dSBXc50X5qggNLQv4eT
lnxuswxiFHwjt4bf5Ba2qmdVkDQP7bRUKABKTNgd6q4IRQIVXiZst2bmD/2INDZFyvAnrzwsJEpt
9f/qIG2vU1hTlONDdPSCn3+mg5+xLEeiX7UdIF4UPLGlTFNiAmekKC70ttdDjiWQRwvRACqYPuu7
b5E1GBMB3CtSJDvldTUmZBO1XEXz4GTVPjhjO5+ilxEmziOIXtDJowq1LU/dFMjHuU5xG8yttEmT
2+Cd7aOUhzz5DlleQGCdpnu0po7fA5S0MW4wXor9peT6iwsLG3PvgC4jJz+uZ1/fhtpdB4OBCTgu
bbKx/6aloOY5xDqn1LmkK8O1dqftz4MGVPGMBrCKmmp4abtGqHhovB8JLCbSw8P/1XTLl6U7pbbt
3mDXefjZOZpTjOCk9u4Sh2CV/alLITggoJG7gChpM26V99b02IoPvj/q1qXHi9OJFuWwI8MsxsGa
9vFh8I46MLiP5ycna+OerhQKb+2q/4OOqbuhHnq1Rphr2Xq9FE3l7/uUAQaXpfpZTPe2tYee4+iE
FsoXmQ5nk/gDXOBbgQzPyPVHFm8XbINqPqlBhvxbD0yZjRSiMoukgUE7ZcGUEbr5nKbrFu8xl0/z
/ij6rXYLXbDRHPDq02F/S1Ljpa4OApCUOVrOZgiPOgSPOQ5XaqXBp3YgQ53wzJfildq5qqWwTAXo
XWSbo+f9zsOvTQ1s5yhmJAhgM03nP/ko+V+H+Z1yJzNWLhdWI4x8lNJ9FpnAwUf8dcBWjZtOvYGK
Pg8/t7bGxM6y/SMe13nUWq4A+myXr8GduJsDGxbmak4286LBECKAFhH+A35q+6UDjCS3AQWyt8cL
NKfXmG+VHa6KfH0ou25gmO413Gjc3Dy4zsyBLJncgHKLL0A8vApClRAuNHIw5pu89rp/KnFLlZHN
27Nh/mGANhVx2pzpZknkqtxmulEI4NR/a9JTRzcYorTLK5Rw55TEA6tCIPTHsWx6XnPUM+d8yEET
5Zp9msIQfX3OGuPFIZGNhAU4AuSOcLWQ5w40m90Wd2K9F+tDy6iqhVNUoSU0taQ/J9zPpGPOjv+T
46EA/H8qY0/LMv3mRQqWzDcLjfy/MPunZnIVjDSVuq0XQHEeRF4NH25Errga3NEOLUrEW4BWOOMj
GhQEygl2MZcrQUv3Ve9I1knCdQQWkDaM6L4y39jH3gpIdZKwzo0bH9l0N4Xt7wPF3cBCQmgWtWh0
QQvs37Z64vjwnc9wRMXtX7jGP9nj+tlTAKmsuV97Mdb1HlH5VOKb+HkEhTLXn6oLeiHyEJxo9x/c
T9QyIzzxeB3v2J8rHw3lkb9cJ4v0AHsseix1eV5xJqYwoTrgKApP2HaTAx0+BWJqlvXCKQHVp7Wd
HQrgvc5U6qLsQSc5AQEQsJLpytG9CaL34qapTDOx3F+2OXrOxm+wLqsNbeyAEoAMy5lCRhJabQvX
/ZN8fkJ62SndfFs5oW7TpP6VfSpdhOzvNfAznKPwa0+eIrpZ7NS7OckHi7eBXmmW4ZnfkbGm/sle
YSKt5hr3SvSAyFJBADqj1kvAoGEdAVKD3aEP3B0e+4b7KLZIER6ioRyYSyAvdcwbp/PsDRqhxQpE
g/aJJ+ut/lKZ3n84dZPRsmFaaS8pG4bJuScefbE7mAfnOs0+yp+ZaWaSMHFPuw+ibLBICr+38UKw
DvaxjkCr3B6A72oVW+tf6nEA7h8ThTHwMkWcWvsx1M79JT/jfGOS0LFh0ZPJXWYNgN55V3yZRL8L
3y4hs0icVWw8TNYd8MuLYae7JmGfIbP/efDIwbsYKGg4oZiq5VoPm9YL1kNtS0pdY6QraPpblfAG
F6BVolD4xR78FLbKEi7ox+PLI/u15VVOsLjTdHOuYWgPlbaEmyBlYGs4gl2uc3H7s0M6PZdCIuE2
blP0GVP/umpxXNmvDmqnuBBZpvBZJxfGZ/kDrTtGthyGJ2sA3mOS7LNxqyvzmBtaqmqDY80HYVdy
1X2q7B712Hj5mpyQjN6bPLkHMRqvRxRnhEv65vn2sscm3tTM9LaIDweYCmpO3jyEhMqd58toMxMk
xgHqY0moGY/45es+8Y6ej6Y1CPd8U0YNtOnhRmrt/y/PmCguLiZKf8V/xt3AAgPuW0NFqBbi92OK
L+ztpdjveHYOaXJs09NdQ7jW7AypQP7pOGX6bz7mrFHDp3uJsTOoTkomIRgp5OTd8K9M6L8sup20
jiYLyRsIqpOv04gdZBBNWXomp71vCIEbO6nDqVFga6r8AKeSbpfIyj47shA9/bbQsIilFW4XCj0r
H40xw5ilFkMKcW8tAX/w9pZZUgu13/g71KiNeqCb02DkXYFgHi8oapm+bbm1fvZDezBd569JNE0p
MLLs7UMVbqthrT26v8vXowSxA8cRvfvHIM/xxXr82xTXsDvLzYOevK6Gi2NhsElnyRnEa+ZHTax+
K/ea2wZ7BQGQthhby3vHXvg7yptOJON+RRU+YDZykNat3F5NpQntZRDuvSMpbxR4daOXSRV1uehw
6xXECHtlyTAKr2k9+090QACJSjQgSZ45l8sRafp7+PxqxRX+BMDLkhKJ5R7E42/vzmErrkja+KfX
w38gQ072M5ugHF3380v4twSisboKH5NeBig5n6IMFQAhzfEhqk7pQUdZcitrCJwX9quEKHbKH8hE
KHBE6BiIxtzolKhFief8755gyF074dzpzi6tMSqj4qMNeob+SKjSFRsqSHXLDexE3FuGmabhEGFk
N1EUJRMy2tzdD4awq+WanxohgJ+w4A3KV0wrxCog73/4/0eBeoJo4s+ZHavkz6oNHD423NWXI/dQ
5BVkacWkCuYy0/95dnMnvSLNbIPaShCuNygXHcR8qsM7zira1ZlPMvPuUKcPUwEYQbZAUCF6N43a
dvFqqOjd2no2Bj6uSUqKrGYGZhOv4I3PZ8mDek2yy84yS603Zc2H9DG0sw8ZJXPbLv74uC/3/CYg
sZHqXK4bhB3TzPTyVBh8Qp7M6vvdaZN5/FYXDsjXF8xVz0B1D8J+fZ+tHLW82fjgOHWU85bl+sU7
xZEa+H/XjylihV1yVpkzJxRkgXOeYpz29XhAX+4Mj3O2AQomOOScRBWyFWrAwwRB1rSgGwfREh42
9kLGpD966kVAWNHPS9yyFFbdEKpqMHRTtq0SLTW6lYy9eJHmwAL6+BsX7DBSY+iKlO/O8/AV46Zl
f0AXWVB75mi4CU1uZEp4F9nexW2dny3RaWWBhDHUVLrqv6TYArnT926iMtTQMowGYiP/vvSCvG1u
DY05TAL1erNz+VIwPozeI45n/lR0FA2HxVMIF1oRFvWGsZFC/ZhvnyNwsRpEiP3CQeHD3C3J5+6d
/zy2q9UUmIZ+iMKuFnOaP0wBQ7GTwhD2z3pMxNlKBf/4Ot9dzQ+X7tVvw39GhXyVFngyqJuzRe5F
KCr7YVoXTK+6j8QBJRKrrR2JETK3iNEkcwdfo74i9q57MegMqgC+jtBxbeEsfobV8BLmwZD8hKK1
K2kghdEPjmX1tByTpIkyXxParRTrlYIaGmNufhJ9bwAAZT2+TI7igF+8O0tt6H52+klhENKFZrbD
F9e/87FBj7uCuMfkYQYduYmWpXoJ4/kwzDZJx4xl6J5z64LmrxON2+8M3r40CaFHFZSwB8Q9GCHj
5IEB7mw4d1NVZZERyO3SUhLwh/T3ix4+v8C7H8uoex09hDcgWGWAjvlR1Wh8zyUUu8ky7GtMf35B
j7HFsOL8qWJzAIxN1d6wm4sirE/7guQ/AyYgSqfeVzNHrr4+660UsIdyrh7Rv5KvUeQnAVs4OxTp
ClxdTuFIV2zwPVPA7YSgBlFvVPUCp/iHnqcQ8xoVPfRvp36tSV5AVRMLk11y5frRsTA9DzBgvPzK
6ed5j/SQjkqqw/Q9Zyx0C8l7JzAsDVUpQ0UQEqrqk1yPt+ZQskHCtS+DZxDf3mQ6BYUHS95VeCFL
lqBwqakG3VEDc5MRe+2u/uPa3fvlFNELMMZBmLG+G1Kk8KxG/s95n0mmiuWtmNp8Gzw31aWq1ho0
dCK5b87WvV16PPQV8IZYfnzLRTTDakmn/kkBRK0awEY3Dy3UlTfAlOPMacXOid5OXLaDyQAtvtnd
erIdDsrwXMawZn4UzTQ4wc0uUF91k4hb3Xs3KhS1bmnxMBKt+JmxMtc3QYFoIJ6gV6GQSSyQqk1p
JgC3wfxRC7tAhrtjHCQ7aRDXR+2+DXPyDf6d63u4l9bf6T2ehgoUCpbhgU96UZIlQfktlNXo7AUz
nn3UiF/DWCQ9yDcz+M+2agvXRoemQp3l/AXcs4W7+JMWxlUjdyu5cvAxZJPglAib4PX5U83H3iKU
I6fn8eLLEHrobuqprbShEqxIM3r+HKEPj0Rk61drCYsD2DyfW8QkLXMNu56LIn5iUhieJNUeCHrW
Np4VZDiIm5vGZgsQnwcVEeXtmn/dJym3Kywjp88h1KYjSd/9sGCWE5vtXRU7eEv0AUD/+iIYSqdn
EJO8YR3nCgiCp1yNIulsV5FzAMwnkHWsvJsqLu1VT7j75QYFoZCJGSP7WOdfiz7hAL6GV2LMTws+
HQZMMEH3vbBCs99h4cBy0KjE8ZmBzcgxRiE8czd0g8tHl3/E9fdgRGmWoCnSp9Icn6C3J4Q1Y52K
pHg7bsxBPwEJkVqCH4HZjjTuv9S6GlDhSAZyYB9d5qQ9idc6mKfbkPmifabH03tMud9eHtfB7/hO
dFHXAKZudGDTtY+lpNjggpbN+Tealr2NLXLGqiHWJnwm/NCOsskxnN+dohybLw+wmkJK0FN5Q8+b
8aBkl08FILyjtY5p4O7tDeZjBzO2Qj1o01CxoOmeCqeHwf2YJX96SnETvVEdhR6hPdMbFuaeyQf/
kM3+g4YsTnHqv8oDywN6UbS/S3zIta9yaonm8t8TOI8AqTeUXfnyxI0aFrb7KqM3Y1Zp/DAReQHG
FaUw7muj0nuSXxV7Wvejh7VS5UXH8Ttm6xRddUeHbcf/PNAKiGo4k7niW8n94NjItOgPevmJ8zeY
8EB452w+93VWxKKaP0vUTnp/hI/p3Xwbykwx9TUDzIRbwzj6SeifKbh6QP6o9opstuPDFsRGhSuX
3oM35SvfpJmyrxXoN47rnDBbVE6KB/TULXd9nrKjN07oPYCHYwVhvuhhmQACQK/bLihVCV1KYEEu
KdC4+tv8Fc0K9Y7hQq+lPlPMAD6E4jcjMC2BFp417dlhlkOE6whY5iEbgi21KVk7D5OmOIoXpURW
5kncxw/Yu6uTsTJoRJY2BXA+WBhlrZ2GkKaPKrUQWxnfE4pUB6wIY7IfLojfjn2RBuPtL0q9VaUM
SogAhjjZTzZqaFQIYcL8TUEoSj5xjVu96lHlfpMMLnpGGWZIzJdCLjPXMlfnLIv168jO9eXfOcOL
9RUUA2Xzjdc+NKmaloqiqMl4tsx7jfGu4Tge2sp6zliEdqh8twped1LDMrxAHcPHCA1xITmTCN0Y
OvOcfASY0k0y1pLdvaPDH5Fklgm/2+4E5awce6Ji9XBkrwwB1PMC1iRKo92vUElsfa0c1zYgsT9T
2wCYemSWaQmMsL6SMd9vl0/37ziIK/ZGjdoG7L/TLoMBqZiHlsMKcuGs96efgZaaiN2EIk6RQBtf
KDvQtjhQpfUiL1XMmnj2/T7LDOVAkK9FknxC5UASa+6JRzCmnxZafQRUkqUZ9oKJbiQ50ys+AdI9
1vWT6xwcmhkaDjJ1/KJsB9Xf5NRWDpScI5UStceQzKZgseIR/MHDQAGS5QCHJs7SOHYI6Kznguhz
EkU4GbXwfPbMjInDTTPN19zREhw+VT7CMnrVjtCny948GnUp6iNk9Cre7lzEeoULDPgTQW/BoFqi
8W+ICc8r3Nvy7EQvPrTHLX7hmSc7wMO7xe3qidMlWU7IiilOh5fbFfXS2KSY5jkBy3kFxho8Vsg8
tcRTaLVE65DILbl/jaJ9pAIWW1eMAEM/aGhBC7OrUePQ0zMAvICZ9LtADA9YmffO6xa8rwv4n4Lk
TRCztbFYCDAnFvEEkMi+NsQLDm3kLetVTeRFwXSBjkIlfvhsogQbll5plZUyqr6dsNsQuBgam2R1
H+kf15WialeFxTJ2C3hmSfnbmr3RAaE+FBjImITOKQUzOZEhG2eFSsCUnNDiZMROUeb8dQLgNRqH
K3PbYA8c06rJCJ6ZODXbrF9ck4jzwHKyOzWiYiZ6/q69aseuVsympjv/Bkk+xHO1/HyrmtgTEmRS
3QxwjPUSktc3Qj5NG+IZERUBnLTFe4RQ7AmFaswuxGQmxSdfInP/+Nbu3lqmuN1gFs7EK6pkBoOE
F11maMTZPPoWKPZ+ouz1U5h4yxquaCoRlIlCZZ3xEuv2RCCNuT6r0S84vgbGfZNZD3ce9ZWn10F+
F/tR6NK+HCHsQEfwynLicnXCKvcNUDEDZVB1Z8Uax7DwM3J9PJ+5XLw86wHeuFY8wmZxG+3uGf9I
YcLcGoVAUnZBM0hzMU3XMAsMDUA7s2Cy1BqCw0R+aPR/OzaUQkt5bWHqJann0QzAfQd5LHeXXzxe
f+aWh6uz604yoj5lLuFWdSAG+5hqcyG2B4Tv2N6CL0chQeL/Y8sxGRWXn5/zy85+Zugj2KkkkgGQ
AFY1/rVx1n7m10TNnypOCx17ZQZ/kt9kUHnLcMJiXeHReO6jPoeeozMgW4Crwih4qVsCSvCueLqh
6t9w7BUx7Od87cQlof0dRtQrbUW1FJp002wQsmEAOEricAFA2ymOvwcGBIYSekDj882eLSx6e0Ql
bXU6H+bOhqgMfmqy7UrLrucLRNdWQGZWm5ubThdRb4sJs9+pQWVR3H8zqTGvZ+Qcl7aTaQ5nfSxt
xwDosY1AtWl5xnpM7fc48KFRJkDUHtTSvLAhYnar8Jz3JztH6UFqbBQ3UNW89/JCJ5XH/1oMCSD6
GHPTut85U+RKBdNFqDuirJ/IFFjS0EM6/ILiH4Djya0X1QZx+0kOHGKzMWIa9/rBR57Gr9+FEzZI
/Ry/DQL7f+mSkq0uDrV7wljL/wUVSCNvj4Ble7Fh2xfUVbbO1a4a+TaHCZE53/6Ohw437Llfx2ra
xlHSCJJhUgf4EoYUMQR1YpRNYWdSSgMAX+rD3uXlOR1x4FIc+Nd6ZFrQZEl2XgXdqyQO2/Rfy+GQ
AyuE+uHMUFBJ3YM9ztgpP6Nep8CFHxU5Xx4YB5ftwUEKhssuuWC0dmnZ/wi18Hk2PFb0ufcvTELF
PXJm0UQID+Syazu6PiS/NDmEJ4DhPvHbfFL4mZwj08li2cpJ860CQ/JfI2cAY+yqOLjlyYSmTN0Y
BJfTM+MN14FxtHHYkCEwa9s0tz1pXFfmyGTe3e1GnVSGc5fDGWaE2kQa8mHEkZ97XPAuVvdsCE0z
9Wx3LS4pu/HKNypkpWFy7qQlC4yzGOEqReq2hzeMu/QQlbMu9ypg3zHHb39oLtQfJGLoB2cLUDeh
MvZDmHq4M4DBbGR7Y6eVEvlQzyVJAcxXSuN2uMBgZlv2jt/0/W8Q5kwgf1ZUloWJJ9+HuSaPki01
pWVnDW2j0KZYzxbm0y0crOtpDKLQ2xg/xbx3EOUFdel/dqJjzZ/af4n0eIvfUJZu6O77px+8nT8Y
4yvAMJqNSoEU0XNiyszSr4huOKoZd+6+shOhfQIDs9L6xQJoVJ6VgI5azOP7og+lCFuV7kIX6NTo
dYuSICoBNdz1xtNRpkJNt8Bdo3qT3RqOabJPy0oFEbhtmsruukuLqPd1bPRM6fB6FMd42TVOEhj0
R7XEK33QOmIW67J/YpiV4032mHj5BWUjA0SIWmxdULWhz85UVW/b1EaIQydQOzoAY085hs9L3Nm8
EXSMT5S3BwscQk/wZH5JHeUQZHsJStDyEnzgUCCcK0dcuGhevdoYdQfTNNlo0M0B1kunUVWjIsEI
IY3PCCT5Ii6erVqB81qo+AUy9ksHqSf8TsoTLzyni6vfM2oN1eoDx1JsXDgEltE30ZzwREHJS97N
O4oQS9X40Mv3ERzCM2UOjrGidFJQ0CB3bugHb0r6jJp3wjwp6BD3OKjgoW/jx6FgPbFIZxwok7Sz
CPWf9s+rCl/0h3liZICqNmN6DjR/FdtQaemqt+FwKSBShhD9U9zREXD7ZhGPyOGCcCwFAsbRM1gQ
7s7k5JZahEu2XmxCsm0M4lDvnkvuO7R1OLwagB28YvoFA5CSIpuehbnsAVeHzp8FK5B5tzYOXjRX
LEyBoD07yLRWc92oX5+S5V0ewiU/Cw7vBcXIDBO9g9WOO3Bwlxho7WtoCne05Ds6EJiKttY6HCHZ
zE3D597cCBgVG1JNjsmZCPgyyEha40zRQEVc9yR9PXsDxUNEZFopnDhXBxAASUq2lSxTnquiN57D
fxVdAiHWA6cdrSYcMmU0YjqOJb9f/i02FRB7WJyvH2KR/AJeMupqFbCGOMHGZLZl4yU4Rg4tHTo1
3ykVLCYSWyMGgy2HwPI0MlpJXw9cl5Ow1lXtTFiL6US2tXV2wB2idN1bYGNeHU9CE0a2DnrDC7Qn
ZrxQz+5zQgnQMMCqgvjgLDlKKGpQjo0ZGJBIOp3WZXDDJx53Ka5UJMB+FQHp6WCNb+JLwPwAlXYL
xXdEYoaBjBN2ygNEggr8sfy2SQNJVM/oYyjXNogWEw9BuAstMX04x3oWWHydBucZAvS9ZGDma5NO
IHqE1wy8NaoW6E4mrW59T2ubcWvf7ql5Kl4OGf3AyN6Jhvnt3LMsaLES88mg2ro+tFLMEjOyfhVa
j/Eqe2IGn4QgqAROvrXchlccyoTFIL53szXSTXOmH1gG3DwxF5/xNIIU5gAI29rp/Q554TJ9dJzx
8MyjEDuA7tVbutMFOqQkv/ftZw24Fyg34Gkv8gLWf4e7oouE4CQl/5UCAWpCcNKdMIy77B0aUSQ0
NF2kI+6Dr3R+SR488geigor4cvCo/1h5A91iu7yEvF9QAVf7vhddbIA+QGkMdyYDhhfx/MMp6ABg
NfRF0DKRm5RkothZl6UFw+6lX81nwYnc8m3yCZhnFFTqaPzQGcGq8HpSNM3Aju/O2TkhtOAt1UAX
aVXz5WjXDvxycn1Fev8KMLtikBkFGFvcLlN9cdjaGo3p6OgZKG3Y53eDneo2nosSnYlDe87IlMLu
1cRb/rwwiip3tDcMaSiuxTs3vEYUmQdeFXlsG5FpasxrPevsYy3SF2zRhTNjKrRmUPsiEk3cW8Fb
HrKELJPL/2R5e9dfYrJ7BvNKUyjbKLDVYEJ60PC/7DpkQWYM1f2yiiM+3V60mOiSMc/w94YBU2gc
uUwFwYZEsOQisV3TZ9Q1X8IfOvJMD5ESlOcAiZrqucOJcVzjupsZyy8pRlmdY+uIFbQ1s48l9yns
G935w/0NtF258tshm9XEwy3tpITtCUFQYJ216wgroe1pbgp36GizleL0YE+/xjMSHZcygAQNiSCe
ox9mq6FWrs/sYnW5/HOzx9x1UIIeWDCBP2/IfsQgJhpnu5usb/2Dv1emvYVD9oPVmAJclaJj+O41
l9TDb9yfXRZg02UzpEA3h6v7mlkjfHwy1L1Ifnz2PE6xAwpqj77h0UdbgdOlKeott1qUPzGeLG8V
bEh4xWWEBE6wTn/GkhfLNW5xWjuDlV62YVGKhQG7TxXn7RSkW9GfW/7ol1D7L3tUmocOEXXIHXKA
zUUXaTk522FMV1/CIgcbL2AhzUghggtp28Hj13wwYnVjYxe7Ty/l/UTii5GqSBCiaduGxE+suc/S
80qAfmwx5Ym4cHypQNdV/cMAvqjsOBi2awDq1jGjIBJBiIHSgosvM250nx9JBU6cVTK7TFFsvo+Z
rFZs0jZ/D4fDn4CylbLMrmpc0JZVWP0SHy2m4euOreON/UFR33aoFdoKIjl28rUei6UZwZEtxrZO
Z/o5r7SdsJpYnNpwabOLsMIepcu1su4mkg8+C1ro1OAxLgsvT2/UUPfbyHNGYKiZ+VpFaiF/7r1d
a5xOWt0PIJFHh0zoCsZvpYf4i9+HeZWVaG3K00XdPdG17edeM4NZPMp7y/g9lLNTblBAXILK+goB
KoiNFfZl9d9Z/iv1FWedKcGKnnpHcWTGhVdfb78RKGGFAFU2KAQ2Pvtfdvr9mzQDHEJFI+yyptXe
tl5Pcba37/NswVYd93YnyT8v65xyMSbmB21A/yNAWBZjBIaz6TCGTKMCad41fg8wcRdu9oQYMtoA
8+T7iRPyaTpXD7Nzkvtw3hPYEju0wXdh01wrbFN/NRPSD6jmwU5h9sifH+3Nb/JeaRDsqvNHpw1N
JhvFRzQah0SGpfsscrx4zVeCxL73eXFdYxTY9AuXWbmFwuaFUkUZQTMhx3iaQvyi0U+Bn+VHvfmI
B9t4bZEThN7Ob3NUw0bYp0spCWgU2zGi2uwO3zXmmz5/L3IlrSnLie4Cc1MDlIlTb4kFE3QpVRTC
7OZWupXhylYp0eEMV6F+VoWQgI6NJziINnriDACkxUnB+vHEE8ezYJ/y2dXOoMpE5MQKBnZ4d4mw
qw41XV6M+lkiK34dbxW+7UvsuIg0M1ssveCF7X9WMOKV1vjA9YhsNZVZKmaIFZHqJcF62CvXbkgs
8YQlEUmHbfk+6tAusgqPhg0qbka1dfBwBkIozw64+vW+PEDp7Q/oqx3agXxxZw//oReH0X56o7pO
wdplz6HBZh+fF1B0EkCU/KOtBGqjkqiIws+CR0oh8NbY1DfVpcRMC0/CnMxFy+OVkPzLrARGnxdq
xgQnHw2t7988d9XirSJh8WLE0KKXvSwYTWoqkJRrMDe1pxP2OgqffUBz3o5ou9zptOQJdwmOkRt1
4bZZUInM35kx1zqlaSQHBP9xsw7rKIRpKSrGlA9iZ69wF+nDuQ4yQNQkK//FNi0wHCFpBlfjLqCt
Pa4vTEcuUqA5QSkhISabOqXo72/sg1Y6hFTZFP/B23XhWG1QdDb8/nwVrtWCKZGazMao5oAxOXSo
t39W5eureQSjG99i3TWFO4CcMuNnBBTY0rQ5NBcfgacQb4oL0R79KUu98Pv8sY9EDMTihpdW064L
Umhq/8ESfv8Xzea66pQvWDOHiNDFbX54DcTgcGT/9phzh8dZNJM3qjAT76f1r8dMUcCtmU20+BNR
RbILnG43cbWznYWRZ5PNbgc0LBGM6J1rXJUzHj5/MJUsCgWvLd4MG6OdpJbusiwZZC5LCCa020e8
Fz0wllqz97p/RQF53nyyw2I3hjky8oHnBvqGsZggwM/VOBmV9nIJ4M4AETXMKvTSTKB13aJCNU3P
ydDorlTRj3e7po1EIopoarDGOFq01Bv0SKcEHe3EJxX0JFW6dUsVGOO48T01dmk9VvNZt3vNOTqM
aUQnoht12RbdoTJGJ2kPol/c3mgTWM0tLiQcqoA/mOEwMdFtD86GkXsfnbU2oXhKT0d0hzV8AZOq
ox3Vt9rva0C6EHmWlO7OU6vlOeYqirnRR3JlJnOG+Oo2jtrlWMtGd3u99iRxHTybzZeu8nN6YyiA
UvhYHQUpsB71kMl6RF4v8ajEmWcTwlJzKUBB2EJywb20yIrL4q3j0Z0lStrskFKiuM3HkQeIvd4q
/dZtfga9PV0IcTuD2iBf6H9ajHq9ZaWKDdlLZ5WscCuJXi46bUDww7Pjv/OHDvEN5Bsqj4lnpAQA
GV6iqKFG/w+LvhPXczkmLBJv4MBaEjCU93dJxQWsuw/x4+X6vGtloF46DmSm88EECPtyjCqk7InM
+wQGEG9slHs1rTcpMGq3msELeejz9XOi4kCDGxrYNfTIO45gl4AsnquSO3bDbt/8+zRl5+KSKFA7
ko2ZjxvNO691ege+v3ovIkkZNaupsZhpGT58h+QE7rGb8zxXAsMz6zBUksK9j5mgAzi6ALKpQPzH
7izLrNYjkXaFMseBtO9C8Il8HxKD2V0jfHdb4JoUj5BeyfvAgvRmi9xO8wnvQ8UqbMNYn91M7y5Z
LkZcUpvTorokk7TIHzBbfcjXapv+ywLe+Kwi3hnRHxpsJdDbWD3Kp5D0C+IlaS0Ih2J7Mw+2p6tu
SDaIlwQ3GBPw8RylyQZiX7F3TtYZXjPsagSZ49IYKZMM6LuM/IrJvNU30lCU+uaYJcZ6ReQS2L+j
h7+1OGGWnyMcvv30JbS3z5PJJv6yFLVk0h7nw0paHJoC9suhVWHpP2k7HsDUiq/Dqq2ybCsN70xB
iDyJ9Ckfc4b2aHd1duGqMlAcqNcZHAlKGql95bZnSg7LUTssYW+lGNhCfO26Ug4NVzPHIMpK4haZ
xQBHUBI0MGcg4mRnx3qfwYc9C3GB3kEcVbC/64ZYsFKJZNkenPsWCjdxajjf+SzkwLPIgVFQ4hSO
hG+BekwlyMS2ZtnAuQKYwDP1VOzceFDJ9zSmOJ/1us0i6yw1OrvONvpFG5abT0pFlFEWjcwTNftE
aNt+LsK5GcvUMBzdZxGW0h/h1npdTbULLuURYS68D7MvTELgNFfG/EUHjnbMI3DlJbuF8iKxj6K/
hKWLp6DLRo5YRTwYqmTRV4fKWd6dKgMgkEflSm5jKQxGggM+HclEIzCb76zwZTCgQoPb8EU8ifcc
9vjVjvTOscJ6b7tohT83Ii+3gG6DmSpWDYyS13GmYwBCYIqmZS2JWcJ9cuLW2+Gji8ugCCp/JAFz
dB31mBq+Ug++u+z0xfMpUd1EeWvAjwxtyLablUalbonOVDkvgrzfJm+2dpLtU/T0kMdanz7zW/rp
oldIqIY4zJn4tPzuK9RQATClZoU/v4hsObd7ygB1+Ez6JSZ91tJAd8zBszeV44ZygJ/YUacy2VXn
Lzyj1f6oM6emXrl2f8+iENr3+WSCVfLQhxK8DbA5sgSwRTsIO1iH+73ZJd1vEr8LqCt1n5OzFpjL
IIorsFPuKrJHYEn+wHgyb0RtJuaWlG2nJxfFAk8BU+dviOGmhmvg0raOCcQyW8A4qYnjQsxx4v/F
tSN/Y6e07N90oEtE1uK/Ltb4w9g5poB/eotAQw/IDmpDS3JI3+1dWFtWG6q+XN3o6f009LHwsdgG
gyu8yzjAieaPFbtMYeq60ew4UMARx+NwOv4erzymTiFJ3tO3BLZ7dNteCY96qES5NMXWvVpJKUoG
M43UlPgu7NeL4HQhJOMgQtbmSsE6GjqxA1m2CWvoDK53JtEWf2i4DZ28nH1oSOF/ZmpbHJKfzewE
bA7zxO20xUQ2lt+L1xec7ZlHeFOxm0XarRITBmNtb+iaeAS+vVydSIK8Q6VQhld6qXUm6LJ8lbH0
sK06o6kd6Ot9kvCZGtlaAUGgECN5BgB3RnkP6/gbToJwIwHjQ1xMJwM0oRhnQkH2blOnGlBxnlWe
2TZyL1TJna5+kDa1wl3Q20+E0Jtu6hiT4n8Xh1mOq/aIhk3QxgSp7sJiOxhGI3HWvEZ69SrF8Zph
s7v4ni/rMBszSYB9GbNxPqvKNt4YRWaRC7pWpPJnaoRH2g3D6ey+bm70MaRF7dQJffuCe9pmbvnD
uWeFvZHfh2cgMRjUOTa/uLPoVgisosSl985KVTt7fobWrzg4ZWqnME2TWx/LLaQMzso97jrkpU3B
WF1JrmycNY2jYkjjCpBntmsKwdTFmfnLt10cMk2R/H7DnoMIX34U2EDVvBALvc7F/VlB6aLGanGX
qvdxHyzPwv0uCvN/OetUR+eCNFqseztQKy/by2HRG0V9UBBVKBmHUDPlwnDPArpMppBkSPAXMxB7
pdOOic1sCjnKqavgHGwh6uBCsVOG5wVVYkVNhrROGiHLoytaun7WNNE6buRz6TJvo3qPU3Il+WYb
Zr0YjcbO4Q+HlUmo6JZ6puCqw9qTnI40a8jzNQvXRIgiD9itgt3wqsjNrJwQyWTKdnZF8C+mkfoU
colrM0TDrt1dJzJbrZ+cIAY2GNyKcgEmMk3qXuGqFYPLR6N3Ee/qsqbIgdZ/oHOK+kjx8YtMnOx2
7Mk5agtRmMJ4iqAE5pxqxy4/CSLja010yjGTnPdRIFe68vt7CvWn8WzesxFfwmKbJFGZcCGC0Qqb
/KNKg9IEWIN9F5mTk+MNU27mFxoNLrYY6MyKC6BOvJLCT3kJAjgGT/Hc9UCXKl3FItCdZw59ScEx
wdjTfg9+1ZrcAPI4FKqw/7v5bceQ3ASQwuBUA3gkN5oL7QWkGj8zqyrkSDxHm2iWtNE1K0fXt/h4
+uw48Y2xsEl1v7JDUyXd8BjhDHbwbSKNhLP+4YDHKWIC0s14pXgejs+jxSnNw+M003rs2cvcEvMZ
lSkcCXmLKcLiZubTS7u620X7QZrkNHFClIlEUYdjK2M8CMvEHDJdIkwKFmajCrr+Af5jnwwBfkE1
4K28DzNcLzOUMro8/bRS/CSy956IFqNxilLroqPr41Pt/WBNFIXFztt20qKPwP7b9a5Bnb/KK1cm
ZKIq+0swcGHRWTW274+Vbb1kNJjzl6DRkpAUxvHpiQKBZZVMRKAIaLptZGcqJ3E8n4Z2G4p6hjwh
/EXQi7kfD17ViHHotLj/NrnST5GMaBTfzvx5EyqLCehYwEI7qh5IXWcqFyc1r00zgpafnyJnAoKq
TDWUOaT4jCGRC536NW2FAFyJC0ihgdv13CH5rJFaDSDExxQZleELyXxjNTpc8473ovVC1RYyevBw
F2+854AcPZq+1roX+aeXqzRKxdwDAruKXwxhY1XIrwuTUYAX6gBz+t6KF+l+aFaKXcNFQisKGO6I
5ctM2UZ2CUAGM7ZgxLgcViKXNsdfzFYNqcpNHusdZGJTMz72/ulskAraxxjP8KTZpukksilCrV/i
9x3XUvkgKfb3M1w8sacHyx+7ABUNFlryNk7Gt3mLFMZ5zmbyZOsoVuSD4L21NneuoWN34ZqAStpv
vuilkvIlTsbOgeM6XuOMc4mIExQ9e6bZlKnzXbknZU5xv12NsvR4ZUKBLoeaxGIJtqW1ZHPCGKIh
PJK46IvJHZsHd8U2xNnJvktBGB4RRAbr5ZQjckq0jbFQgKd+IWgne/f3tAADewUmtGLVH9moIILb
/GvR9ASnUJrcJenk0GmHjCH+uRvNh8cXsrbk5IZG4MT8eDOwgE7FlJwoUXJwwmz3Hd0TkSDgIqaW
X+hZUQvtOmNhimkvch2i+IjxtHBPQlmxuLcrbZ81i7Rq8oHKjFKsLsxHrUNx+xesqgZ0MYM4SIVC
zqJDXhGpGlmTwHKiAd/P2WZK4aNry9ZtX5cz/QwJuftflegVvzwTCEqVfH+HrNmxS2Huz+nUAL7D
XeGt+OYY0n06nU/8Tp9JNU2IGuOJU8WaJQG7e8KM63LezLEdWr+bvcEOTyUB9kdmrLqsRDXm41Zu
nfq9cvQDPEv55lHPO5MgZBg0YbWboxPyycl3SUJPtSU6IASQcEKmbv8Ej5Z2tBFkFxhOUDOZuOu+
6ZoR0rigmC6O9krJZYVkW77SDsqM+GSGvAdEKhHXEcM07hFP03EFpd8TKxtj2Ij9Dt9T7jr2Cn18
BYLHcuTReYKYGtqxG6l5M/0tDigeHjSK2eoTTpPSwxsZq9hAd7L9Tw47v0cd3f5s3XLpag5A/CYP
kOfHy88nT6CnFbk/I128Fxt/8FjyfBNo/L2PkeMMvFnbOdLxfaBvndkQXV6ersDQOMPGjmCR3A2N
AebOG0EAtjg1T4J5TsQt6ZvTqTNXtMkmA90tYwY87X/aD3LAxiIZ88p8+zYgcIWmu2M480H9RbbT
Lp5puaDoOv6wrxPnmlsRiq8mHhNhIoDFWxTSlpIg3aIur5sUEPXGujFCMFzo/qpmzcdPembT0pGG
4aUHcy7SNbVHUbIsdivz+tgtxnGTwRHho9ZzctxBbdmhx6jx6uNH3k7p+sex/YcknVkSCQNbGtMa
U0Fi4+izCuFuskd3UMb5413knn0/XZ8T2OFgGMSDbGOIbLcS0nWCGloauRiNrH+kL0c3WW6NIm0H
BuwUw/oU6PLWasAgE4Var7UM3aP+TyI+r1Ai7Wmidl/nddWDvozjvuDHOsQgSgb0rXITalMR8JSp
9ig8ABLYnl6rs3UcZ7HMd17v1x1Y5KEKXGrsPZvuhxKzFgWsAhcPYwssKXCM3MOR26EHvIt7plDy
yOLiW4NU9MwIuM0HQgrQ2ouFWsm7YWaM/O8AruKuV2JJj2AC9uaEIn/MTpy9tmy/poWsSB4OckLx
nga3p8MwwwR1wF6UG0NuCmWJgk7Nux0Yn7HRAZA32uF2yOPJqA30DrMpzx9qEbxUJwCKvyHR3GdI
GN2yONB+quNBEjakPPPOuVqv4M3xXN7odWL//lilvp2ikVg/pz+0RDSrArm97xB/iU8t18Q4arMM
+N3PboPk0t0R6KbRUjHOCQBBrNeFfN+mVmvXxRQUiDal12qOJy9dvhjeL406nVK4QJ8l8S92JPRI
ZNreGxsK8J1Gl5l0K2saklhFht8ybf0ViYlFZbbeOGNG6RGZqt4LlmcZzTkb46jWtV5CyPCvpsfR
o/dQH+62KpouLm0fZJQVGDLCvWTZt0vobDuXVF6Vxd4fAjIA+3rhchuJEuSJlc67V4/uMWr8y9a7
cW+HByk6wcUOolw76U2hqWza109wzb6LhSwEctxtU7zU3sAlFhQ1dIJFx0Ba6wX027nZSCTJszbA
s59UeocgTkUy+wmHMIQ9vqC67GjyCj60Up0ehcnzkveKRhtkuMVHftYBMuRzIKxNwg4dnRpyvIT5
jO1Oeex74Knzn2bz09ttiIBdoMF0a6v7G93O5Ub1TfB1mhY6HW/V9jOznmKbv53PZpvpaP3xIS1u
CzePkbgmZUkvI+FyFDVFXtGtU3w2Rm75E7a7Ue2EvhqowZezjycyaJulBqORGpjZOPVsPPOUMXi/
dv0pM87wG2tnGBkmpIDcwTSqSgyNrRkMIrqnKE3gB6kdBDvZkLzCuAxnNOK4kyBEUTxuuFvaD5fd
qJ7MKEj4pzHEzwDfCvYkwuw6ghd2fYxTr2Yf2oDj0yYC5KlonCSBB/tbgALK2VQ0DAko2Ph1aqrj
0SeJEAr79k4dM7RdCJJ5SDjWiFcDwM3JqYna46Po3SH/u7gXEBD+oIkedzP7i2hkwBsQmmdJxvr6
SF5nDMzL9rpGRKtnwmJJkJh21A4TTACs5brInqGnXzQvCtZ9uAsfyp/wyZ/duwvrbpggkMcIbbUw
7fQncsKjletf/tncEJS+QoSzMqblfntHvC8YPZCT0Kq5sApheRSVsQ21EsVcEUUqmkYn6GlV+zdw
Rl+oh20M2w8/yTV0SAoPr8vhH+rA737CkBVM6twmJkRd4mWBatTj0pJaBQYhWwKQrHXJKoy/8MwB
bwPgPTruepTLDKVBHLnNmTHael+ETs95OFBz4dQbCPVI20EGnCq8kGAc0ntOQgvlKfErWjvVspfX
sHexmw/gyLGGp/0uHr3DEdBQKYsGUAysz9XfFku5RwgAQLqJXEn7LvnJWD+0qLrU+h7alit7gKLQ
jzo2RY5sBfWTJa0UXDb9mtZLb8zfg/TWNuw8Ca2C7UPJtt92KFxT0rK+10ut4tUlhYmxWi1/u2Vt
VNr1F1e39Tv7Lr/6pwDNUqUktHzU18I+DOJGl33gXFYqCzaM0Hun9SmU3WIkQoSs5FvTZ4eFEjRG
R4NyVcc7Ijf7abwnND3becJiBPgs2WkmuSbtsyVeqKNXftWb5qwJADHlwlt7ZXaBfDOXKob9Tmas
tMkxFkcL1+GH51qL2Sxl6uvBHu5Bmilq/CND9tm8GU+V4Fc/6HoVuX1ourD5pGf89U8OISzMk1Wx
lh5dEoRky73wxXvCUamvsQtfyswEI2Sjne/zNxcpxU5U4fdB5+B7ruDW+NQmC7ismIktuzfGmcb9
Ct34vkZTacqkkgg85xbEnZG5Dw3RT/Osyd/2+BbKQDrXv8rn3+U/CV2ZlQpEQkxH6kM+aEQ7obOb
0EjOE+qYXOCCkZzsiVMJgtOMUUwe3LQIqavKzgxttuZCF7Uy9vRWJjMXj2uSyxo8IEk6iQUF/CjX
OTGiCFyXVPedwFfWRvx+2cAnLHa6GsOYP+kbGJN8alqx8j6M5acmKUdx0SWfzuMID5kydLVIhE+/
UrbblvY5KWcy70uAKaTSIDzqyib0Gy4bZ8YUgCGJqGMIzNoMB358Sqi0sg6Rz4jfV370glmLl9Wa
cULbTIDb4NZ50hIlgFY5V4fZ3GE5bCqQ8+onbtQy5pdbEGrAEoyqC3FIuAMPwWxqCXohUVDUJSKT
WugOO9lh0zE8lyHVRdqrPlbCv96HS3Yy9EGesI0OCOwyMS/esOdpyO5TyiAf9M+W3UJHSOTDEPs9
0aUp1vhrq7rl1fzUUDgopI4BP0ayNAOTYdOXhnKh25J2DA5e88C6QNX2O3dMwT3i1yqFhE5oNtYr
VC12r7GjbZ7HZWn7WKh8PP7OP67VfJmz/uU+XecTCwa9HByiuz0El576WuMsMYwCQ9gml1Ad9B9w
bJaXj2Rdvyr1EsXgyt/qgYC9E1tznjRyjXznadebJZv/m0NXQl1HLHx9wciREvaoR7PhkYu/iDol
Bf2aQ62cKXGXreVxQY4MI1CAGTug4XkzH26SQZyREsV3WE2CRz8DZmAbq8TljrqRyjeVMxUlzyp8
PK3ib2Qo2Rs5BsqQC2DbQSUugSUvar0w+QWyJldrnKE//GyhZzOiw4MK4IKi9MLbp6oExumEZhup
r4hO+AE61DJmd0EuM6hQ4RzF1OJnj7raZn+T0mZv4iMmQ21F13PB0pYxLDnvU+aNKSXn6OHPMxIp
FiO51YNlZS1uEM32xAAf7PxDiMlnT0HJTKzrY02YnCbp8bZfVdDVBtrTLIbhN0pugbsQRZ1JfQSs
Ey+SFXlxCeOStEqh1Ch6V6tn7jmanqofnjroXFKiL70iPD0Q1uviyccVHqsxhWrxZ3aOYXHwrRZn
9NK3LMR13qRB336jEUGrTYhhxKERqytSIBeoqwIHlSvHo971++LJhKeuZZVYopdn27ffxbOe9Nq+
jX5F+W34cjO2osTEkSMfDLcQJkw5N4OIS6X+aPxJcdhSEmYkPewPqNL1dYx1el8skm95GoeBpAAF
3atNx7gAPL1FJyqie4BfC6M7e+F2azR/a8btIBp8c8aFVuRE/iAxstbP7DOSOFDdW66WIX4jRBz+
nrahdcQPTkTx5JArvDSlif1SbMKQTB7KCKFpkwVC2zfpfSl/ev+rdL2Sq6pkCNz37Idqq0R8TGyj
VHBM2ro2B9ORVn5UlwL9V81wp5xZrf8xu0/sWkEsLynZ+HszwMXrIQ73+HeV5VQSXd7m2j6rP2D1
yTCfkzdCkWR5I9rJNCwb6ZXzzvVoA+NMUJaj0/OqVcBpEm+Oqryxf8VS9dAr/BNFl7SxN2cTc5Sh
JL+vm/DSYK5AhAWk/PNsYPWACf7zgnnL8LlEskbGLqoyAIVeGpeb1loaHjYhOUyTrFyTVv224UY5
zQiW025A0Zd9fUwyJSg0vzaIe/Bq7wcvvDyyTVQOBMM8kcVuxCb5sendveKz2hUGHUyfedBQ2Xhn
ce3vE96pGUN79Te80f78hYNXGcFJimu9H5eqd93OwWpRmBDtqXhEebTU8MMYMidGMbJp7X9nc6qT
WN/0KQgypoOTF5wUqfh7U5TTjFoGuiIJeIsJ6KuRfzVUv2mEqbS/XMyOk3OurgDX41EBbHLhbu/S
Cw4Q67Tms3CpEfmva7Wm07Iw2cLRvB+Kv39Ofr7WGlif4/h8iilnUD09deixIrmuf+3acivqVDEG
4DDqDuFBqz0CDuNBIiQgmBH0zLFZVKsG0xi0d5HLaa5jemi7GIS59A32FH+o2Ylud4/OZYSm0sIT
OGE1QqvPaaHPNrtgY/HAspskiZohhSl04QoL5qZn1hVCyiOnKrLjEGcjD+OPgu+5mdGH/cj38hqn
WA5LKKO9WNp6FywVfxEV1cGQ1ICt0sifvnHLuoP9SSvzL6ivZr3KRo8M0OT/XI6adQHP+WtLCMB6
ClNU3okRmCq7VcQigiBrloczlC+3ky0Pg7vvd1ss+e0S9LESgWG2wP/9LHhDxoxzmb8fJet+QP2N
oP+3jxxzgnLGODI1I/Bs4l34D7W9yW1gkM7E/2Xq3Er2pRSby/NvxWD0nGFB207uuhuzJG55tdbQ
lakwZFNZ9sKiARHc3Nfdpt3aWgwzR146r7WDxjIKe0rp4BOm7d9w9JAe8kooG6xZjg4llZ+ol//4
vUPPxPY1tbgvbluixk/lFY0h3e81HYdv29e92YE8kQ/GkG+vOhnKnzyIhI1q1vFdNS5mGgPX7Nms
CVNpB6l9EbLnBsUIdpIaoxJ4mHGTstksQdOiKN41XBTbigyTlvPIDNaVd7a7fAX+iZsKbsGTljSy
bvwBad54wmBBlIYMeMI1lilDVndAYWnx3aYm19ayNbXBmW28I+cUJHZLWDybIzfNdBOUMXTb65To
x3MSqdvhTaZyAPwxPYSG++lnDzEmDlqoX27Qyon8U3X2W9RJ4J2bt/6kScHH9NgO6vE1y3fLnaID
pN7F7JCE5u5Hgm0uRjsvF5UcRizyxuVv3FyghbZLqp0OacRIRLPcO+1glu0UJavXQFtoqtUMmW9N
sgvVZVy8/kvQAoK5oKnM2bYUGne0C+hJmxiC8a92Ugokpv/sUZSWHTuEtK7ap0rnM+O7z3Tuu2re
bxTeeDLBXBWHkfCFmXt6n8DY8KTlpgmmWRjFNPZguh/eEWa6S5XHN4MawIu4+khbqgO6RODQIC5B
xb2o83ICCQk28JfBdkKY1WxzNno/XiaJa1W3XcUKbsIAjcAcNVBOq9kyS7NyqIPv3cyfgLdoJGCP
pbyxM43b9t3sRthk1sKd5c4HVA8H2YbCehtA15IEWaZIoe/i0cjx4JunwAUuOKr88vohYAOUyUtP
fOSViZPS6g3l8uSIdSSyIg6SJHP6C+y8gw7Cg26HiKr4Eo0a1B+Qi8rLcHnwtbq5zF9bXrJN6PTo
0W9/+DymJ50KV3por3tygJbi6oV62WAhEDBRB20ucty0TlT0VKMK83LYGo+4ULs62eFb16WT1Ir/
PpFbE9uWKkcVEOOFlpiIvQzAbvvOfpjpL7H/HQ3HP8FCdl29L1x8H7MoxWrUnl2fYEwIDMrrSMcB
ejJ1dFbQcfCeGYTeENizEyNvdg0T6coix71Ynl1IJeZBAHzSDGCxUtzcApQ4DT4LkebuBO7uDjfD
p8SXOqYDTbxgqE9sJXGa6tdR7T/vBqw6hrEqaIiKknkq0wSG0+xNuSM/jmIoR4hnoTO3rbmSg7s/
mnNHrK9M7kAkQrDmH/wVRyj3LlKIh6QmZeO1Lfe61ojeUSzcy9Y8a5etUH86hKte29kb2hKbCyKZ
aOyzkzPMp3oqhwibbbwDjipuDNIl/FmYpju+Ontj05+HJBufqIakLZCPPblqpVxGOyYppI69p7W4
4sYLJKe3ncRNe5kqgjAMXQ0SbwJUzO9817HDdBnq09D2Rs2Nl3ZeK2g/bpKJTiZ5xvg+9yqPtwlu
qkWEVxlGaSogqa0lNSullGTF5tPxYSmlfIbmjR4KFXsjcrm0A61I7318Vtv1M6tdhB68HcKtEmU8
I/Yo3fCd2PyYJkpB0lTt+ffB/v8sD0jxyaGjH0aRge6YV+kZdQm1FjUCZpMUjPukZnp7OS7LZZFm
k+4LWhdFlUjw0BqFuTrz53MwDeM4qrFfOzyUuMaFc6K6UzfeNs67o+/tptVYc+FHy9ch9+e9Vy/1
WPe2BXp4drZ16/duYBeB0VabRSm1NzXaSYT4qREXreylfG+iTQ1NgzXb49wDyOdlw4xW0rkKrebx
b9O3fLTmFSmyVH0DKgensijbYuFzWsQ88rd2dSJbPc01rTzsim7Oiy/bFE8rxDwNkgffDIzjjjYS
36DXuf5Mc0zy4sNDonh8XWPAIoDwKf1oW96turQT/rcMGFa0kuGFVqD+4Nry5R159RrCdPMfQ0hN
5xmrpHhXc2Yy/jinyqvvqSrgT96xs6EZ3nlwRHddbOEtpLYATKxaSZ3miM0OaBujWLSjC5/JiYjj
HMdZ0em2aANfs6G5DDt5zHQ4vzmq5piLKjCwyXaDT5bK6QzicSNsU9vyNGuPPBMX9ZkUYDwDec/1
jTRHlzZRxdRAIt2PS1tpfw7friFXKTEcUhv41NJAcsOnokxFV8MGXLoQa7JTSUTJNOaxvhXnfM0r
ulpSjNVJsoHEwOJL4NOZ7bCpH8LVXaEgrosRxLUY9U9zK0ZmTgjJowNj3cqON4AYz6xZ0Hvxx5n/
e60vrxTO00M4Y5z2h2AnC+Gq5G6zeRMWNbXvwDLAT6jhF+yy3QRHpT8pivrOm1efNN7qKXPKYVyV
rG1qjrCyKW7ztybbPzSuH3hGRNojwXFaDaSy3oQOrQqCo7NDNAtsijDctAcCHdizShgQRxKgIbNN
zhj+UDAyHrEqqTyUzP32OIRbIPOivTFnZe/mg/5x3ZgcNP+OWGKDWUTtOVewPq3Q8HtXpZ4/mfHr
65wOmT+wbLjLvy45hm1qwISYsjezQ+use0BpO4YRzQEmm3VCySH0iiNPPULLeRm82S9V8JtE//hs
bhoXPUq3NuAV3U0AxNvUQ7oAhvFtA5kp7UMqZyV9f0nyKJFvXnlLAePyKWhOMGAGVGkCZ6s3Qwtn
xugeyEIAun6vyQO1g9vOobPZmZPqryYr4TvqKgZSu+obswLd9uRFfXxWMlX+/35XfvD1mIn3G1yC
qqGIYC/Qnb1IIDo7EqZJpR/+uINIdwFuT7HpaMkin/B2f7wU8U7k3c9kgMwB8lvp3SM0i6HlUE76
dzifsUAEO2YDLJplT36eMhaG3STE32stRaQBQZU+cWah/9c33DfOMJhEUMClHZ6WhJAnBYbOsR7b
fdu6DE/pH/mu8ZqajToRzpRuotJZn06Pm/sMCHViZqTOCq5NtN2jGyIfcHuogaWes8IXhNnlxh/O
Oybet5HYP1ujtp4Jctyr+/K9LsmJZIa+4TmlqSjgADou9cmL8RguWSPA7+OoF9/7ROw5zg6Brrtn
D4OBcBggrDlIii8PG05RGeWj6HiUBTi7fgDUdnLmdRM0beswsSBiCrGvMQhsDHlZCxQbf4CaZXo4
0tUOAqF4ZeFKz88mCo+gbQyEdMbsfkCtHe4UN6it58cGw01J2+8v/C3TRG/qFmJGvE+uJEQV2nGv
/MDEJ1SiC+bJyoggrhaSJVMxWdmpIX9wACNGlxaFURSCqBaEedGMI1SqDpPlul4hJyqt4WrJDNeb
tLiYegmejkOO4aU+kUt+YAtiZGbUJverwzfitKeS+yn76MGqbeZTqfUvHxFpniGfPnFGY5YCGKWI
/Ickzs2lXK/EsSsrgU99rV22xBcdOM9ZAhca/72ZPB1E/FK2nhTYnhENUuyuOzmgB723bGMNGIDy
AXtmpF52+PesjA7pOD9+Jk6jVb61tiJ3+Wh1ZKjaqJtupdh942q5HTDsYX0Y0DA6cjcRvjGswnfQ
ioe9yMWK/tCZ1k0q0wCVZDSyUD5D+tdMzZs3b8ovxzo64H3FZ74WUol5Z+kn0rxWIAyG2ot3rw0e
w06jysl/AyU0kxNw1ENvraGlyU1q2gIbreMLHhz0LUgdW6k+bGEYYM04QcXxcQeK7LNBML8YWwHq
KWCUY3F0glcOjHp3qFix5G4P0WH5OC5vRRjDem01Ev2wEFeIaG0FwEFfVBNGWdR2Yb25quPY6mb/
pWTdbUONF7DlPt+wVlrqNi62ggH5dZIJmoUhfiKhciJfxQGfND9RfVXm2Xk1rnxq9BmEkjZwq2Xr
m/TCmgtk+DPKbI1rt9nBlTqbj6ijZqY6drhaJ5uDXGGnATpzLyTQ5k7UVxFIGa6Jm7mHtLHo4ga7
w+zttbcIzI9unLsjpYoS8hSVaHCD8l7qpGZFi3+gNEjQqvALZXMe5KAXcANYBg6pI/NYgoelOpxH
rUta9CbG+8udGdtOrGgNwUiTCdeU2LQUGfZlsniznMD6gtsEUqcWlIE8RKnhJLmwnTLcSH6nGDBP
bVdY+H7pBvoTVkOcU5pd2BiRZr869dArnGzeRKAkmiEY/W3hF6uFtXJE9rYC/5f3AIzpiAKI/C7d
Yu1JmEqFuW1F6wn8bvQJDgg82LbLmPr73of7MoPz69QEExijVb5/ursmz5FabH625TxeaWA7oAKG
AIzWZ/SbJtM847oImTIOZ38skrIFJGt836vpmjo/njcmy1/M72X4zoh/PesDU2LfjRBtLK9S/zVo
JS7B3rQp5Enmwqkh4bSiazcjgxyt5AIv2Kr9A02ZHwoI7u99rh0njnDbByrlDo2vCzwWUF3RdWle
kXprvG21nTxWzO+cL0uoQYiqPPB/7IASR+z6mrjsD3abMSJ96dlsQ8/rBkd7OLxAdVLjo4fKuOv9
R9/xdFDnxqyffn52EWKRjRQ3ikHlX1k+nJ864pDvTcSiX6bdoBKMHyt4/TCtSC4oYQGz5zf9OlXm
0a/lX6vQXU+7NQ7Jdk+Khqyx9jjpL+gus0ne4NMRCmWKUN3hkR35s8NDFkVaqdJAfucrMB91LjoO
y53oE0SnG3gcFbSH1t6W14oQZjb91daE5HoScU99KwvV1BWErr4NdSx3ZuAeMM6D86gHiyi5f3+b
n4ZC71oMSEFKWP/YVSpqegiYho/xWG7U5DEBHZGkfaKWJc8wd6hnc8UzuzKSo8gPDr2r2zdYMYSi
cavdaqvEWZSPdgqq6e25+ZKnMF8ew2U95l8WM0Owc5jqd/TE8wt6FzWiGJDHh2fbRyyzGE50dU1q
SJcHFKQmqABKFuCHk1W3bZS5Lhjx2KBPWgSrrPhZiP/Tnx3pVPIaqbJGlbFB56tDjcn0BUtQt1Ql
pTdvZp1H3Brq9ovONCdUNEgE4YU8GqmCzG71yL6BKMvDn85Ejv3k9h4aDsNCPS922TjwRQZq5Zxx
3DedIxJmBOFWMyhOe9k3L6Sku9cs2B/3q+Wqnin+wRuBE9alzcDVdDzpyuOcDqL4y2rcUG8dMSbG
SSHIuoiOfd7ZaGHixrotqtFPXyFlxSQlTa9YC/SePJjVLP76gUVYuwgYCMi/o1f81+mFhStLuReb
Dnta484nxwa3Deazrl9NIysmeu/8YDgxqpw9QC9E9GnWIVz0f2DoHAguV1Y3P2eqDFoI1AbBUDEB
AhkB9dXFyTXFXmG7U5veAA4iuG4Z28hSdON1irIjfOTOZxKqkfrW6KrmXBYIqHmTKevlv3M8fo8w
2YyHHT02U3jKjmR/NAqJQZ9XiFeUKGK/vMzRDLn5AuNEWt1+8rf8h1ZNdQqzzbHR3X3OkYBAI243
GfkbdMC8E3o+yeEjU4ZAZ7dqzV80ZyHugh8GRGyIV+HWZQZX8/NcKmlBhuGoPzv+v+IJ6bv7Z+x4
T65LQk0sPw+Z4W9ADOAucEK/8Y3svqPkNkS1fl2PrQOUEvZByBtp/0XdiA50GMTO4sWyjJ4TxHNq
YqClOiwGQtUj6GxmSqAh1R4inz9rYMA03Y07LLraTPOja0tAFudMcFulukRUVqO3tfETiZbvfMZu
65KkOe/zW7agPa8lV0x+gR5WY1eEU0N+v1C95U6R5bFdpevLYjWg/PJyPaTxXBSM2SKkfs25MFFx
QvQrlHr4XfDUt6l2dGsDcZGBB1vvdnVZ/Y4qsrdfba63J1zil0GJWaMXao0IpMHX8XPPN8t4CSuG
H3Z9l6k1h/U/iHgb7NhAQM96gq8X7gqFwOloCkMQWwC6YuNrq9HoPuLHoYZ81fK475ihv2y6XXVY
tJzSwg1y+P2azQQ3qW076oL0R3J5mpnWsqRVbsCdbj3Xt1eHdcJBTf3X8SaVhlxesOOS9himpOql
dzxoQKSP+5UUoHHS8u/7KrhVkEMMGpLjiLuDN4tvl1JjbWvhu6dbIfvHQ71FJDJOAb890ZOzc95w
0xI0ZxKzoKMPbYLn382W/73J5Onc5e1LfzQX/OZCq4gUW2sRCKnPefBGA/5oMw/eVpvje0LHgkkE
lu30eOa49C2kFOoYfeKLzr70UesJxQbTJ01BxM2y4AH5JPwYpQOKijX/9L6/oG5HbdJsRgyFPJfO
7KXei+jQhzHUABli+w1hCOF7pauWPODa9QAO7H2Zofl6yjX+t4pmqArL8cAMngImEJyjSOueBpyd
xklMIUz4lPJSV7HZmsbTQSTXWJOspCI/fcvyMMGC4bUZo05C6BwTWsZIb9BHThOvkn5/iTxng3Ms
1olUmtfs+bGmm/Le+SkHBNsvUB64UHNLHQdp5ijubuaLmoRnIL4d1tgYvBDS1LMQE18nqLfKn67R
xD9dRQc6vZIkMFns1RevxgVnNncGw3RZI9LFY5KC9QYslHC9sfz571n5YAz8GB+iVF0UGxEGJlUW
wMTaserI+2hWTVHapaK8ecwN3sbyJKoCbSkY1VDV850BpA9CIDanwWTjZB9V2qSSGAV6mg12P/of
5M0Q9WRdJVh55croei3hs7x5b6aUWwmDcwJyUxNNYiz+2hIEVJgcg/DPlg27IMXG+W5wVESAk8oy
4KO9EqMbP6S5tC8vHtTKH1HAHnuw/KNACrtI0gdycK0ofYw564Mtcj94EK+NpASsUl37dsBH2cCM
kZItbHPAXSjyfOk1+tm3CT+essCUhRz1J4u3GV/7woFqSw9+Su+/2UbNq4Gjpxg5lqRi+c3w9sUr
rfrS7faY9lpZzh1/7o3KmUftWlf4YF/ElMeiR7ubsM5ddlWuIA8WFvFkOXqamc17ORqgrGDpzPAj
JXiDBv4Wx0wNILPAgAApugKwhR1pwIPNEyGnck5tYD2EdqAn9y7f0DfHEHlw4PPTVEhtdzTr3jD3
eMa/Lmvq/k67oELt61uL7fVe2TbC5vdNWNof3u17NJIA2vZmMypP9+fenFt+so8vuppdT76kaCA0
z+DANHcNQ/L4XtdnqY7Uu1RTPQdqndYz8LaTgsp6CWlvzirgh0AUtaOjRM3q8jn9vfMFSUS2zwVG
c+Sp6fZWRKn/xoF/1i+sQq5TOvZVLl+RbulqpMuDXjJj9I7as9hoUY1OFExbgj/SdvarkAKaj41H
kSqn4fhtKYHsi3TM+yPzxU1F9NiW1QjVG3TBTT+m6/Y1KaMSf+cpn6L2WCl3JLg7mt26cZzDtINW
gQpNi/2PA1jVQS0RSTR+ZBTkvIMMiP8mjTPfzcTAJrru2EmHi86cSlpVqSUd4N+5mHwOR1nx/lv6
gp67wxjpHhe4nrfV8O0+kK17iCtjkKnf4VmPoRJgJzONR9OWEATrLkZPLDIsGWkqgGioQqYqyyD7
xJ0wXVzXqhkXLgvJBwtAQx5y29WdaXM11GZJPYF3bwjaSml6MnZ1AmLsxNa84r3eadPot0/t0iHm
dEjVjh04HZPO6R5lHsEOql0YXD3dnBJnxEz8xbbT9MhM/+5rAi6X32ptwglDDuQW/VqF1RFUlez2
RrxmX/oRBvaGSh8zS9krghMmw2NGZ9lYaS8qCCQFlv0sdOW0NzZ9B8x0fNFBA3FgqMUKX8qr8NWb
2y7dg6PqKfbfaJ5r8Rn8ot21LPLUGLmbwgolZ1juSdPHjZoD9luC7EqHuoyp7lC5EZY18//Vg0YI
BR6gs8IhZpRTVMHtso4SDtK53V7stO5vunUiMe+vxbM7LNIu9i/ipxmBJW/Rr49+YZNBlvspsDKs
Sb9cBYa0cvk2pWvYwekQvbUDxYghmLqyhaYKR7AVN2VyIIdB58ZvRJpHiej/eQWzgVg8H6K62R8Y
QNNDUEStbr+VEjxtWrA70+gv2CM733WO83hPeL9W8z87DoFuh7v0lStW4Naz+C14wBGrvATPnypg
OcTbYc+f+xNmzyRXSbcy8WVmi3w8JtEVHfQWxmGrhHXdrNd0QRBCVCLFDgHAaqG9Mn5WUK0/creY
aRjovglq+DWB+BIz2Mw2KPrVUOCo/CAyL0zqw3Aj7w2V9il95O0/EWO7aVemWx5ACCu2t703CMLE
Jr5mTq/j67DHsRqBBY1EGNJ3p6o4pPsccIypbz1tJUi4nNexyX1f6DZAOcMh8BjiadnfGE5MIKjB
vooU95NUe5lIIITxXDGAMAZoysjbpfWCfMUwhjqZCsJu/BG0HCyNWISM6+GFBg3mxnDIjcSkW8bJ
wsf5adKeEXmxxskNJYk4VF6bg9RKdjRMATZNxyMziN0kSQn4eloBmu3KzUVNpdP3UgSC5a6yihEq
NwGhIM2lu5GXXo/z5A2hLoMXNG7fTOQUv9YPWVNbA8YptzkZHVpPMbyLMRcmtKjZUWMUkECL5OQb
D5UEtcSn3K7XkYfjxi8NjeziStAjUiY7IL8x00dtKdXXvQfQ9lm1N8q00NALMeRwcYeoiBTER/4v
VbdpITlU5Nmq3eameTsZVabxrcRHTF4YdygBHMoP9WN/RmuFryZxjr7KluMDn/oOETfMe0w8Hyiy
M2I8jHziPU2753Rf9WIpUap50ZH3k2QNDBoqV/U0K8ln8MjpV4Wcz7btPBZF0K4nMB4lDJagrIy6
0f4CuyNttd6167kKC4ZtvPh7OAsDqbwoUh/iaEQ4HmVEIdl9mLu4sg2qPyi7aOS6eTg7tdh/BpGE
jjr3ImyomZ+X6tmFt+d6E0YvB0LpqO8CLw5IdWFSePsNiKluULED1FIFqLnG/WtdRd/9mvKXNYbS
KLZk9Aq163GnM44Uyp8hDUIQz4ztpH9ybD2SM1XGj7VMUwp6ylLPwd982cIRbmSSK7L1rcycsceN
bhr4T7KeUsk2t9Am6uVlFI2hjOtHsP7cV46iJoug6yO+qsql5xbHjGhYn/iyFurX4Ac4l9eHUS0m
QnwH0T7K1aBclbqyG7fljTgwGDdhX1EoBUjY7dyASum9c/06kNl2I++7WNZbJ5e0Ktt/h9b13hBL
4nHMk+PnkjQm56JP1DAGutSj40Pb5f6QCSlS4u0liAlavyaMz/bqoF/v163i1GURgfCNkjHh4EMK
IrPt01LYOJitbe8YbH7CV9/UvVxbc455p8YnIoE/fJzrs9g87EabV+VLMwYaAuQWk5am6zBPNByX
28PxsswN/6uiEm/8wZbWWlaKHSa10bhpCk534Er8DQR9Kge2K0f4efYJ7GoHGl6mTe2AyiN7yLzz
9s5djWq0SO45/32PrlP/ZxH0NUYTTL4so37Xqvil7Zaq+Hc9wSpK6BzEXQOmFRtbHS7Hh3JKys5u
kcgyUIULoyGBAYbWSWuAIjbc8oKgck1kq9FGDU5ys2oVLoVc+bs+8j36tZnZQebLVclkymTmojLC
lDEQji95Fa2E74QSSYaxrZXyEn1BdqJWNtmznhjhsKRFzFxPIWuRLxKWc3b9AKRUMybc5ZAsrEpz
zWlgCDJzYx7IzlEbmyLRrTI9q76uxLbyO45IZJ5DRsniR46I2+GxcBrnQYLtQnVHFPiojeb/nJSL
KyTcqzpNBDKp6alwNUzKeBmqumZd3CUsdIrYo4qfz+F99H03Y4FWrylR5V1bkfXjpBUlJV68FpqQ
s0sCM/psn51I99pVNhrSctA7PibIsql7rgjoCvjd4qJR/OtNf5h0HGa/F2KAvgIw0iqQ5FtUzgQx
lym/yWOamFLL1VGbCx27IntGUNfP7uYnt6RaxRgHxEK/Abyfilz9OHqXU1rzwRmoqpFNHc+vXzVq
uMwF1su+fEGXVCEHeQkXhNKxVFuUAy8aPn/TIdAFF8CxCqlBZRhn8KtUFbrjqCqsJUMOOhaZbZoz
jTfqfaJ0R3RYyzA55c0NSmyCfMjGzXcdaMIqyQVNmVrX19zkAb3n5UAFgn+ngQNOA621G40F38Tn
hl02ONBUoKX/xB8wWhslvHTiSan9nsA/1bxhL3X2SSFZ+uuUEPHtNlR6LtduW0eAjgS2jIBqa3LV
5yFGElHL9X7EPzvScTTXfkFNTUYOnedqmw/idV9rEeHNjODOo4SO8AlKqCHUpdSrbgw7+rdohMl9
1/fO/18jUE22fgY9yAAtZJ4EdThuyj8dNqPGwZ7RhqSmEEjNtST+ek0YUpNCK/s0Yzi+vIfDZAcC
VKHvT07hSq4rL956XuaY8cS8RXPh6M+b0rHwkBLwNL1ZX08E31xjJW4dENEw+nGO1I21Ov5+R+Ix
XMtZDUBPAPiXX1zviEi6w664BpHdoCe5WCjWGT7Kb9sewwJslHBXoO0/JME8UKS2+H8sQ59Du2gb
YeyuXmWHFnVeDKBTUW/9yeF2IM96DJSnZTcuflydHjE4CkuZfkQMHPqcp1f/281TDLBXdznSrh4Q
2U6nodWRFHLOQQkplomOKayzRQzeqoJWmxlK+WoghzaDn7Qfg3h66LLXSbbsCBskExxIYCmDzKn3
5lZ8mLvJ2nh4Y2yVx1xPguaEiUO1QBgsAbrw+aSMMkk3NjwmftAZmmv8BZW4qsmauTW2YNJEAwc7
CXzx+iW5x9A1Ag2oWYMKiIlS7j2ikedSJvFXGGDOEhLdCfGPDRFJJsX51Bceg9cUJlDkEZkV4f/1
83m44/z3AJpmvcRI+Mi+BWzdW/CycVJ/fHtm57d6ihMDa8qmxGidvvm8UkRwYm/ctPZ6DEy5FXWb
9er6yZK/uiKWuJ4gwZCZBfEU1wtN+20TZLZYoZejWJ3FCIR2mURLvnZPf8sq01jxsLSsjtyAdfR/
0+vmHw2C33Lp6Bsn3usf9wDEaCRIAoUptRaCdktuqONzOopEIinQJCzM8cZ7udX4B8ZsWkZvpSOl
KA9gN/Hjwa4yK30r957F/BOHkvBe1NUQcaGnkv95/yg7hMuwCV41RTE8Eme+nncOtNBWcNdNXDd8
pa/06/0rPt/0rct5OLsudH5cohImpS7J+ZZXFZ/NrofXWm4Gqfk0oxwPL++/wR50uFtwcGb0cc8a
L3k67+u+VpoLCam7ieEAeXSsTnglBar9URaWfOS9tf06lNkFsA7WxL+g4Si86aaF+/VmEuIgNvcT
j+P5f8DN8jqxAe3ulJmYMyHouUBZtQEarl/v2D2FMxj4gPAi1p4Cy30+XWLoJ7dcA/qeIlaLUpBA
UFiOE7YqAlg7ZQuYSNLlP/hOIOaZSogQ1eW/tf3csnJCEtGNnkKsy2xxrEs45h18VITgPcQg8lZF
DZ5t4wgfDGsd/5WOOku1vI/DtTKdf8tmbmYa1JPkAFB8wonTe5y+25YAzQNg6tkxJbFNuqOqRQvb
2g3PqI1R5aqQ4jM82MSVd75PfWizlxQ5btAMWt6lOF1Fo0i5m0fEebE/imlD0xSaQ3w/5xg5EsV9
gRftB1B6wPKhf01yoyj06JgpZIzeKY9awYn9jvBURiVcksgMJkr+GHixhI+BeKxm9tqKAsLxnNNL
XBRA/JWrERt/znLfKzp1VZDlYvaFfj0LbQE0KIuvh7j8XpQjgS+WRPSVF0YbD0f6H7SlgZqLRDPp
oZ+oo4oU6Ta+QRH8IKOaYcWywvXFe7720jPoli6Cs23x3MuKrdhteTa+/NP6LPpM8bhE0oPTc5KI
B8iP/jYk9w9lT/CrSM+1XGpFH54JAqFuIRY+jpG6WTWTf5b1A0ZfOijahUr5zCcWEZGtEDyTiBjr
j+4V33jZZT+AH5q0eExn2EMR/p/mEClDf1X4QHYvX+dQz+IHoYJNrMVAwXIBUQ5J1XUHheVopSzw
HGtA9a2x2nYT+YpukW2m0suGOE/36NmyTaFvg8esE0AJgS6uwRfUdnTrA8Dg3TGvd6EvEgdedo12
yJjN7nt1r9BBHloMG/wzo42AJoEWWt2TolFfT7CItl9wv0h2Z5N4JSlFIFxhOqxsrGB1PKXuQP4u
5gd7t0+sg9OpTqpUnIi2aT7sfxMyKeVeVA4HZNdexE5Cog2SWr5+OqUEJa0jH+cdo+YAYXJynzHw
clI4Ly2A0Jz2m6Oo2IIhmcm6v2j/HH7GUBMTa46jzhGVzQd4C8VmbqGcgiWZJ3n2OrzO636N8R5d
bHaxCsOQMpb3XRxZy8c6ALpBt25DBCHt1IglZsglPETCu/Z8j/28qHMXjVFXYSnjKgsNSb4eiUPC
01UPYxZDMhxoBGm/J65AGZxyTu7BWN3PonZv6nXU7h59OJNPo55hlxTJigfSI+1VV9WXp8flhi9U
CRIWHjVqRVCG2LSQqkIlLjNH18d+3EaPo0kXmGxSAlKZrhpepv68d95v42VRnJKirf3OKXNiAT8g
Hj2JVB51/888OmswFaAKQGYnOy5kRP6gqu2b7qhyxIqIb5CWzL/rZ6gbqtZPRT1Djh0EKp1o7NwK
I9qh4zcPTLlKeGHCqcsPoBSKaXs1nCTrZI6S8+N8otu2C3hukrPeOdjN6zglVr+ivWCRlw3nsILd
xMkiTA37dapvbhLcspEm+92OiQ/inizI7NuiGFc2kbNS8v/l3/EDhFxAekksWJhAmf981UoLEt2K
eU6D1wa3TwAaXZ7zIJ3waTlsKa7iUxzL3N/5jw0ldS21P21WgMsEl3wlRjZJQzl296bO1+MZyUvR
TbE8V16tQLkGxYOD1uTiIJ4NDR98EHEBga4AoQrWw0P5uOvv3aQNCPGUQfhNDuhJBTtgMch9VUfv
FSRy6n+fNVTc1RsgShqlylP4kdpm7IJVfkoQ4aEVfesdwdsE5eyYxhKIhs+T+X1n4FZvFxAY8Yai
NcC/f1XfbUurFzUQU6T3icVgVwSIGPraBuOn8Y3tcx6gbju6QHnP910W2BpSGsgJqLo71otsMFDK
PHATohrJqz0fo88Jyf9OTjHQOqm+F4bLAdncZcyKpQZMjZrDgP7+xup8o5Kisb/sfomV8X/sXT4W
cL2c3IyG5ZioDbU4lVd+Gye1k8UPDF7a/r494Fl8eUfPkQ/x6Ipg8pXvPtET+QYijlWng84VUuXp
YjDB/dp5ER6qFIes5KNsjCvpgLi0WDALTDcdapW8ea+gPBcMbKGTbRAp50brZps4eCDDsWdkVEl7
34uqY2e7PFLAcBZdG1b1/HYDt07l8obQBRUBUnhHdHZyGavwL+BZfxGF78fp/bQJlfiXjFXaysB0
+wRmK2CQDQh0aUZGWEFCGeQskFJj0u8N+2MRcpEqzmY+0MvdTrs9HAfCJdIk3eF39giQEeldogLg
MupdaOPi68a5tuJakXjZy/bDG3wx77/3Ob6it26pHewS2uCs9P0nHctdy4R4gNfBJHm7r9s6YI6U
RkVjJAcrHjIz6d1fuwKoSvhI0tCwcVaEPefvHW2jn2/Wt1Mp4lAzN6BGXsY6kG4iplFD3LKbQUBZ
QZ8nPsTQFObVNE1YCqzXn6NLre8s2sOS2ic4iU7OPKZqluUTXIWCfV7HiSyEjrmdnDkBF0LSi70R
lKFEOgAC144AJEpuJSxAycHdbIB6cofKE7TDw8SxbkMFAKstwjUotKy3fCkfkcQtubZdXCe3VXH4
a17mRjyWuytNdMVKe9q9yyOdoy+FzA7CxJYi/S5/1FASSiTlm3yug+DZI7y8fp6u2DoHsryAJVnl
1jVngFhrJMAyHh80dYD8QWSzxjFPDafncldsubbud6Eui2pXTfL2niJd7EZ6r1UCCFDD73R9gNya
3RUMQvbRORFtp1MjJiDBgYw5qt58OxgMWst1q26DkR2ZdBKpMiqxfQsYLV1Gfbp7fj5cici9isps
4MtZUYo3TqOqdlA9UZO7TabIZX8CiHdldsEL4txEISKrp9126T+VBj1MqMBC804UVzcRbLkXhsQI
RykUZ908/PPjG2K8JDbIyBiJ9dS+J4a3I4DVhM/Wsb/FF/FNkHdyiATD31up7G37m+vg23A5zKwl
SMrVoUVdKJkrNqQxsOHzppVFkNi3Id0U81h3oR22r67H1Cvd6GDqvMvaNDCSs16usVHH0Am4ocr+
+tIy5qWu0kx3ODGRum3cKw7wpzOWS61tec4xPz99QwOU4qwYsvuUyvsipwDENrXZeLl4mNNmsZaa
lDwBt9oBwuTg1o0beKHwqCQApsJwzQQmcl8NBB36uDwVD8KO/PYTns2dEwxlC2GWZtqf+4HCx3rr
QRWk1fxHjKtQ7AXzcaVc4wDduIC1W0erSVY9M86wjFySNEfhz10eY0AbK2q/0ej56yz+IaBJhrAZ
R/+ejrv9B5lh867Ud1Fg2JcDuGk4Tje0JvGd2z3P0rZGR0SoLU8UTzRdv0auSHZ/uMmohr0mHdYK
ZdiNE0T10dAWBtVfO8bcga38McaP7lJGMik7bpF0i58mQhqMrkuDVMiIBcBxwGfpJYTZJMK1/vDb
4SIPdMrFUKNhT+znMdjMciLz814gBrPjdBn8U09yPRwKhyWIfqBi9GkcvrMoSfArCeiXDNdx3fj8
NP8NX2EhjKunFjvV9HOMC8bR/56hYgE3nPQ3kwGdR/i4Hxzk/OO93nZx3pH8DfKpFIOTZ95Cs58d
8Kvm2g+g2LlqOSHgAaJASarjzMVW6m/vh3l2orZK+dr2H7qKXtR+54asFW9UakrL37H3nj2Lzl3j
ana1Ck7g1p73HRPaRlGUu09SZxCe43K5sS5O50y0mQVZWjzcqrN6rtIGvCTJ5dfIi1wEnOUX7/W0
0hxa13NTnyWzl9qBa7KBBzrrZHVGgFWDq0oVsOTSTHDkR0bQNi8Rg6U+N38FL6xtB+w+zoMC1Ep4
Txy6FhazoiWvQBDLhxAuaHG2cRjxPloNUDSgzj5q60wGK69IOymEmNqNOQh6TV9NkROae+UwaVMx
wHKDURBC58Ngr6REEXdG7+Ct1Cv1Fu83dIawVsEPVeeXnvSR07j/b9xPAdor3cExdItuvXnWKzaT
Ppht3pSqR60z2FvtT2BrWbApEH6QyUWDM7l3rvviyznok6pdqjowXbZ7/j7LQ7CyesS9yREZ/B5b
kjc2RKzvbx37hQ3yZvnWMLLZLCDUfo+Ake4+SdZigmWPqbqsCpf1m+maMR3ZUH9mSeLZ7N5wOiYn
OKCDVP+idzZsQ5fMaHBNYdwxztAc8r5m9OltQ+n+XaWqVNJCAZZRIuFOA4aVVqy6/9aco2FukNwg
NeBkcESA/wGYwwKimcFq8tg4CmxWy3dpWBB+8v2QyJy5lIqNSR/YdNFOvSaBBJYlpByqqK6iccTf
FV/yhyAbFp2dMDWsdf+azRimMPmYAxh17xmcPdQv0emOcmDQ4eu+1HvF/4MgLLWTsKi5u92oSpi9
rsBEAiuGOA3NGIIop0I3JvRmr9e+Pk1RrHcT4j+KtpnDdFLzrCnxPGHSLN1Nv01yGiH0Gv257eAL
sr2h1ZifE7XIgfA3EZ5/qUqdcvVLLVOTH/3LYgVpIp+QGwFHcfVL2ubmVLNFmPTr8vJ3a1u9/IMu
hxcfizgE+agUsrY9Dh1V5IeJTItgbQqwmeI9d7ATb56u2d1bKUT5DdURlTZOf8Bkfb09mIh3VIr3
Wz9lhl/NXmcCdowhHo+DCRTF4Op18qRMlqtdHjDEFu6oox3lJMKCltT98cqcG+qIUBxssLlpxNR4
vjMPcGUV+YjzpKHS8Wx3z1z+x3z5c6XgC1cGsFoOqkLZb4YY9cpExueM49RhnJpyR8+n2hhi8TmM
EVK5jgqlHebGkrW4vmqMa1H9PST/vs1tiCNCIIAjpMn82qw9m/Szj8tqYnH/BbMFIKx1pdgeZMKc
SRWoBeEW03IwGZO/AnqbxR//Gl+VQ12plbA2JR+Azdlm1hS1jqtWoGeHeJV2E9YRMViEpFmWsNip
v3JpO2JlEyo7mEDbxWffI9HRZqO49lrIrGtNkP/+0qolzAtsTe85E398HmSjBzeYowD6AXoyFagB
W6XzbXV7LIHqUqCRmGWzW1MoXT2s7DWDYqzMnXHTO6Xt4LBCNP5RZ+prl+hnNmK6Ewquh4cvDlVa
lGvjFdJvh6ILIrMMgdHRTlT1LSLeY8Sh6wJveSuljofUYcxoDu4kSq1Zr8GthzwtXUIcA5Xu+JIM
aAggHD7+MNd4V8U8MqtimeLWsWIUk/AAojMwAXp3xp/uyxO9y76cncN6WoQu1NYXqtqlx82k1JPW
8DvSIIzIAItX4DB8XF6eV+rsKZRjBmcYL/NLH4MhmCegRUOcs2h1+svLFRiqfBjxZAqtm2Bh7Po3
AYxut9zEKJVHVIT1Br2iMAWsDGAzzc4HUf30Uv54JtM9HsJXF2quXaBeaZLBgFKEtBMvYktpUVFf
2D5XDZTTdHq/xxGOA9nSHu1lXQkABn4l04pHbN3H1Q+c6I5Gl2g2vNCWOkQelPiFo4bv+4TOm1z1
vIp8gclGvbUtjSXwdz/4AzrUBxJXVIkyw9HJ8xaKS1CJJ8h3qggzlam3B9/XEjEBTT7m+2pmNHTx
TX/jLAM0mLUeM1zMfV3VLmbFkOf13Q5NfPxvBziZs4AiLYqRyFgSXxj945JwfGLQJuY9R4gURm93
wtLBo6tF3fzaOwAqkd1mlfi5BtS1IqHhYs0MoHRUAwqKoDNIUlgU08PWcG0MSBMnhA+FSfufyBCl
pH6RzQsbN6T1/DS1WN2XOM5jiGABnSzUnbgWX/5v2jLWy7Pjk55cuPtmxxi0z1vJ3TDXXf3iuEwX
6uX/5wkTrNGNWDIUv46ElINJJikZZvocC5qFPfX6uVowHBv9bPoBd397oWibqij/0tGdGXPGMQYT
/lOqpHMVDVSSJCjd1Cuxl31hhBSyEmLBePEAihFMEBa+bBKtdp3BcnrTbTvDybZMpmTSD5WW3kPk
m8oueSMGgGCmPwAM4KBlTCBwpLO3iijrN3qggDyZ6OXJki5d7zya3PLBxv/DM082CaYWs4za0xKG
RJyy5Sze1V7HWGnaSpT9uXX9B8R9uRUTuoeUnxu+h9uAJCnfmtVPNYLVDru1zSovXlPkCpq4xHEP
TxOD5CvaiRHLWKCoAJxbPVxSL733S+zUOH4SobiCXlm3d+KDtqR9UJFnkEeRiu20OY9JHhFhe8zW
SEIMsleWl+HOo8B3cAiyOht+pZJ+xCyMDgkoEsQc9oxi/17V5uozo4W1ZW6MgNRT1+ceiaJvIlTF
hOSXqOBEiNugmktjj6lLVe2rZmjcOX56MmU0YM7BG1XwpoIi9XcVEYFI1ophXkEij0Z1UXxBxwPs
Gf79nREjDDVaMyhavD3P3di2MXGXAmVJlUueK0Tvf9+EG6cMmpImlY14UjURLHCeLfSkI0PGkypg
14Ihsm5C5E3QAezzV1anBdtnZLSanBhybOqrQLHurFSg22gZdxvNQtMB9W0wj5u/Ahouu2BD1Vk3
kPC762Y2kjCZnYjhnGR9tThgKAIgz2mKwQEbDAMmSZZv5g9YT/kq9loCBf43CG6NVnddNhs9RVdR
fENtCf1oeclNQzeX0x4/GgzUgYGDwyQXeNaR+K7NZ32o0niny6juSUZ+b/OwjNd7X8rbwXnzZce6
8YoGnzH51OtU1TELt6425NThuGVOlAghRa/FKCPkV+0Kc+uYOIwmFsAfIq5nuhqIzd8Gyo9zXYlZ
szWKhUS5BpAiPe5+mDSW2wJx6rrSP5N9o8N3AKlvyp5HC6/hyYoObNbMT8Phbicb7s1wGA/tf4FJ
IZgp55CpKIKGezRGLzRHTPgMcJBL/9cb6vPpup4G9r0EQRi3dYUCljb4/1EMnhyc3GYoFH9FIao3
ihj8QKILUfNY2fxvZ07aOAlkrve9y82+oao2uxhMTUJBDEXmcq+M+b9KfYxD6F0xgC77HhmYcy/V
m2jSaxVeYg4KjdWrwcnQuzVeZHX0PCJ7TpKRx3ZrQ8zLL10Ei9tgBnI1q85rgFmVl6g9RApQ5GcK
UQXxNPQdJcqMYSrxsJAmUFD+SJsTgbftzSurEL1mNybhLW9dpq8WIU6cphlsN+5VWczpdHQ+DCWV
coBXyO/HzMseEjl8kSRv+gd/7i+w8qMxjWg8tClDNrGM3Dl+Rzr75iroOo+lkZK/i+qvscVGM+KJ
yhE9e9ITRVW+hpdmsi4QmU9wbrTlpJ48qOSSJvHUJrpoF+uq81QaMpJ8TESpBWULURaEi16sK4Dk
9MX9PbbrmFaHo/Tfn1ijpetkAcC5p9PV79j2kGA9uXgr+++57TNqV9tJ5+QZrvExn9TEIkb3Cori
XAPT1OEeya3sa/acPu0acaW4YrbPGE+MxzKxYjVIX+5v5TLVdRIPqURtlg4XWzuBxI/GEUnWvAhS
7c5Gub6ojCODzxQEGKVbiuqwDrHkqYGlrrbCghbsxPTyhDS18hKa3z+bltLOAKhb+qavYR4PxevQ
3n0LHzuviKj4/b26Z9GuYOisBP2QKilNESuEXcqUknlzOl5xZ6Bd1dPvrrAW82EkUUOcHrCgylNG
66PeYZrZGLlYxtUuOECmf2HC2M755dwk4WakL/idF/iQKdNYNywVGJp0GRhw1foXuyqntxH15x9H
Fzj5inRc2wMBqNL1z4dUEdANSObnIIJ2o22uj9IRXjQuV9H3Wb1Eis8cqllrYlqhkO9s/1FiUw52
HtUtEZrYvQM4/+8tRp5Td8ypK19PvC1TkWFsn0K0GfqPedTx26jv7DSX+0t9FXwi3X8bp5tBOxJz
3bqzlB6d8fyJkFQku5gDPhcf/KmwxED34+SUuO9m9DQN9BbWZYyN96gMjs0oG8EblSTrSNesb3XC
9FJCriPsZjv+Hxh3BLODIyRhDzKy8Ebk6bFAqgdm0zBDu2wM99UHR24DIDzX8xHsgQOZ2I4WQ1HW
A9a3KMDkaIgTNPH7OfqjTBZeVZfdLzeraDjKdC00pq5sAqzqkGfZXqM72+Qx2Bs2g71g5eaaaUKX
9y+u3qu++21CWkdNdbAlY1u0stJBD71pQpcHZNECZffzmYsegCq3pIhfWnb2865haAtpCNRwyepc
FEKHo0JmkDI1i8oARaRBFNHLl178+jNTSvKS9d7NAO0jz5dQG1ZjcMDq3iNpvMa5YezYcQtFf0i9
S36FYkXfO5FQqJsGNUkMYIZ+5BSj2MvfO5QoOsjbDaNYfzUUOJpaRU1EeHqo6nCcMzdxtx9fTw6K
aT0SpCrzeW0GfrT90zqpIjrQ2JFZrU9T/4D27MQwOkMrr/u6H9O1hpgwMT6ljGe5x/6aD0Tz82t5
xMnn7f47RPiLAE1GzCozyNhlWLOT9nlXKxRC3u1ZLvfH5XgUn2Sd6+1RmQfbGdoKI9bcp7OkRAPF
WnI8LO6WaVHU5/cArX+gZBgoACTuRYmeHxDtMaltT+MP5EDWK0SF8s6EcJsiSD4rhzDOM/R6cj4r
ggOx7xvikzOwQEIRBhsitkLkURLb3l0agFhD+g6x6qv3slazsTjIjV/vuxY2XyNC7X0BBJKjrY4b
vtlJ8yrK1svVPujre3tSHo29+r1RX8Db5d4d+3p1o4Mwf/JG7FwQqnhwZZbFblaXwWbmhZ/LqQ1u
z407+gmNMGTcMl2p0kycM9F56YeFzFE/VZASs8/rD6cCaPuLtX8tnYn/m29DKk0ZCCk/LnV94xn5
b/dcLVZ1Cckcxzd3PWyJkviKxH/NaUQo+64Uy3HzCR4ARdVD5Rs0KObNTUoTnVtagfQDRrUaRzFg
Dy0nGnkcPx50wneyz52iaGCgKuZ+mvJKj5ocs23HhFKyD2XqSxVHq11XwJ4uSMrX/M+G2v6dJrY4
2gu/PIPalpxecYmkRC3IjsTVncD7ZKKV9xA2DGuIbOsIoRFm3JvtgL8lrLeNAo0PaaBPm5vdWKAP
uPdhivSGaEI01zt7iIH/46dpaPFQACTm1GH9v4IWTTNQ76nU0bknD3HIAW/8k7fjb4VsgGsmT86h
stYESxMs+zGN53EVAqKKGOv+bbOqZKR5zCbnE3UTpg4fVz12fe8UBOejqwYbCVJ3Pc/Gj3wcIfCv
2QEe0W/lSJ6pbGVEZkpeS/tU0lxc3EwbzTSX6IN87BjfuFTiJRlOokyWWBsGtGZeAntvRbpJdHKM
CUgJrJKZGE7mk0D5NUFsUq3uOzIm0Yj4hPz8uqAL2gHVluZjj/bRpSySLjyHtzCLbIxQssuVQgbN
Hn+1fEPllOrfTO3jIv97eewKzbqOu+f2BWSYz7U27bh5lsy5gcfX8b123XSJYIIi9ToMUL8KIdli
aheJh7bHcRWqroYwuVt9XgSDyyBJIAgv/2xhIAiVs5FZgnf1jGi+Fp/bdApcSKc52BOPf1BS7WQQ
wTrI6hJzvIafRkWloRcwr+5pSFcxKNBZmgJad82+N4/GvGOvNL/vmP417QP5wgvsstLBKfrmTmji
/hz4CmyqJ/RZzDNKfDOvSMT5jMV7uWWk1ji/GlTqtEollZ+UeGwS0aA7CiINzHAfmUv92BI+To6H
7ZzSjp2x77UluDlYtIeJIGwDVgQiit80x3YP2h1ot6x75V5MiFyMOSaoX/hC83QXiqNxO01gsi0Q
GNqZzkN12FvegjTGOxpdxi4D5TtIVxisTTpe050XZDshJJgjRFGcaHs0TuYte6UQPFjZxxaYKwAJ
PQaMl/XVzB/6ZBgtElbSMxwHUzSTwNKmIRgpyBmVYBdZGN5bRO/s388OnxtVUI734cEErjRhDJ8y
sT3bgLvZYLtArafdIC0XI5qijBqkmQpWIcNz43Sul37ihYfGmfRG3XSQsC3Bpw2n9QZ7WVgWrChC
q3/JhWsD6WcagT/fNEwxfBEn0WJ6V9Z+ClK411Cwm2yvZupjeCUoLuAFaP/KpUKmSVkSvauwB17G
kZLNRKexsYONiQv8kFLPGetpOuUwy43AC7+tEfWcnBTxZFwtt4sMJatme+uXsU4PD08EFTVZFji8
e4HUVzPexMkbk/8fnTw/f3cq85aewrD0Ys6Qffnn3PwWnJRyUpFBsxAxcox9DAsNkC446ggpJFyQ
DTF4XPkfPl1dPNPsJ0WlZNYLRpmnWEGC/Nh0lBwC2UdbgF8/sWf7bQ7Llnx9ptRk6laKj5mvhnL0
zRXvqrt10aO2KcWGlTq8CsYk+fo6soGxqIounM8BWMdACZuj2ZEmO3MN9vqUDFXfsIk+q1bhqdnr
G/f0QFXTkhMX/E+gAF1Tto7SYNcSyXb8VPwayWRPl5UWvJz85r6rpWAvHymboisPoU+7pPwXu6tp
qWW7AxHUDzDlKaTIbptadwrKh8oJxHjKg1mwDxpjeKcfh8lCNpkj6ci+lThnXz8IAgpfpNZ96scK
FYbYWD76MW1TWM6X5jtc9Xm3KQad/NMCouPrV7Z3oSa3FiyjUseYQ40LCD2O7ob+yKfJ2TAKHkOx
hzqvRvM1LbAzJHptC2OLbIX8+Hv3BhSLcuHMTMpajVJBew3oPDHaDC0cyvv1sk0NpxaaspWLPz0s
VdMOiHHi9cfNzFXhM6r5xNzJESAuiObqd01bWG4zDYQViVyD9fPOqhIqQccLJyyxKYQk8L42+XB3
6pJCoNVLSysg+9VzU4CML0FhmLu33KYyI4PbHaoAU0QMx+ZnNrwEmv9VBUuswP/Z6Pt8rzVUf0En
fVQCnsZK1yP21VUX4kkxfOrvbpn4t19s4oCzYGlSVCOSn+ewFz7qY+WSDUnPfykm8ntpn2/l1Eo5
vpi3IkGj/AvSHhmn9EYHssQ7IYWJauwR/KTaHjMEMdjbXjMbtW1qFSGVhMigE+Wq51R5uGj0DEF2
k8HCmUYJXU/hotv9RQW47buLJKJTgsGNjbAP1T0rHekxUf9g2hUJjNbolkaPS/2IqBbQR3ZwAIZI
GKQ8jltEVnK9hGd1cEHB++uT6VOpJ9b7UuCWS+U3CS/5D1wqY7lgFu1ZpBFRfMkWoAAW615VUdLR
KYgYznYp89+ql6ICIQRyQD5YOQB8Ea/tqE1Ysskt/GyApqT2yG6ypVankcogTisk8l0bomwOTmPW
MwOuGIxBqq54jxhIHOXCpPU8HE73nk7Th8+sN8zLiu01m1Qn3k/Y5XUImjNccVg6kx0Jyb76GJP1
K0T5nWPR0BXOFevCF94BL1HnpsEdSPqIN1jp+9RHwQD3h0QjCY2zSfw9HZKRpzSgHI1sw0wCq6lg
Csk0ew86gYvpzMK5WswUVWY+ONdw7ixyWWVnRmFVWbvK9Ep4OnNVJyhgqrmToP1DpYlW6ilDzdna
mltvyCG//c8iNiHpvYBlsGDmFE9sd5TnoBppXXKQExJa5DXl2+/pSFCUtqqS+nP1ME70WBt67Oy/
uvUIf/97ckVRqJPdmqvHQk63JUXnoCx8tNQYERKoGYQ1Kv3FmUEO0K9K3d/BlvYc727Y6l2RLgOm
K15V1JDNTnTBQ+Ks5o7J3XDXHnT6EmQDL0E+kEbR7wlEDmU2SAixFqucoNkJC6BzIyar4FsOUxSj
1yUfZlrxE5h3jQxvEDGweQWcVL7KCQYP4bW4sL8wizVFZyrhwIOVD6A8iUuE6gySMApFLSkbpTv7
jrJAxlZTOxTzNqPfewPNk/iIp6bpEZdSIXjE22tbPy6TKmUzKfWGISY5UB9jYQI9rpcswckk5k93
lWwn1FXf7oeuP+IHlIkeCnKkVOqzNPkqm58SIRT/3102MHeRnA2KB3UmLEFx/dYRZrIGQEjqWsli
xbB0X+XgtBh/ZnWKYkmeuTuBrw+A6mxxEaA0UNeRvsmTu7iZwsFZ/zfmQKqNFAJP567NPKQGYxjA
2FZmN2tuRL9Y2dkDUAHOInRzsGI+na38lit934McmEKdA/REVMK0vWAtuDxy30NGq2W/W8HmCBo7
FdhkHRqDcxSFvyXUoAWjS2fIPJ4g5U9E5l5ugwhQksZ1+Tu1l3VvorgG8Milr3j7/oVJNiYOaX0W
nN6EFAAiKxVUrNRlQLXqn21Vr+od3NKdwoudhkhafTAFY+5ZO9priARnY4lwZVLz6iRQx32VviAQ
jFSArBvCHlRFl27fBWQ8707f1S8Lk4I188otvKpilzO1nM9Kf4I7mKA9wkjsTzIbNCB4N5c9LNYx
9L5ydT9q5CTZ56m074XBBDMGoSEgp1yFf9wPmv97Quhjs1xAhnaejCjAjjo4PHNh2icFmTveL5HF
UTOp5nRPWjMFagNr9B9C53x9UHIO3Moz2Dtk4fkiCCr9B/oaLiz/WKZ4zJK5HY6DQmV6kXeyTXcA
XtcRHGzxrMGWUVOnvYbdcTgOd+gvRHjYuz8ekSAFqAPBTzQVp3SXFLA5puPn4AGeGWFEfh+bYLNz
wFB+wjm6L2m2VKbOawGp4TQ2GorolS167C7B8m6cChxt7XzWNsPWqcoLdhtcEW4cHEJ+CvD5YlNB
bSHjJGOzrYSWLo7smVbn8FO7ZoZVLuoJ2jkKdAALaEYyDFaeEOmgbyjoPFPEhhNya+74k2JH6JjT
snjjAj1Rgk3iuoIBGMgZneOVP8JZ/r8t1WSQPY78HS6/BOUFSBA3S8e4xnSWm/aNAiY3/0G5ewPJ
KbPvmYnxEMeZJBU5TEYUx1+5xWRG47Kmv6jzav975DoMdLzDkKVncKtEXH2ky0AEq9z9hRKXdaGm
0a9eCIBUuXR1sQQTNAP5D8Y7pEuv2UohMB3trLjTZnC5tG/CKO2mxQtPqJuOJ1XTNHB0V2WueEM/
l8cW/bxjrFn1mKFIAkX5urVY181tIDsjzPuac7EqdT/6pWITm6x0Iucgz0QrKeI1EDOnpR7Inhfr
3rg7Jlwagu+OuCxIKMaZS+7an/JLl2Yxj9FK/oGfZvnFmcCxtWWRxEWM/cFD17U2IGFquFAeWjDj
nkfu56lwcwfGYUsRpbJ5NqTj1j8459/8GojPFFdRp1mrkYKOONjyHIsUObhfGgpLhHurQ2hVjjMG
UJR3C2Z4uf/jMv5D5ZlmVDcIo37XRxZKwAd6sIsJc53hphggYFZoJocIxR/s57+uh1V+US3FX8HW
Cp6rZAvIqR+bZcOq84Kk3DNA3tYQUv1zP3z44cj6Tuyna083KWeawwz5i0ALoV+0gbcKFnRBQPZ6
H5PrvkDus36ODOb6+YZYLbzxhhcipcMnlc8J6V0ocmxynmgNCHqRPu/h8ZZyaPRN0vl8GXq1zbCD
7FOn5BFCpw0bka79my8b2W28EifFTciAM3cCLpSATq/bnkH8NbzpnuKAcH60mPluDKbXsk2+zurp
duIlh+9XWPjMGcCd6IDAgMsoZqmX9c9cpjWGPfRGRAJ9qOWTDiClLd4U/h8dyEe3jxWsBKa084NK
OxdcTFN7WbwvxE+ArKoY8nd2Rhhk9H4k3d4KuWh62yWpgiyQXfAvCb0E1yyYlE2E/V5oT4ppZM4l
QrNJWDlWIkrxbvlaktOQ5vf2X2G92fFMbDTMljXk/746Rxxqk9t1gLSDxTfDnsvZKB3rcB+BLQzO
H+pRe/94Amy0cmoKJC35X2ym0chyTKWdXFHu4MW1i2JrMY/C8zA40Utmv2oQNwyv1bWpOeM8w+xw
ghbrYETrfR22n1F29njXRQOBRP952dWfnVkIhUOaQQGDblA5TV8ClFJJojfKRobHs1KOLai0sjqz
lXqD6ew2JjP58/eJW27UWEnPh2raoVpJSQxNUfUCwTw5ofBmlGwQhXvli1OpVtwXnJc8W3DlyRtd
X+j3sbIOqqP+C2ymSk9EftoPcJ7tnNsj0kdJ232p0ROQAPV3zhfyfFKuIqVwuSQsELeHL4v+Q6MU
A8mRylusvysd8EdCELeULEeAmEyZmXEMtTIDl0Vd+UjLHL7qjQjzRRAPxnSM9wL2XDhr4Vb8qeXF
Egq85qsAdQCKo41UkV4Dv4Hrjc67AHKaWlnpGy/1T94qcCxI5UPb0wURFvN0k5XavGw9Rpt7hL9b
DwpN/RsCmJ66GsGTFy9pbd2blSj08BFD3shVJkcwjlbn6neaG90QYulbtoIMcblDYyfBwPgZBbnP
1nLo2s3s+21BYpJGO+MiBx3e4fIsk/srI7wP+hoJdI+rnpY/Vsn2J8uOBuRmgFusglLaJ9b/5YhQ
SFD3ox1PhMY+uhF/SbRQEr6cVCrlISajk00ZzbMscrstidq6dgld4/rZACyflzMD9kGukYCfTD13
czuO5dkG67hIJvd9kWZ7oJ6ahc+/mBzzfNj3SPpV32n4KitcMkrAc4ERAEWUlXGUYotQr+oc9AcF
CP8vvh6NvUNOWzmskXJHracxWCHCfo66gxXMTy4FsrQuSLleyRZ4BwwWelBM/cdjAfAiW4ROlZv3
s+njRYNJZQ++M22m3zgNct+Nbc7y8X7696IK681UgstpISjPWMx1Fte//IESHbaomF+fFVkoHtxT
WqjdAGlcOWepKrL08V1JiZ/gXpJH6reru/REpt2vcL1KXwjf68iIXCRTd+HF733l6y+lWH8eaUFq
tugao/Gf7jhTHf1yapyVvMjuhrLPEO3QFgwnY1I2xORrXPFbYJ8sTvd748pm9LxVhy3T6pQ2OCl4
TmwP+CUo9QMJkYdwSEviKu66LaTjIrz+R5VOl8nzYlOBGoH86XZNIAfNHKiDHa0VsaWB2dWjpNDi
BM+e2gEGMSz1Wh+drnxRyhM2y6yCQR0HUNlSxKtIia6KF02gfvYuVhzSU3GG5OvIxXs2NqAZCJot
gmLYgr2d8opax7fm9tCFtFLfpTUo5iw02zY146igejg7o3B6Xp+MBErSzUG4beKdUn9vlRquhaQn
Iq+f9Bxu1noqP/vtFvh6emAzyF4UGH53sFv3O657fw+fuLYmQkS92E/XUvwGPeRH+SyuUaSvkAk1
M17Z5h7sg6zl0oC4VkVGwAb9o1HKlI3WEufS15Er0ex2XomtM5oZhYwCOA4OQlWKJsGTSdufunQ4
HZ5zNOHg38q8UXFMCQ/QVN4IU9WRyYKhE0mcUf6WG8c2FUd24Hbo6dGM5pGBGi48qkUygEFo6GXF
+gko9y8I5s8m0160zZquolhBp54IamKY4oGu2hth9De7kEq8ljY7m1TfjxYhvzSC/NBFWoFiBiCB
ewcjl8acuAmSxfQSK5j3Ngbr7QMJTSQghIIr9ONv57H637XliwZfyLyJDbrq1WIhm52dSozMsAvt
NkPVFFbUm5HjJCg/EC3jYnGoISkaFaw3dzXOKxmA8MY4Zl4HxtVn8kv6dlXpjtLN9Nyq0pB51Oqp
cnSAqE/z3cse++i8iO4Wwz66nHbV98s3LGM8DOmFJfbbY5/M+WZABSmoICIfGT6R7jXq4X+Q/h9m
XchO4BrY2VFXSs7M4oKqzquGnOu2kAh8iJW6vrzuJXjNjFHddPEePooXS4i+CTzU2BB9qh1E2zck
4giW9ZYUtXMPypTCGt1/NzRKKa0UfAJMRqq/7PLyRaKqU4joci+EMwXf5XxqJ7xnfPY9bZSKzWc+
h+wPpgePQkH/f6GqP/+KifCodv2Ac9hqESarCPVD++ZTS7TbMl6/5dZ74HiiKsLcwvSZzVPGFRUR
kH7VIsHuni0xKmHx/u9SC0fXjEFRBH75/IUByT7aiMfaLI2Ck9NyhCFVyjyoOHM9rBvdF6sNlTzC
1Md8jjtIJJawFY5y/Nhho7Gsi8I4uEF957K+f+xWH8njkf3KlMbPzelHy0owyM9D0LIRbxv4qypP
ikQJ6QcvvrCxbfmAwIXyZhToF5aVEbEzOW7w628FqnQjRpc5JoxdCGeZh6lxYZ4q0gJ+bZikM8/Z
ue9+37RPJJfAjddcvZebmItJKMi/gmrDqWCD/H/BLycA8yDLQliTF+6g5mdS10boyvxwmdFCwAgk
rqnTU140UEwcK0d2/Rq1nlllNYLLTHMB8LAFHM+VIa8cGI9AcyJc1dRNioVi6UuqbYZoV9QHqa0f
T6/cqsTcUOX+Zi1JlXKySvxyhPCyTV1O4lut1R8hPc1VFeEudXieKVnbFPSic0iiMFEKr3SNmSwE
uusi74wyxsNNvCgxW9Z5OeUiOMvm6ILV1eKEAYUQDYzbBdh9iVN9QCJq3jjTL6j5dF3aXDmm3qBK
BSXWKaLBtj4uXxanM5q3vzZ9pI9BiU4ZL/Gooc037N2kYgAdWjET3grqbzyeBlgoN/Ap9bA1PxPW
nbYA940kXG/foqcvYRwXocEYeJoG9vbZu9ZCCD8+I9vFqmyRIfx+u55p7IAdmzcRVbPpqX06nYAN
1VEr3qwlkhmz9MJ5NoPmo3+O4coSeeXGAnMlSFmzwSoTacoTWb55WPZLDp1xJu5XMlLbzTacDobE
Xc50Q7XxvD0S7Og5PXtGCKQmWcep0SrXvfZZmPpPqKsVurdM4giE557O/wBcT/E8OmMK7KCoIFu/
K7QQ4kMTnINEpWyry64a+w9wd1FC5l993II8lap/lz5lwTuFsZ++JdxmFkoSsn1f0b8Op1y9Mw+0
+vgPwHIof7SknmzBBvXjUbrFEIINgKS3texs0w+ewIFdpI1eUXob0yik9VRZ3qpm7/48IOTmZaRd
Lq0/SBpx+q2JM1ww66yYKpK3rLojpWPJvw7hIg+QWb3eXPzSN4ZEIVS2iN88QLIxoy1ote8cB1IL
iUDhl+F1/4qoiTZi421Q6wOQ/DG3wpBzPr34I9qZk+A867lAzm7oyaZ0rtPcdAZtiZXCxTrK7axf
tpFIC0cfGZH9lVmwCH7a7l1x0+oBZgNBdvnzTNiFVIPHtvsTHYhEJGtPdk6JzMdozo+XLucKBU6F
bjUK0WanljhFHxf0q2uDjefswNJmnZqucA6U1OcWoLZc301qqAtNAbtyrWJZax9DveapMyCcM7dQ
6YR1WrKix9+8jCDQCq8X/7+51qU2LHQcWDAywUnCBshoCfZIz+lmvs5XRszc3K0Bkur4wwU/oZQf
DRbNr1T//6U1lWkLUtfM/Eab2WdpJbtUYmohSARmA5bJ44zHlYAQV3/Yr6MQjiChEa+a+nTXBj5/
GekYJ2m8Edh+zuI4xgMD/P5R13TMcjrOsBpmNXj8r5BMaWTKr0FrnMWY0JMSsUKl5OCvGL4ZKP/H
5/b4oEJ0jgAe6VvWTxFl00L+ceeWkQFliMhEIvhIu6otw3d2DFWYJhxQ8a/CrUjNuZLAOvTH1O9o
4KE/3CJsxlncG4icvA4mS5Dx38zNvespj04b/cDKca65QKUIk5kc83TvXJWp/AfMvkvaCvXc88Py
0ot947FX1mirubxbMDN2EOgPThYYuO1nL3GfkC7cVKN3STDmNho0ynQ714BLHUtxCAI84hFKtFe9
RHffkDftOFycsWTw+GWTpRg6gLD6i5sxeTAr2CnTbcahN32/oXnBNh5nXkOXW9jTn7D8TTjv1k1T
zWt9Gb1oFeMQM0HZiFH86BaX/7Zw04HS0uh4XD6e3WN6nwudLAxsllAnAsf/84/gZSfulYpjGXqn
wKNtAK1B59OsU6ItoJYjZ2obmPi18GvmxVsnwJCzvpvVHlBmrLvt0YSUTKeU1NvgpFjXTx/LWVjd
JIiBmELeNcToO+TE3vOHAA1NBJGK9aaNeqg19CxqKVIrH/wU385E1p7oRikAYprc1/AX8FWsK0cX
MbtRSLfw7mVtiP09w8k7LCNfOjvT/CxHH+63mxtuDXpx/FOY5oadfvGjb7AudFah+Z4bNA4XQ8ME
ATYFFpOdzjbLO+KLw2lPAopwLcydKslP9V4fClFPG0ERxfdflDoG4eiLQOEVJ76oqNTJyGuvHs9f
BJtrkkHOfFx+S+crQ/IZ+diFf4aK3d4W5pfLwzVYZxYxsykK7SON1/i2Yodn7wl3KiCx7obwhg2e
/ny5XJPDX3Jan0qj8pxzCVBjayOVh1QxufzsG/1IdMZhqfXwDhn7XnY4eZ8AeCYbKIzKCRHlQCpW
Lo9nQzIzKfLlS/Xku5r0v3VuVg4uOmKMrr71M51BhVj2tD1X2IDXSAdRXs19hk9PpCxiXWyGO/oM
C/grc/RQ4uC4+kqD4g6UctXaTHgv3bL3fo85IUjzXwHtBUOAoPdMksEbxgbbb8lj90fblhZce5hP
OMbD6QJCubD0rSy+F7Cd/a7/sShiyudMwywWLZ5/vCUFG8hDWQMtlo+hL/ptD05iUN6sWEaH2okN
I/8OoaeTWAtWD2tZgFZYo11nmjADHDpnr7YsREvXUnB5GGNey24buV9h0iq13Egx4FvDlBl6Xd0V
fttbY341TFJ+Wd4iwfJ2xR1TyXnZ90tTADO0N7s/Q1lF3FeRLVwXC3X9HXLj8rcactEbNLEj1w2K
nV1zER0bxoF3xBLAURr6dz/R87yXOhLHkKAywspKVwTGDg/9t8+nC4SdSAhTzL+HJJ7L93TjDVLR
GbwSEMYkKiXi3LiJpbN+NKwj+d4tWOLAYNQiXyaoEFMgGGkwHQcbk7TNXRoR03zWpPHUZNPk3MLN
94AKW9jGbEFfCih0zKfw1OiqUEcvDFzn/73egKIMcrf8G3VdKa9+hKgs5gLebanPEnM9ujNvGwT6
VpZ5zAPs0yjqeeF9vNLuzW5JE8JIEkpgznRsnTl0kOG/Enrb7EjYozBG8m3pEABpHa02GnQUq+rY
/O9g/0ulIS4OgJUyx8gtyxqhY8difoEZp2nyi8wu8Be9T/DvUC7l/ilNZTD1qSylDguIhh/TPbFU
3AzIvur79IAIC1g/9yIKUpYaVFFXBIZNMogJqITbdW8W8Vcq2Sb2yk52cHRzk4TbU2Dx8/ipTQ06
tBtlp3AHOpB3HLqiUNXKk6gDPDp/WIcILBMYxrDBpsyZyw4jcI7ijPeT8uLHMYq8UoKq+4RucsC1
5VfZJcqDJn4kymelV+Bc/s7QScgaHi4dDt9uAznbv0b0/TELaUeULWNcPg3LbCKvuGfRrsi/EiA0
KIOOFs2ePoWSd+aC0KC3s3IKy3fY6xS/IA+J9uSY2CyZ2Znfgp7so4vKl0M9nmvqTb8lIkt6QdlR
35RTUxnkMz1vtMpmjUqWf4EjyCwxndGCtj1yz61zRJAb4XBwWh1LDXJe56VxWaGkOkmb1JiZ0eAi
MDBFMicrue4RFO9q/NKiszuxOkmTQRQnYERYSS8wpKp9X7yrBvvwfi+sZJzGkBCeVvjDMHRjjssb
QtO4s5wSj20iXnbHOi0WbFUZ65toHG2QVTYgTYBs6HMRfFZvzCmEjg9AlrnPOPs3ilo7Z22N41aR
jLeN57en2nibT1yU9LWWaDEjKABDoOnNsINcFzRGAFza+a1hNleiOOliNbNWglJ82SjiMeoWemrp
sAl6J2DrRmDYVRsjKzPhjKL5G6JytAyWGCNLQWJLScL2+kACMPJlGk2B0ESiB9CIuBCR/WcpriSI
SCCvsdv/dfZBTW+HC+2sAAilVi3zUsSaqsxSo0iM5kYhDnnP2wJ0wTcrVfajO4B3r8wM7fm2l8hs
DJS1CPnXi9wSwXVpHTiF5MB4ygAnAnf1R7oG/p+7sMf0/wrGrgUMQ5WFIkzY7gz6gRKd8xuxy/DW
XCpPOxIBMm11eGG9+yKHGypBYrNjR+1xDQ3UccVW23FPQttgOmwImtb9vqoeGZmmB8Ny4VjDRVkZ
We2EHNkAqT63rYnllgaG4+/WMsk7/ZSbBOC+3t6TbhZ2rBI01QUmo4eZ6Eywhfy5D2CXMudKGj+d
lNrvynD1vUQ3DeKwQQ5d2o24SI5lJp7tlExQz36mAjF4g3ssMXQXJ/MhS+08Bh6pkOBOtua4wQW+
9dDSHeACQrfZTq6BF4ya3Bg+xDKJWX47RR67DQ4v9ezqY1biOZSzDRJXGMdwEt8IzNbXdfOEbOy4
YEP5vQxyXWBxVXlkB84Xvzq8JkXMCaZNwoG5AAt269bWqPw+zgk8MLSzYVcG8/XAZBaz+7fWye/m
PumuWh2oRvxat+//N9KgsIBTrTtqlZLqwvi63IpPpeyCTwNJrVAz67YNC5BwDZ08QuG3X3z9nXWk
33oObUdfj62kOwxzApR+Acidgkg8maruYH0b2jT4d1ALUvax4QGaC1TotqTejNblwHY8/Rz7ry9v
1vxvcQ3H042VTh0kqDNslnf5NsArEqtojFGasV3yUGUsD1U7puIT3X+Ob7pg3G5/pNW+s+h+HH+2
9t5eEBKaGK4nrJCyE1AMEDrhNXYaLBQJVedz8lxPv8jtw1W/KseG9q+xMdnAuYfNjyaG92ZPoRm6
y9WsCOoIkk6yHK2aHFrF2vK1SFQXCIU3iT2EOFLp2dXBUB2wabIF6yNrAcJx2wyQa9w5+E+OI7/1
g0O7rvO+wwSgcOemLI7QrRS/I3xzE2duj0W0NF4ZkCTdc4KziVe2frb1Hf3FQc+XN9or7EcT5gd3
XP/UoDrEdL0BrL392y77sJ3Ll1tepFYFmIF7z64f+6cGgsw9UDY+2TP1mytE7EIbfaMH88TMYLLf
7GOQXlstm7hCrGIyOgVU0Vx62MRblz6ST7y8MkmSmPdlxGW3tcNMufHbJeBGnpdYv9k44SHAqq6n
2maaNc1Vs08IXZnw1tHJJSUqGaymOmrMkloLfs96CRQmMnJwIWZqpF54u9Bxhq0kCs5f1PYQcLm1
Cf3zAKdKAidKLZt1aYka9oMHjTylRXFL5me7t8H6eU6K5XluUUmT+8lFFsZAtHbil1nNL7BEU9G+
U+ET2pYiaudgt9rfD65mq08O1oaE4Tx9SKamO+krVclPfOU11LVYwIWqN6EulgWT+Zdwd30EdM5G
zTIVj68lW6YxIxUu6ll2EscVu81N57oBS7kH4romuS8/e4Y0F9RUvmJaojdnkc41Lj7EV15urIWQ
fhQt3a10Y52Vo05Ssesv98M8oZzyfNlaVKzgOvC7roA0JmI8nc2Rrr1A1UtwHZvxPcJRGklV4wpY
YUYKPHEPmFXZ/6HYaNvqsw/wmW5AD8Vrj6OeJMKiB9y0FnYGXTudIdipnzP/xYYkzyaByxJRBYoj
00M+GIeJSO9Y38iXk0gDBSRssph8T1tR//laqVmeuwZk5mDNr9T03KaPwjjrKWbKQTVRBd58BhIG
EM5AIvwlpn+45G3pCdf9LOjwhIEkZ2w+cHNgFK/cSBwmn/6v34bE0E5/agYSBK9S34samGf+/oqH
N6+XG8z/IZCP+1WXxHeE1TDn3Lp5G6HnnvKaNOMAQt1yESEJqdddGTso83h1JfEl1KQuWRR23Msu
bYXeftgfKXAhaqPLLFBcIR0y667VdOAsnS2vhSWIg7hMJ+5a7HzcnKJbFNAOAwLF0vHZQr7CxG+3
e1cH5WM+d12lCrXSlg3sM8FIq+a7T1KGaMPasMjbfilSMJ8eqoRkdSoQFUDO/CsTJqbKUErculGq
DaUlrP7cUV5NpRpRxJ5x1NjuPNSCgQWAAjFc7kW6M5fhU8NfkV4gEkkWymLzZD8pUjgULZqgDOEt
T1HsAEx/5AGmz90pn/1XwLWYDRA9wFfECIyAzOXAr0ikW04BYmcjs4Hfg8qhJWutCZbzP5u6msEu
HejUShb9yOZKoyLSgqP8XBjg5CfoXdfS8vkPnV4c7JV4+v0ELcrNixr6lNxroWmPeKYNHvY0B5xX
uksD7J4yzCM/+vp8V+ZqdjC1/rMViaJ50lD0ttvEX9GMquVNsrdJGHBBrt6/IOrkUMg629qropmk
eQWBU9PjfpZVShFcS3gfDsKhlM0QrK7e2ADVucL24YMJwwm58zxHb4myGL5iBKSE6bxbLtMSwmw8
fIuYBqMk3Ezv3D9NsnUAe7AlIo2msf36ts2NgIE3j1VRDT24z18POejChFh4uE+B4zzgpLZHwghL
dh/ROJ0UY8LkFl1KkvB/qdD4Z6M+YT/S/mI6SsUI1wJMOYdQw6t16OSYPrT3bR7eyPgtzbKQtASS
gjR33JbPenLS9upvES+alK86kTZTyagiZhbTLoxCJsWUnrj/CEjmNEkhv4CvYRXRhAELOhX00NZt
GwMlr/kWKZiOUmQ1z63mR7nrb3+D333Q4KLc8pPnwFbtxRvAW/2y6AoSxqlxJ4TTdTjvK6t7aLxE
V2+lbZWAZCFS9v0sN/6nFwdF34pbu/3efUtJ+amgeVYUkS3JziuxcXIh2XLrvXzecGKHfk8xSQo7
XtC5kbwSF7H5caLhQtgVniRN+5TrLOrxfRyH56cIRoUtQnBKXPDl94ExD71GHSgoMUMLEt6QOsHm
ElUppw616/dYqtAHRBOUonQcFR3Et/6TamgNNiXfogaNYcwKCcqnzTMz0dCy9nNJyUrCBkl1FWlL
VgbCRRezSbaAKGzm5Z+koG37CkXL0Qk9QGz98k/XfjWKDYV3ZeCWJuIk7fLNed9SzcB2JP9/1dAG
WJLjs3jmUaEL7DsLovIXc9uxNvLHGLhBTQSnSR006UUGx+CAh4l+IuKl/r2+27HVrRut10bqf1QD
RSDDfzmE2pN+Gz7sYTDi40N3WG1a6Di85HIDGJyTkN2zKfcut1fbCYLOOXm1IHX8bafP9e0Bgub2
y/5fMBLXrvgJTy/5bzGKcCNj2Ylyqe/81+WYocrcB14aNHD8igTtYaaJafbUhDKp9glAAOpkZtbF
OTsHFocLeJsvaP599sqeUNkStZvTm3nJwxUKR1n0qymcsJRVtOCUcD6QtpGvJ31REXXuV1HIxIIp
+AF8Qkd9JnfWejSyZrSywvU4IoWi2NduAly+8IMcspg7KzAGf4su0xxMGuSHtdWxhlFwPl5O+UzY
pHeqrDaKmpgDKhTlc+SawUbSsUZa+rFuCGudWIy/YJHFkNSX4cxvudPogSVoIhcR7wahRvji4tJf
oMvItxSQ30t7pNauIbkx0UZMQyJo7ZccS1Fsbekf2iMXmInbYrdCMguav4JXtHgWlYHwuWFoQ28T
L9WZYw0fiOjoxWGCURk5vVwb0S4G4hZikjySCr11VWggc5vsgzcTyx+i6hIFLiCSziJt0+P8iJSj
APNzz/JzqdzUueeMWTKuXHy6w3ESt5XSEi/+sBszEXM1JSZcBY+rgn0Ne1KrSStHzg+NCg6M8xag
uhqPB8+h+oFVkUZQp/O7SoBgjRbLw/xntKh6mgbde3Kyd5FZFCEghZgB+jUGb4ldSX1KnLXzB99h
ieFmQqcs9lSLYTC6CQ9ezEESqPb4MkvkVQvwJnSBOFgUVLlVBR5fGzGgObQ08O3de+hfw7ddANU9
JX33NMn+K33842c2JhXtSS0elpcjeG/obA1bIbuMNkZeYDvauH+p6DGU2MF/R5p+lNioD5WLzxPv
TIqKR1OnHe0rqFnLX2GkAOU53ax2c4Izw/vMQvzeHfqU4hzx9lKiOR5ydzw1WStvYpXfuHnXdjHB
ZxVzCyf7sPBg7MPtqNpYJcZMTa7uYOclCiKbP4Em0BgDjf2AtKHhMl1Rtqs9/jKTK11P3FHYIWQ+
c4yJxAI+UHUPoXt4r+wsUtJoj16iE751LzHTubCmYoS3RHxbnr3HYO04LPeBRiGp9KLCImHXV1cS
8gGoaab34Vorr87qVoAWG2GNzYSQhxCyvcuAK0Ga7+YTgZR6wuIDXduQtl2SfeiDEBrmHIst6mOD
GzRxXKPT2CCt7pLs+CyPdCss6wJGDTARGgE9OyeLvbH2gSoJ9OOak4CNzQmWqBuOE0Xj64FON9xf
GjaS2xk8VzgegmLzXN/WQ5PWl37+6BekXnIlQgn4LbM6Ro+JxQtjHAFflPFpmP1dnnk3660vIZp6
8i/EjG0kx7UGQGs94ZexDwIQ3BQOKBaRI5AJDcdPlpdVQ6j7U1iI+zqGtQlCaU4ZirgdB5YMezQk
o66W3gQjXl3P+H2lE5Lm0NmoVcpjZ/GQTCq30h+IyLeX/Ot6+Wf7lFTG961CygSGShBwGhyUJZyo
7FpD026QHUr008i4PzWj0pfWzV7Sz1u1L1ZpLP3d0NskIYY2XdoR/qHzXmY57O/bxbbB2LK+UAxe
tZE1rqnr5pAKFZMJl9kHUsymVwPfjf63bhxmYwDy+2zdDl0saUqlzWfYTJ70zPvxX88BtDnUcjqX
jvNa1ijpNo1ctnwSH2lOtyHHsC8zRVM7JSa1MrgZ1qro3Cfw6X37wr09syXfLUPNo6v49ahSKCfA
Xpu6M/F26WY07gS6ZA6ig6XMFd/lRZGSRxJUiJYYHEO0GDDq44HGe6QzAFLo4Hc4A4LmhtLUtZGL
wEZhoYqVsHT2aSnP99mvhdY2DNRPaQr8EqQi5mtx4s8R376f52Z7/F6DvO6pBoIptBVCEzB+vgxk
Dw5mFnOlm57Vf/QMoyIGLMjwirzGlB7Pa9d64hT+fGYigae3dmfCiAs3rcgKGF1pQRyFe88bzGQ5
vQRdw6r59S6+AzvGqbn1Y6MycJkUwGyO3lTSv/4zhdQbsTRoSEmzMnxPP1ytD0rdDBivKqhosqU2
LUKW6ToB+A107QUbIK4I7Y2wPHkWcnQQuOQ3FFSShD0l043LaviCG+tZwaQnCWJcsTD3NOpnwehJ
BkvqP7VGa0+qglUPvnUY5tbPfkzxkGe0NVWjxexNK/bskQ6jG0IwviQZzsxnBx3GFmrlYtnqKO50
X+LBU8u/RGxpNz22LRSFuBHqPNNDwxGzFYF/+j3JXIsIAoK8KmTVEY9q99+4pVFPwgzFDK6HItYj
LIyCezqepgteEQDVXbM3QsQZQn/CDhE8OvW5yRKHlSxUlxd8qVPE+NUvp7tWIgLT8iGBw+ILcxDX
fTwGxoGVP7fN10nbtKmGURUqiPTnOYVxFln0SC2N4iS8vu0PE14Duq9WIA5+5jKllnqCA/DuIk7z
a22AsdBW5ptZIdBO6zNCO3VdC3pK0gN+9k56cZJnZRtjg7K8NszOzSug1r+VVZqgBoWe7YaM+Y8/
1wG1R+mBy09gL8mcgUnTTjK5ar4fn1BDUCg8abxAUQrnwnRnyuziB3cGwdbJO+f/7wEWChRQI/l7
6G0zjudIYRMMlzFp+cjQ1JiT9RfebaYKwa4NVqJC4xH1xwWAr3uo3Cupao9bfP058XZxRh7l+YS0
N5IHfdmvm/nuBQhuC9GCi47MwZMhf+BrDbdgMm6k598HUW3xBIzyA030BWUJXMH4XV3Mlh3Tw7fX
p8IqAwYxAVnDGGaARnJ6csDHDARfO3lQyYkclzT7ReWDlrKr1bib8WuuhJcq+amp4Mlbv/nhvDkN
R3CYXUwrvLCl5R4A0nO+fCM7KrGE/eok1uIq/xFuYHNzLXMS8rf97C7sO/gZ/hZDgGstsnzjDHcT
RudzUey9O3QCGKer/EO1T6KUPwiVh8usAT2Vl2pXJ4iqXacMTV4TL6Rr5tmLA4hO95HV+EoeQjjd
hQEECiofgkQG8V6LZqZilyV+qmtbjXKuPxoqWShjVHI/3XEOWvrniUeyD4iMS25e1m3cQNbWg/Gu
VludluIWvMkz+mPGjazOPgj/8XZ0CRHviXt8ujAhHlOC5zbaTGiRzzcEm1eMVzBcl4DIOfo0Jmye
QBO78+AluRRqv0k+1LDngqKjes29UCVx9hcFiKOuNm/KzdyqSxWeJQg05ttCDILZZ+ksYlkgtmU9
JAiw7PBvi86IMM6p0aOHWSGhf8QVsR6ngMY4NM3bSR4iBbB6CotZwYFH4px6xwQzgBS6dnLXFgjo
2OgIMrhgX6TbkcoQF2Q1FCMSy0P6wGLleTSL832HUel5hU3k0unFjrBhL8rfzOwsZVp0E6oQ0Vkl
tbiecJcBlZJao1D0sCwd/XOJ7pT7Pgh5XgTuJBBE4hlVtcxd6T+3owf8IejBu0iKUAxOAOSLO2ml
CgtKh6KL4qpjy7QurxouzwxTP8mn0p5st/8ME/FavUQd+ZJkOmWyRy7fjH3SLVck/gdvVzY3VVxt
0XZ5miexT/L5xn+owlq+wPS6RIS5Gkw4f0B28F1KXoDrkKfeVsWV+KDOv7jpRewtYEI56SAkRCBz
nmrott+BRkeLsYzMJyi5kH3n0Wsa+0nDhYbeOD/poBYhwqBPrODmS0LoY0aXf+5LsRf0oboTv+Qg
B2LI10L0C5IWfrdK5c6SerZCTK+a2Q+dXj2W4QRfK72W1jxzKDtsrcEyLHRegbg/nOKrO2ueX8a7
xb67tByaPO0cMjJSMqzOSDga7B4syG1vX+uN26r5M/ZSh6blKAp82JCP5+Zbt48ach+uWYb931D8
RQRQEuIyCHvXFaWX0avHiImwWoytHdDEaPo0Gd6rJZvj4P1xOt8fAZFd9y4C5F2t0kFfIhiRk0Au
TWNPY04TdOo88LHqgh1sNXgcn9PV0dek+k/6Jz8kRl2xg0ZAaRXAJOrU5MP6/iE69/LBT0JmKBfL
jMVomxR6K/laBR5Bm/Cm3D94h4ZCxYnuUnvlEXpfDrEwlwVOSBBBXPRiZkEFTgNq0ruZM52pL+z3
gFCFyGYPbWYbIEBrJ4WBJliPrigeWXwYa3ngUavk3lrn08Z0QAZDeDOZsySDH4qt8Z8hoNSJeTBi
2ZCVQUhn9Fgo4KldB2VhE2eI7cI1GwfejODTZw3DJcV/axyxGAktEnDSVJIqXDiJCrjskFS9cFmQ
DDbOyCtqwjAKBUxWMpQDWXrGitU5PqqjLtv1B8IgrAG0w+cJc9AFLrUEDmCCLo+b+e+fU4B01B7W
gLvL+9vq3HROdUOjYpLi/ue+G+mVuxMOPrwHmL9IMR9dvn3ilIn3PIEFtnLfjYiatgZWm5zGgiEH
pa4Lk0M2DjH2+Y7XL4FihxBsLHAePbenYnP0ehE95cdyJ2XqlWY/7AOjAQsa6xc0PEkub/3l7Z1K
x/Wy9zfYujJbregAK0pRmoPmLhr6q+06MKqaDRTx5Jm4C0EH5ZLONlu3euZg8EDaJriVjYJFxU76
PWV2TfL2fOR5paAHfpq0r2oN1hoGduWfhuHaWuDjZq3JPJgdnwrts+1mGSn+2456JQGmsQ2ls0kE
vqYM/tA9/5WXicootAAnEUc8nokvg7qS94ZTraEhEqGRWpcfRk8vKtAIa6b3+hjdk2oekluYshwQ
y5IvPonOaO6BBr6LVkXRWzQoKHgb7cjhNlLgy2aVr2TFAW35yqCcSLXapH1mfEiG9AkZ0eYWs5m8
Cd9UMr6JTjjqMNPArmy+rZDmsBt4+jTtxzc6cCzzacI9x4/uW/61b7zwMtHGLiwCHwvuUYgWrUrd
7KEBedaTtPpe8v8xLnQNXegJxKDcqSqOYS6X/eRFP7/SYy9Mb+wzMtuLBwPvQ47zrVD2EE0c03WI
iiVx/5TCDnqQ1HYqbjbYirBPhgQTYcHUlNKTR+/TgCBp8RszWkNhGI9WfFX9Ci7HhTM9t2a37C44
UEPGnCIvAGprCmjveqTCuJ2f0jEOicNxwSiIz09NPeaDpVokATbqD30sZOCT/GyRlnddDjKrca3W
HjmJMFnKYnVQdg5ZQcXXy8+DdhwutxC9E3E3YJ6YV9ZbdYWrcx+w0MtR+jDzHEy+ZLBHZxN6TMEP
G6n+o2JLALny9LRLk2JVq4w2Ln0ZEOkp5khnkWF0XBQieMJ/oMuM48AUpkpDp5jQiXXQ5dDwLeLr
9yzeAoct5LCQ+g+4banLeRiTzH7Y0ouxKBS68mljZRQTT0Ny17U25+//I4M5ktPJlT59BJrdiSeV
6+Sc15cWPY7e97vb2B3Ykt4FDiJ/dmhCQBMucKukDBLEdtXO55xP4ndHqNbpoDTfRrrSgqM+Jw4u
v8Al1C1/gLYvf3zsbpvy2a5PyUby7alTALDMRh//cFFcvmycBsyHEdhLAyhYCCHOMycBileNh5XR
HutAiGQ1XMz5Zs3vXWIjqTNPsbaViM8zsdY7D3R5+iVLgBMojRGuWtnB+iLSuS1ZBg2xWcZnxM0B
Mr2oeh+CSkwaJH3w56u5pUkDSF3a0xNFP/BZEgYU56jmccJfMob0gQ4ZfvM7l00e/cMr+Qsr4+bU
OwbOFnqX9xs7LRKhJ2200WbO89o2EjNO7P0+uDjluoIdfMflLrfsuYz8PWJ+zBt8v3XyrXSTGF2L
RUd494GFz5GvBhpC7hLiCW2MplX7uV4Blwcuc6kRXXo6QmaD+nldzbjHYrVJ9MwIuJtorGpRoQo9
Dw6gvuQRV8lBvaDcEZWWu4nQUz1Z5kM90KEsTS4VpoPO1n30hc6dlkUEcxXqvR5SXGqkqIeOnbiQ
2LNI8FvgV5HYqtOvDJY4NKAcq2Q4wqOedDrBs1W017oIlhnKszQLl9hCofV6FKHO3lx12yzm5blM
281nuNlqNC8hFW81wamh88Z/L0q3HmnqCChFxZEB7pTdX54WDLT94QFwWhZXa4HZUhHG55erO8Ng
4TyQBjYUL+pxxTqru3MXwEp0MeYXxWi0W/ugaH4WjMMLOKAmnpEYfGEZKwluyx8LEy55PdrPtcPJ
wrk2e0YNftG7WzbZb4O3ld9BgkaDYLN7uLoTfq2jnQuiCqJE/0PPMa6v29TEgn2IHb4lojRzg4pz
Og0hKdy4hwClq7PNSanog+ldyKVxIovmZefNPtsYluA/2nNToygwBzmkYID5fQVikcX4Tfu+NR79
iaRaZWUTECxL9v8LbjiUc1ucF9j67DRGZuh25xePVDGTqKE4+sRSlZICQeMdnqmhURCp1HZlZwZ0
rCU6PTzotAXAxw+rYETq22Ip5wWBVtCiN3s2p3t+V2K/4D9cga5fM8VMQOKSe0gtdAq5iD5YJaBI
IMDD0jVXTORvDedgSDUrlW/uvtljXNyDpHovdfqKL1rjCVyOIowcqXZ0SNiZAbjptoDNX//pna9p
Mi/Bx2L/EQyOj9/F5YgP/MD3z2jT8Y+a6OsJlH0gHzaJ3denmRxCTQl5l6RtsMjyBI7nA4jJq99w
FleBwwQHQ5WqGfc5eyM2kQHrzJd4I7eGfCM6QAVkpUTOY0BMi3WTzDEELfwTnt/gzoufQEmneY8E
ZulmBGSlc1Bi2uJVjcM9hLGReBUIXqZlNwCCnIXSkFzGYCik3Q3KcRrOZemcmMJwXU1TNysoA+nQ
2ejeiTjTFC6fREFfXqqaFhsRRg1fF8FnPurIczZ7z/BPu7VtVgEc0OnnKxrf0MqTFpVYd6DfBrC1
F7MyfnuTBa2vh/X+snOOUEL4pUswkaBxg9shIpJCyDldR9BL+xENf+PH6wBilSIyHSlgt1rIVBFv
cL54ux/XlbQOoOBHvmlGGq97vQBYO1/JCydPw2zyaz2d02C46fmxH3ZQh/he9FTxRKylGCXNFsDN
nAP5snfAOKGf+4+7LeArOohKUywq9mwwvmAA99LhM0YGY3cNJC7Ztodco6mKrJScolOzU0uqbRVf
nj7fLGEVOuxghskH3aDGEJw/k7+Y6HXYjW2l1hmNcWTr52+sZ5zmlcY4JgPNNw9h9IkBgkQPRB+U
jJsCQZCAEmlkIL3lrgxve1FRhs8Nmn/VbI6h9HrNCRkHAAwwsRO7DeuSLFrP4BYeta6ki8dJrr4r
Q7TJcg0dif6zDdITalr4a2sVh3juDQiO03wbf3KdLKMGwtmo0bVupC2yFhh85zg+BtCZk/wT1f3b
izoeNJXBIT2jOgASzQN/33giXPoyxyRgE3WsyQAdJ3ZTjj9LucY3ydy0mLQLqZULJ/rKf/NblST9
dXUR9xS1DAPGLip05XR7outXHWCCvcKGXaBZoxVR4kMZmwRkSon2MBrSD+5xheoqzYZLK+OpPkRz
p7CR/YUEJTcAiAHl8EoatuNJZjBYhsMrQ2sR98d/TR9Rm4BJez5LrEVB/DVn6Htm5C5wbdW9lMCf
Qu76jf/o7tkeJWgmr5GvSmsxeTjLqWP8486PtL06tRN7dYaxvPHFIyCTLS/bOAXJGJZQUrpQ6xUG
ENvYfLhTOfSTKbRdIkAoX+YCIXtqZatMAP+oYr8UU4whoYFbY2HS/k/a+UcnPFs20BHsbQ4qbCDh
25Pk0fXa2fJvsq9PGf9vTY9B4bfUHimWcf42/D+7oXdIxFmzQYhHI5Wbwl0SLe63r3f1H6bVqM74
OlWSFLkezsuxjRe4loWlp9cOB3Hn37HXsmaOivF6dCFX6xI+CvYzXR35Gz7IxqlpCNv7KCIEKSX0
LbIVDe/JYqsuCw39bcQ2XSrjcxJk+wybIuBiuzolgl0wcV9iUzGugswJxTzSMqOd17YMdO6OMBOH
PXS4tUJPl2wKIgZX6Sknbf551qqp6bfK8GSbvLJ4ETRGMrLHcewHscsqqTmZsgsgyWXeJ2pOs697
UL2vHFsnp+GElRLQD5R96MCJZmyl7Anxc2cMR6Xs/1a9WP9TRX5LCRQtoGbvTYCfBRLo7C+HccBy
LL588FhjEo3hN7iDHS9rumK01u1iqgQwD7SOSI2OSDqssiKi9ERP26Sq0dMNX4b77lKcWCGfFwiO
ieUaPS/MrBPUNYN9Gq/CJKaPPg0EjJoqVaCKv6+GmtFqS47e4utzJ3caAr4JBE6K506q5R8pCHwW
3rY4ozjnI2NcUcfZpNA+52M7/ckIoF5kcph6DWY5DXMCIilBbWYaUZlbghzx9McK7jJ0XpOsUdlR
fteRmPZYtdQa5henfxkfL5mZqgPqIfdwq00zN+HIvTQYWUCl6sjvh0RCipXDZ0XyTgidBGd2+fUC
u8O416WLcyEMT3t2Q6JY2hzDNtH6ZZW8yF7Z/tnFKNS3KZlpdcyBVuTLlzQ1r8sN4/0HPEQZE4/j
l4pspj23bxwlum2KRTL1IhC7ol0/v5YRR6M3jqPFoN1Q2NrKTUcdQT0+f9l6taCQ4aPLhGqPzhBx
CWoACdljT8qvUhZOe/1BIvppVvTVVt29jOxQL2QcMDKyUXmyNqrnICLXV/7YWZzKPrBpLuW6XEkS
KZ4N051Ll7QVGaS1sUJOhAG2tLt+O0FJR3XgroybIk6O9tJAWvBF2i8Ib2ZphIoYIMc/pbeNPJ6j
32aFkrZPussOd3crkSP0iQY6UpbLVlhJBgGFcIEzn1OKvZw64t5xMMjbuMe51A/oACw5iIhYKf1s
bv0xGlDnIPvK8gqJwTzHn6O3HUulFe/qdQpnEYtxNdEW4EiU6YhlM6JPA3cbaFd70sVN00tce5ZX
C9qPVnWVPrCKb6i0yKC7xdnrrokXrPBodGGEvlFfTpDuHYUVvel4WQG+Dbr8fq4I8wT7xBuC2WzW
B+5RkzUvSodwSzJFDz8Jqdbb/cddS9TFnHtrVtH4F717VO2d5b3sTom3yH345UVJhnlGZhSz/gVs
XMG+/SELxFnwj7uSVfU7HXsJn0T8Y7sPCX1uXJgOO/+yJdCm+iUDVDzh7YYXtIcZmGAIPcztSH+e
JPteDzRqMQgFrZqbPdvpqHVuEJ40Itq7OGhYCVrRjXRCA9iqk2Zg2Cc4J3SgsgQ5c3Th33udN3+U
073Cr0jcoHBIuTxRwCWYEXQQtyuCncVaNPUgr0imFyygT3OVL/TLGRNsepEQdE5X+6jXTEqNyx28
vZEO9tnv7N3LxOr+9bAFEMuH4U+3H/3ZCwstirR7zym94q4dcwaAMD4HGjmoc6/UfwKI1bVsLSdv
95CBkVO/sFEqjBvErWP55UfbnTt54tPm3cT7acuXvFUMuExNKXjjQpWPHX9J1uqj5zQpHaxpKkT5
pLT7T/J/bZjCGOy4L/pkGZys0tkluYypeG/XXTTOkB/EI0VkR09AZVvaYso6P7AtwnPnOnXIrFag
w0sxB9Xtk3LKqbbyIk3qThU49CtqCMe4EOKFlR+hdEYyKCFL0TqnyB/TN3HCP69G3xY3+3wT5foA
p2ojjH/Dfpf4UpRSGPBW+1Iobt9R0Q7+MjcHHnKOtGsjVLan1P58Mip2cep9Gn7j2dXZ1dcRACj7
7BjrjX/5nCTtBamMVflNYx7c1n404N/ikIrq/nlQMr7g0x5Y4sf+CtQV6eJrVsdOZsJFMZFu8Zru
kcC6WhU0kzeF9LfDZuMk/k62mqmByuu3AjPO5FpPKY0MweD0J4kC/dr8Mp1tySC0MTzHDjEmLgO8
BQqUHsFZEbN3T6Y4/pZJfD0D2MJ9oK7yjL/trfr2m4ioJGLsernGIs3vNWAYmtud6CBalOMM5leN
8eHAsF4a6vxxCocFxUnVF8QMsDvY1BueJWJYkp3pcu2p5vx8/WY3Za+vb4ROY/Wt//olnl1OMLZI
VxESFO5Ro045T+8htpBq/dfwv7YUXMHyKHNAsCU4+G7K6zVnRq13poEVHz2PsjW0TUKVGQz1ZVed
Kp0sz2Fgqmc3OO/wpogXN87yWF07lT15T04LZZbvqavVFoXvDkmMqc/SMfS7PMONE8BoucAwEypD
o0bg3kNJRsM0ygREMVen0JIPxq4EWjGXCGGIPsVxmuYn6k48XECpEgTTMTC6mpIh4QysK8+ysZSA
ewStJDm2f4jstxhGRphxNKb1DudJpFtTf37itRi7YxwcGV1b6ml7WLsQME0Q4klla5M8qf3uP9iH
/dzLz7Rcp4yDXQWFmSkIiw6fAt238+cSitielT1QXwk2XpIRHWMoDhQiM3ItDTLwUMTD2GkkvMcc
LIthRCyVe5vD3y5upRXxXNmv7WOKhKh8ybJ+EB2B9vgNhYOcLxM7XB9pAhyZGghLwQfdv+TXBhJL
uZTCx4UY2FWhfgEuH9IiFeGZGtdy6lEhE0d0kGbMi/vtUuf9BWL36QtGbsNX8stkgWpb05Bqvpyf
BC3wJsO/e2gTRQjDaVxmgMfxD6QIldxBqtfqk3se/RRTLiT3nsSRSyeK274aKouM/2pVZ0y+2ZdS
bFS2oKnGiWxs0CD0sqzxMVJlNbzL/39/d1WcNZ0ff1Hak+VCZvg6c5nbqRSlJgUyA6NZ3/G4GGni
EY6cpkfVMEqe2k7ZPZTHedk41mu3iV1IqjI6vb6V5N64V1l1Vf37HVPORA0sX/Bl+t22mmFD9zSS
vwSeqYBzIBD5smVyHxdBktDlGVaB9mE3pFwR1rO8ah8Ca1aDDmyrmv+gxFb4dEz8sfbzvv8t+Jrj
Q4xhOnHxlxfikAts5iQvWX0zgbVsOwebijaFsomcOjz2PUnJ5uwVr3Cx9NXtUgZk5dBz2iLNl2xr
E9GSGM+cv4s0DOmM+Mv6+9BJyuFHmHscUylpgHsz8VVrsz4PtMr9kSwp4gSdaApPp6GhBGaWWlPV
RTRTD1ZJqajZ8/JWQDagbWgan77B464YnrgdRqnmezv20FLiu9lp/lu8aADhe4ZorYICP2/lDddO
txSjC5jrezx3U2jIWqTZ3GyeaOrBKFbk2g513umm32kPCpxsd4twNMSezeniUSbVw94LOs8/8p0B
CnpkTRH0zvlPAQqCY6ZDtFNiYItjFv7UT27a2muRI13RSlQdizeedJ0WKc/tw1YOU09OF53Hwnik
CKBYITXsF+2fT+8aQ7rjQZg0qdJHjijUuMSjKnw/5w1Wi3aCW9OEZDSxry8q9zE3VjnUc29YuPf2
Tx6p/woA+sNcSfpOHYGzZrrc1TvYrmDZxrz0EivN0dScbnOtTwNsoqyU2gA9CJ86d65MOIT43Z7y
/5aE66PEekfJ3e7G5FYgRzZ5/oXDb2AknZfBDX+E5saYsedK+nET3C6tWbhuHmLg1VkZY5gH+sTy
CF4GtFyV0LmMFsMp+HnIWvbETbsj7+sFu9bYNQTkpXhnTeuzF5mfZjmSJ8XLdK6R0ztPEy2THwS2
VDNrFfu7X4IFQxMeFy6AxIyBe/+hdefIM0Jj2lT2Ej1eHFJF3BVWWwD0yNGbwSAi2qfc7W5/YoLk
cYYtUZdhpWg8eVu6l0ugYoodOTmmOpB4u/BzNzUpH87FVVRWFhQceTczP30z18fJSPe+UhdK9a9h
wA2sElSgjVzm5/kHblw7P1rr4Lln0M+J7V4qxqfZOwvtXoDNzoabvidXDblW852iVuaCF1vWYRKs
yR/BBkynHFdqymmj4IMzQtBIlDFmhn0zFphYam8yGxcNJzP+j4Wxh90xSRpCBl2SGtlUUcrTUwa4
Mf7R3fbN/IN31v/OTNiida4giVFmwSbkUcXFzhz811MDBaj6clYtBijrdg5Xpwig9sUedpuYo5O/
bAbOxWIQKEeaqZKzZpEUFdDtozZjP4SiPFSZbLu4YQNFkYzn8mHSdhJOKMUzKBKoRKKi6ilnNYtv
GdEIuTfmXVYxrLdT8IWQFRRbhPk/ucFqBhn5n9XUOw2yhJZs41nBfNTZLUvw6uEW/Bwgecx46fIG
Y5+wL42nDWM4mGbbuK0Qk+eLZoENmzrCAQjiUQlqVNrCugwskmlHKJKmxy7SH+OezaHAHbyuvfEW
3XGi8u+lU7TCVySOMD5ORXkwJ06/X2Nm1GoQBRS6KrvWrPVo8WmSjuBREXK7rmsLrNT/IiJaNJlZ
TNHLdGKR+3c8JOA+x9qg2iMiJBocUotrJRgNSoFWKRGPjWHZtAxO7wEGQE6llW8v4eZePhjFUzBe
lhDnVS8/sLsZHCaWCsVuxQP72IjSKq/701kZVnNRbq+wS+JyuFAj3NBiJw0PIhEBJuCNjuVFM7RS
M5MAt1yK/bWfFUy9FhpH/Ds2bgkr8GGYJkClskqyM/DC0uatJ4jP5LYbpPhZ6GCT3QxvEG6sTf4J
83D2ki7I0ozrN2Oh111LrUjONVGdz0cw1DTc2lvlGFq9AO5bGyIah9QllDS/aqk/ZVja25GXtn8U
88wiPXI9qzRQEydH8140HLR2WtTnw2PPx+yLpCAK400w2E+Wi+6toxYmv0YqBUA4mv9qaSZj0n9O
RgB93JuWlq8JQtgFhmTQ4NCd5VyLZGfOI+K9RSfT0A5IVH/v7M5bVVkHvhPP/8z77OcD0Qv5KGxj
tuFzpQrZ8hnt7yfudJ9XA144iQLro4F2mnsO79HpaBe43JkmRPqI0UwHHdSTJ243q+I3dB7+Cm+/
KD22ASSpf6xt0uRqPacM7DEKu7r02DckpjjtfBGorLpHoT+RszhUB/h8JkdzcXoQRHkw6OU2eULS
29CL/MQnKewA4TuB/Lv359neHB521SFlVPCwlwi3MOLNzqaY8eP+P7SWDXMPxQQdWgeUTkDEsc9b
pqwlgBVXg/4pfU6F5dzux3sj6AQ1J/SvS8XIAAKE+m0QPlCTVW6YTJ9AgsiJwF7AwgJqVPPdcEEx
hPP2humT/ksWbjN3fapyfEwIe+vUdODbPJ0cfLGo1wBhxB2FxwGtVQJyaZQlWzLeMYJwpMtndYIk
OZ3dLMDTg0V+X25hpXMSL85xOi/Yt+odrAbdcpT7dlj1e2eOFkpdp+LK4dCp+Ps09YYiv06D9y8t
K1zf5b1dp0TBmYPX604KT3R1Law7BalIMyajgOr4ZkpWkS8gnZx4QinhpjVfGzbhOde8wAMYYwKZ
nqKMvdj1KvsWBAHv8o0hjKhcvlrnY42HL3TsGRWQ79zbiDSYMYhHNf/9c2dj+3L88SxroV92di7s
By7lpdSwdfEXOep/nOLW3ODE7v4DQwaHAdDOQLtoFOzhK768QJrCXHpcqdlcxa9KuEVXg6MpG14n
yF0katQP+2dUk3xvzruvewa7CH3r95qgJWCUhIdAhFnyHlODKi2M6efwasBwxlFJzS0Mv+Hw26+r
agJLZ0fprmHWqvVDmzD2mZs+TXwMRehkWGTIP0Mx6GYPumBMvDml+PajIUJUHN6reCjy6wSKx6Xa
e4HNAqGF5fK1gZqef+8WHCAa2tiaoQVjo4pYpBdVnBNTZ/N5aObDqMSwg7mxC37yRCYxQC4K2MFK
cvXhj4jlDbDT+HK4humfgSXSgkYWzS+c2bTwnE95qMjxLNyRdqKAn00BCA0ap2a/YLQx7cSqm0Bz
VfOj0r2iApeaWicgsQuBZ98ZOzZIERpu78dGEUOgy44oRUd/+aFy4WmQ9c0vF2lFK+zbiJbNCTCs
pAkmfKCUW89YlzbIYWlJRwCmgUcuF0HcGZxbqHgKrNb8id3Y/nzbKIfpnUoNsTvPzgV11OfKC6W+
f/pcQd0JXd8pV4kae9+UO280/N5AxAc0YBawiRbFXlyiVUTz1wqGLWaNILzKv8MrP+sKdPI2S0R8
OIlV3z0t7D74v2tMgItOfJVBwXZ0v4AUgYKV4TumpzNq5z8DSE92frkJSijOhXxTdkTKTp1ZRKjA
gXV4Fva5B3N8wvbQBs5Vb0yH++J2ow9wZQ0fIyp1AWwSTZY27w2OXNWLtEH/cfM3qg4vqPUENNTB
6SOtmb6DtyUR8W4Ua+fzDG+Jv4cz1xK9HoeJDCMS3fzzRUHhld32At06WKXgMQn1unkOK3z0j/s/
qFwkW3a3OeJKBcFxDhmhPs5kG4uwRqOJIOhNLUTwC0TNtSfieO2nHAqRwIHYHDTeu9un50pF153O
Y6T6qcnF9W1LuXeH+BbK32j4q+CoACSSixH5qS0dmodQnmb5BmdzBff268az2QdR8Iy9Mqy7ZZLh
cHBMlgtmk+D0jaLkRzCy858YUytuG6JVw1NjFG4gSb5WS+Z4OVvi9ifcmoxkhb1/oK1RYqxQBej4
l12kwnJ/FHjUfEqYSu7QfM7F0Ud0DrFkdHLJA36A9oUXkrHYfRc7feqpyeleDen6V+lrhcdVfubK
q28cx3TZvC3jjw6u/VIriU7S4fr1eTeb4fnQHODTgc6ZrEy5WW3/YzYYd3VyXE2QFDFn216FkWhO
jnmuht1g4KJlKOMYgP2jC6cTDqI82TTKKVbPL9e6gMJICrgbNEu0pWPU/huCFgexpQKW1uqaiShJ
WtbtIRKOq2uMx04KxrMxF0R+Lj/8JrNZcc59H0/nK67Lv5rH3kTwsc/rMg1bsrwIcvmB4xQ6alyA
lku70RvrRVdBqeA1EQANseDP/qqwIcq8Mlo6UFKFe+FlchNzf3bFPP6VzZqaL24cuBP9+J46GRld
qqZLSa591EcmsLCdjiG5BO/Ru3q/5EnyyOdLrkyaPgAGr5btXjoRDvatOBGXtbQVyFDVsfCcEUq/
3IJlas2VQng+4EjENDUN9cBzxOeCq03KpbN58Y/zF6BQcaWaNkw2+YMSIxLpKm+1cu8FzKRYPgmJ
6v4K39g5K0kpT/pQMh7L8DCI53ux3j6GLNvcB8ntiYxsPXOG98iimt8X4ZXKxt//Yfx0wFDVW1+S
BEg0l9emNtXCz/KHwZRakDK7iqTjs2M/Mg9S0fv2hzLRsNo+6kQ9xUen6HGS6yarS+cGpSqv3DJQ
SvEfEg/L/z7PsU6Ot3Qth8zaf1by/f4lrnZ4emD9iWyLdDkw0D0XvIMdQMN/ngI4z5VswE/39Lvq
fr/2c3nWBkTkzI+18o79AumWzkQmKUprNhJNOoTDnnuYngyzu+5h/EqA9yDheUO31RE/Jff6ateU
4wnMr6GOKPfSh9jIQTWKLQ0Pow6duuCqZG923E/ujMNXMJOTHaeLasP183YM5YIEG8D1AttkvKIb
jOiTVMw5SwZj9oEy2wQpIRmg0mds1+YiHlwaTuLgia1YLaWMRlNQ7pK/9NzhojQcF6K9wv6uos+E
SLbfpst+CAVK7HLPz53oevvW9C6p8NS03RCi78ToqHUk8prWIYLBEQL2cJZpnRbDbhV64oDPb38S
TLLlEAW4TQz1ZTCdknlGJIqnCfCgfGIr4yU9KvZkM05aTwL+XBL8GoLHlcsB8BxMdJh9i/z2y6ut
0vFdIUI5Gb64C2ZJyi9Lzw8L5HPrsI0NdWPR8rlacVsCKxN6TMS2mxcLPuLwZ98bqyx5DnSCngiJ
nRdPy/gATCOTtLN+mfLtspbRKwpcWxAr7uivRmOj4oSmF3rVJnvl92DY/v/h0sNZ76s01rV8GR43
PEmR2XQEzp0gExKbG5/j6DGUgzOYjpJu6+9JqplGmdkkyOV7GX3yEiD7HFJfftEIB+2t2u1pMJZa
oTdyBxhgDRvzIjAoHwKbxe5ezmSeZMdNNM66lR5FrqZ3z4cI1Mzl6rv165ilimrGgYZmf4rWec/y
zSgMcXBsSHGWYvj/j0/WQHHcazJgJHADu03Ni/IRl9qF9xji//zRxH7v8B6b75qsCkVWGMXjDKLZ
tqRfKMixgEia5qcRtxr4M/EtZJEV6y2URxCAshTiINwXtxexlKFMXKUfk2967G7DaeuZYRD4jm2w
OCdszBJRC76tbC/GnC74EhLM2dwoyg4YNuIuDEPzlC2pN3AkNByKWzK1T7QgrCLoKplbhFqe9rji
TGll/RNetAg8hg0HYvqhwZNhGt9mhT0UDCMU96+uINg0tfW4ohzPbYr2QkooxZCIYMYXsbKYcKR6
iNlIUypfptOh3dhWr0ke5+kpSdDPrmyqbqVPC6pNpS94gI15DiEiJZ+3C43Nlm5T2XPwhu7aZ3Z2
/bfruF5OReicVfxbSDkbmxbf+g2qS2k2wWOUp97qct+UKTzWYo0tG6YSnC11zxwLdET72CGk32Du
rNk0s1BY/Xu7CEOZ+yAG5VDJGMceshVaQsxLI8fKuwiE90RkD/PzFHwKrno7z3MGFjDnZUhxbXvL
avWTA/tOtTRpgpz4TqJ5GtSG70S1467Sj/eEfoCYHfjtAZyxKeIzcheV1XJ9eTpIxc46quaaSTJQ
5HsxOyNehbKyPs7oUgd+zi22iUgdo2FQ/8Zjtepge37NdY75unoFUAP1VaAmY+H3wxl6sBeYlx5T
0kgU7jhyro08llHQEhfufMKsINqmozT69XOIITLUjKTI5JTBiKyb/Xh95+VzfKTIUvefIAzdJzaa
AnhTYhiM42r2KXozVw2gwrVz0rso2ZYQICCNlweFu9HnV/yHZVHQxoivLZkRi1IRGjy0z0vxmEuV
qzKAp+I8rYCWbQGGzU6BmDsGRSdqJb5KFvNCLOzMgN5Iboxf6q8OVVmqdJFQBgVRIviA+m9VL/MD
2ht8DXd3I15qbCbZx4YqbigLnoEvk/Ue8i5NmNYE6d7z128EZjhNcwyx/VQWIL4BIVT/5DuV2YFu
WZeImp+gon+EVwuuEi9D1CJnXWfYPlxjaMMhCfY1NYj84tlxXY/SUqMWhbAweuJY0rPjCDJVH+Q/
BUWOjarOAGBca8eEt7dSuqgEzU50OMCjloBWApb5RiSh5qEkJbafTfGLquWWUz2vKVDRTY6SuOzY
Sb5aGQesoNMOSI++h466kIOJqC7HIfrYPyyYoBmYoHdqmEqvz+mDxU1luey2K9IYjCJlrCsG1kaV
Q1TNfPhn9xOO3XMQYBx+fEDjmTYmln7GALR4nSNALI2Z2IXSwDl5AcF5YpUGUqH7OMBjCQFVpW+f
K9ZCZdOw8+wZJogSRAkEqloEt9/UyHYPSFiXvMnPGz7HXQvTAB1yueZ158TxCa+12+BV/N0g6z+t
VydwTZjVsLcfj3gb1+55sJwhqUQMiAUFIQFan7MW8PPwYhjbG3ssLRnU06buKuFMDZtL7jv/da9p
AQl4rB9mOHGHJ+rDx79gZVEs4cmwM8FajD+q0Z/+ESdmzGFSojTYRj8ST+yqiuTKlevWaS6coW4b
c0VFYdFtuYMM1PE3sVdnJp5rs8MAWgQVXe00wz24efCGM+gtlUFsDUH/xg64XUP3Vuf+oIk1WZmb
1qLdTEF4aPZtiYoarlukGdSXfAzevp2dP/P+T4j6+Fzapw18VFebb5tYOkyHRfOxlPKEZ6KdVJd3
IkB8lkuoozgstS9g0zqrXolhcVZIWRDRHff4cnvN7okDlwiyc4vEmFMOH4HFPaBwa1BeYc420XaP
Ph/V49xZ7Bxu4GMEmTXS+4Bpw1Ge5iJgS5/f2WoDF0jvipqg5x46h3ZFeqDud1LLb9E7JDB8nuxl
imprT79hqNDuJNw1Algggjc+EPnbGXANIROe/i0yX+voXehiXxefyDR6NQ+GkcOynYMUAhpw9fRM
U8XYkpS2Gfw/egu2cbJIWOPJtFaYxNiZgAZm/yxliXVSGcJIx6dMackuXblqsDLJG3OoJkSrKbSL
Wd+CocZyDqs8EHQF74Q7f4Gn2WfgMSORF5b5Bgq1Aw1Xk0oXVIC1wX7EOHmoy4nnfEMBLH9Tows9
r6mPRkyHF0vbv5pruOav4CAN1Ff6Y4pFJdaJJCdAN0Rq/dxr0CJkJZIWxgK1K7ocNMKb52svNgiy
OjejYYYfQGZs9ZRpQpksARvKc2qmyO/0K7mXSxmYq9RQgXz9QvmZ9IzpMg4tFKUqBR1wyd3STnR8
zXfNbeG5AyEGo5Rl+TFAk6qIeAG+DwGmD0rX1/eSkT3xpuZATx8baViAnj735yJToI/9UqnxM8wS
pWeaJRDLki+An1TKoF5ChTSsouE9waACrjnwDnXeqeZ9eXCsmfyLhfZXw/LcskJyJZe+5E1cwye8
MklsMuI6hwUKPGdC7UQjVr2vNGBve7z0ot4l1fBAoztB0vOu+12tFndZV7XnByavzlzxdPHE5in7
bYwlR64ptbMlfbKZITeJ4I41IXpSq3tj0DXRGXlOLqnVGblUVO7JxzrGElgvZ9Zsncg8k50/YzTB
J2fRLbO7XeBm9wmsy7sMqh49xcs+PvBVQTWQJNy2I2zCirs2PhpULWPTsUFyD896TfbI80O+t800
xmGBLkjUwv2LN3dNZyj3mTDzudITKtkYlrxVaTtF7pI469d1rkn0CXJU6HSHoiWh7rgc9wXeS8hy
KNSH7NRVhnYxFpbo2XEDo/NuKOHrjasvZtnZ08h+kOsoik0G7XgMmq1Ka0Mg5AQorWpzEPLtztpI
KBoGGfQPIDe+UFLphK8JNGNf87d6Nsdd2DNc6G8WlbDNGLckKZyjboE8AFTIl14gfiMF9Kj9tQfR
iUhO8QxjKPgT+NGlJyu4WqQeDRRnhv9Y17zgFcn66NpUE69wyONaDpf0bmF8EbuX6jySi6NHGd02
TytzECjsRQZTZM0l5sMrzeOpkP1SNeRLTPCWUgnZXl0ncnXeTc2cDlyVO6sTGvE3a+20qUohFcro
O9Vow2hMYCWPWmIBeeLu2oHAhnFg3EPHmvdKFZw8VesE0r1hTW8GyJrFnnEZSL3ycKj+ycYLw2I3
2opmUqJlhRNGTT8lT4vCVRYINg4OTNZv+/yqrcR4XLdxkYOwUZio5XuNAX81r9m/VplkIMxgiBH2
DnmIWuEAJz+7dJIWPo+OMDC8ZdOBsY++MTIzIFSN3GG/V9e6i4iNzjsVrzFz79G4/eJ89tBzGSW9
zRB2YANlFZsIRPdlKMJJ43kbNOuiRXKMYMmHXJxf/G1+wK6vY7ZKhgBewrrlQFkkKa4f3Kj7ZvIX
YW6t8Z3UXlZ3Ik+cPSPz+/GWJQq7DprxDXoVPCAOR+ZvtrtuqXbpJNXuy7WBGmLUjzLzosRplklr
Ie0lNWjDX6k4TIASws9ioIaydFAeL3xTSW45zcd/vKiyOaguehwAfWC8uP8NJop8iOupUyRH/i/2
aBFn9Xxe6GKP2tl876+i8HAgvRN1gI1J6YyC33b0x0ZherJ5j0VPy+znurm9pghH5ZDSnS2/A1SF
CdDAfqqoQpl3dcn565DR824zJizSCDSBqEEh98wmvfNByrjSW1sZ/NDKZs5KGm05JRGd097u8Xqe
/kPfM5Y+V4zCNMbw4UEYlFp2PdHGvYYuD9RCcNbwGzP+OcRh0uWN+sxNI7rqOgE42Pq4zKubt0zl
PBZsZCbHQhDBtKy9AVvRatVLtyHW7U5t8p7TDKolekM7bFWbrT8qL68h0/sNwOlN1uMNFAuxLJvZ
ij0RtZ1ZkM/yh/2I51GONToFEqSDlRuvo+/kfRkehc2NgQQ3Q9h+om9noLRk0rt3PuwjWHUnS4ro
GsgJ8aGjYahO33u9DXrKl4hFlcEhgmT0e8LY1OMWrEAfci7Y98e0m+QvCTkqYh0egsLjL2AwO7QN
OzrfAOreQ4dx3gT+x59K9L5xkXUF+VKI5fMaGif+OXgeiIj6hx84YaWgT+OYAD7J/sAzhE/JQgjJ
wXkIPs66M1ynQJR86icngDlSmqfIvHOi4pwtm3OFyAcl+vi/rE+LOLDwJVxLAVB8RCSRDtZgx8q0
v+XEw4gie/qt99jw5LB1EoK9MRImxAFW3RGPGmHcQIr45SHYoOgtiIhJowzL+S8Hf1sUFUnCllwW
upSW+M+2UUPEOHWQJfo0A6dhr/STh3UpdYg0HuK3IMf5kx7EStRXbwKdKaKf/bZy8P97ZWsMT7Rv
lzWOvLOAnhcbv1To4+UBOsSE013wWYGbGlRJ3Xy5xQWXaXwCViiG80uCZZoQNmmed8m+MCbHtddR
ab9ejmgfyU2R/a72CsjR2kLLRKjzcqff4Fv/DxJTiSlWK9X5SI9nMVH09uJT8PKqpD72dm28beQO
HAW9+oDsV2UlivDp11csBEGYOxRZn31edLFqb3oQtyRjrBxeviUStD+WXx9uE8VJT7Y2IBjkz83j
XDDlJX0uBY29tEcPyJNDtJGdHWv/iCot+s0G8sL1OSQHBCVB9V1hlwuONicdup6t644FqVeRTbuH
u7OADNITCb0YLmgHpkqLIoRFG3zbftkY26RKccpW3Eg/3MftCUvXh4kVTlOsXh0UhXgXouZKfQma
Y7WTiYEzhVjJNRHMjiJx6KSi2Lc7ofwRDghYp1CwAKwhgXiuV2+d/pMf2ZwNnHrdZgRol+F0pq4x
gNLN3FKLb5nWh/a7KoLwCj1M7WN6qLRX6t5AmyEebV/a44QJFW9UgpCdUbFADnMgRnTRmgMMaYBC
dyHQaP128uQfDnVCmwG+Kq3gCyaV7WdQ6irRXZ/zDJgXQWVSRzXCHJQTJ7FlBJM0RojC2svgsdr0
oYxeV9bUZvgVLLnQWcNN1KlHcRf/K6y9DVsmSC72xtZ+qgSC+pOTK2IHhb5gVk86ghvzXdnVqpdv
1kBsS1DCIJq3XpYfabiDNaPvjRkWv/roKjniqVzEk6dtoFV5GO8K/M8/SwHEuB7uutDH9+I7dMdx
HriagfmEMjl3up/WcdgmSaB+nBWq5EXdLvXnlIVhFu4yL1qJPohrXVA6V6mWkwFnB3hb+NRNMplp
3Z3lDB5AY/sEg7uit8vxeZt0kEMVaXdSbbzZaJCuN4rJ4ExOgLXYBghaINtZ+Ty5jT4dqpgqr1pu
tNVzC7Gyrvm3ckpFbIGCh9WK4CzFjjt0XooDl+do0aGhGmXW07Of/114EkeNLDxrBwuD6Ih/RiRd
R2WncR4D+Vak7u5Zv0bdIB8cNweMWUcoQy2LzlFO8in7Q1GfcuZ2V2Q3rbgG6H6HaltAYdCuP2J8
gBInFqvg7UOvpcRp9jbPSb8T5A4WwaaeZQTiFJjz6Ioe8H4Maw/qDbta2p/HiU9ovqInNinjz84D
b13yZ3DyO19l53a3Lh723IU35Qmq5LnMqYmiOH9ob8ZcvpfYGE3XSxBKhFONjXxFsVROg/XXCHl4
twuE2V587nbWoeOFy3QbVvYpZ66ZIXhD2YsTU3E1bfcOiIb5wrUqbWPv3zONC/7qtKHfuq1JYxnf
bvhOk483PaTZ5z+9RsypvKZdFMeg2eFRItV6iumTUZ3lptlGVFATdeEwDmhGKYTGZ6YjSjFj8hyJ
asS9a+tFUMvTzDCS//P/kMqNd7pN4zka7IvCAa1Va19/4Bo+Ti/DXp3ja0QI1DyzQwju6THTigCT
xyuoN858RsWwiz8inpxSBOQuSTV8GH3uVi5DzL8KZEAs2K/OmmrGw8o9PR+F3bGH42EuMl0jEB1p
vlUx7Pinqbdj3C59vcm/7B30pbwyvw7SKUPYDWSIkEeseKL1kyvZkTfngDPhu2pjWcVxPembdaK8
hA4edkIvpttVZf06rlt3+lIG4qig+3X4PtCZtESN1JK3GgI6wEpeK1E1BuchTwixVpH9QES6CrwB
UseR5y2Aqvx9dozNEe3ulcZfE0ImsKMf6VKLnhqmNpWorZNRAEK+UobVkhiqIsJMIPBUqXoiw46K
cjLKeKX76UC4n4S0WJXNn+eI01rGiV44VTFspdw50+CrXOC3Iqz86tmvg15GPcqszBKpu+OLJbC/
laeON2UTl2hvDX7uF29KGtvw/oSFzWXbH+k/aXJDpsMHJjtt2YB+QujmpoQEsPG1h+E7ecdf0RFu
Gel/hXq+2omxJF84hz71JjVLaTBPuX50AYRDG7LgZVIuFeyE89q2eH5zM8iKvY62koTxRGdwyHet
9IIa1VOmzjT5nrKluDSCCUgPpo2GbHsQrWHIIbqay1riAkwO5LcMlKntE5Rlcr2gVLxtPzkz69Cc
XDb++uulDN8HB14ewQr6rUiNoZEVvNj67exN/wwOHC/eCzzeuiEaf2O/splF2BfXe2xQqopk3mvn
T30wZh2+5X9pjmxFHvgm5vMR8uuioUklnN2kbCXWBtb37wbvsOtkeuN0AWU+2nW1yS1KHsyzlnU+
W0jTfaiWulL9f5Ltg4QdihHOKi22RDBR7siGe6VCghrds24tD249lXniVMSHQqRKU9ZzKEXrOeYl
gdNKD8CbM0CziITqIusZtATVPS9bYnJQieD83Jm7yniCZe6JKyavrlAic6SMM/HtCNSh1xxc0NmO
P9qxhVmSZ/LgqldmgIjQq/rxUTG0hNYyO50XgtQVTo+xu9toYPk2C5J0wmMcB+csMVwVthCw+Cmk
b5HQT76UQPRKLiQNvHzN/CuvM5akeO1D/FsfZ0vTw7iTyDRV9YLkKLBc6T9o91SsdBSm4MlUtVga
G7UFhYKHpvlvh/VhS4I0fB0UiXg0m5XS18sRTw1Ou1abkjN69CxyaOPTBNOnYZxmBMQx0SWeCFim
vnD+H23M/tqElJ5KvdNtH0++G+vwMs4mJtYnecvIyHOCHmeJHpaiy/ipRvHKKZg3nvQFekJbxuAX
Kxs2osQwrgBBYK/FM8yD/SuRiTyk2JBVgAqXGY+J+KviGUYbNVDOztfcNKCoKsOo5EK4EooNhKx1
VEmMrjCpEWECgsBCHb4YVpLHCibVqFTY3rd10/QIJdO06BVXTnQw45dRZJ59VpFDs0gBze+bfX91
HFzYNpe+0876CbqNNp2zg5JAH6zDoAY1guobi/RbXztNA8VPyWKwWQGy4TieejVo+9kkaaLxBHs5
1iFQ3xPyPt1mXTEMCCdDc8sK7ChwEWoGMgSMfWGGjHmNjxBMuvnWV+ghELPuyg3KqawRgKETttGP
c0CMvJtOwPGRoO004nhMK4AAfJrVrM3C04mhFejPoqkzRTnheS6vcSIQN12rVUX5SO6AD7p37Qdl
1M9nUjJjXcXW/7Hq/yCEeQONnt02S5TV6Q5T4ciUTKmVG9R+jss9b/Yy4VMusUpxNrrjdrqtpcxp
7Cu9El80FgQs8N/lDmAPwo/buY4DS5uBuM0i37OR35E2YkvaMWXwPHNqkIb7iXq6rTf1YYzuhTs1
42rx6/t+3d8XzTEUJf24kpqFqNPebpbF8vJp3KpI6Lu8Bvb15d/NAeJC6TODzGWRsUAwfYc0aLNX
Ov3FrNj9PeTEBQaGbLwncwxikFzMNo+mufyF1+bkEgS33AkOyPsJb3zAR04JsFNyC6DrTuPsVZqH
t3HPB3UV1n5Zu3IttA6Qx9dp9Gxpl1txXcfkapvvYOZ/vYPDvW6uC2B3UJ2NfbH53dsZqNlAG/aK
ff880WHZKuHqTyWjXSIc/vWPEGnFgvYBlq95/p8oMIh+lZOnRFSykhxQjxZD9Bpb2IEA4cllbgxY
PgESgr+XCIOVulzOADLGm2EJZLjqgqZefWvLboPVO/Kho8usyS8ym7GohFOZaDHuZwSL5s+Eukb5
Bj9kk7pOxQ3uRUYKMTdC37v5z6oFYUQeq5HjSigRwq0EmOH7sK4QMYPLdt7x7Ry5Dsi7jAS5bsvg
yUrM4Yk3I3naSJJQRrYF4EoGFGllyBtbWkXJ7wzhjmPtedmBsgKN1SqeBPEFt+q3Dg6Rqcc0MdW0
rYoPgF5aumat8rzTnvmj/xj9K3mDVlO/o+gzcLkrnOOpTwnPpe02hs+E6EOgP3dLm5DruFz+m7dy
uovw6rIBABNaFKD555YeQuUrJzvwmDeP3T7PPvnD69cl8jiGOq7ddNreC2a4CsXeDp0rnCPqCNyg
av1fQepuEdmb+p1VzGeEKE5zMAuqhJbDR8a8XTePY2zKnriuxnyOgEcgwQ2LIpOzzfZp3WbO2k/J
rijlQ3qWPnQzCrTXVq4EIrKSR5i/jWjHNkBPkZ2XnOaTdyRuNIcRVvsWdTOZYvSL/YOY1SEO8YpL
VbH++InRbAaYfUZwnTsUrFJTlBggKxr+JoCTiK/aqUjlMop3Q7Rhm0bBA5snCnwayGNqm2sLi2Jq
YXnfgmYC18uRt4hXj17S2rOYa8y/i0W5MAngC1Smfu8dbOXHiIKA8D3RN5xcl6po83Ge2qN+wcBX
kjzMhOl7qBii4SH8lchbRPTFnQBpJNPN58T812d6LuCYZMtVS7LS/eznjz/qCwvgTbve1C7xu47c
gNfrI3pmgGx6cuv9SjeGwIJiNk6W9e8YXTaX3nkVXJ6m/gFkh7NU/hjrBR+s1I2SFmOZvipCCTYo
/SfbkOMjxlgHuIXMAHevMRspc20jTuXqbVGWUPUCoIJfD1SVbHQPNI8musocUyW/+DfEYYgwGDuw
IJlspjPV9pPUnGqB820jfbH/ahy7cLyZ8NRm8Putym7eH8w6gy8vCgAIyuhNAo1M8/sysMLflBCx
4hxBcOx6yF0zf9V+vPHdtW3Rq2OhtFAR85cpt6aPKBBicGkjjOkiUTW7JVH27ceX44FigcyqdcDH
BUysLETW91xgRpq0VezcxhftV5hcmgxsAzy8L7sabAvJDJZkNjQUIH+up1sYmnN5/MHO39YTgw8S
WjJOAc80htTJ8zn2smP9jwi8OYrgHGOlJNtZSUr3V7/0pzm2V4cbsbkLcqJ2elbmT6aXBxzpgSUf
rm6RxNr6oEmP1ePKe7LKban00cOEadgbZg5a+XIuIcdF5pH0OMxI465ynAc+daDCcMBci38wbNFC
ZIQ/7Bo5ZDMXgeMnjzuPL1GEZZUODTPpBOlJg1Kzc0XKOavpKTSqM7Zljb1BeGwMGlPkGbHVg2ZD
/CzoBfT15/p/L4fuppHGWsWNwJyb66VjPnOWhMUjN3QiMNhM8XPCahowohimIuSXMA2UdpHvkgv9
njHUJCJFXpHUlE9PI5013eFboaMLtJPc0YMQW+7Wgg0e4/F2CvBbBwBS3sPQSEivkPTteLMemNJu
VfVSS36JJ01QkHAxgfIJLXk8IzBS/NLOuNiw4aVvSdcqTnoQxekxyKGhiQxxdDSGvTHSMbAcyP48
gMD8GjiUQaWR3jYk6/Snr0hV43PtDnqmmJJjsF+oLwrDhOoQmijOic2lc3lqPomS3lWNdJ5ypNY5
PlMaeH3bxGxxdO6lVOJwlTRkwDd5/KYU8NTlJwzSiJOzrKkNYFm3kNoQWWitwSeFmBOjlzebAdfX
+6rLVzNtTe2xpajvEpXtEorsHC0TenEwa/sa1xSPbNlbAkvvZnz1HXu6RN6c4r82SkoQymKZeJ7b
61aHtdQ697W4lE7BWfIFcV5cpIdfFMIS/yMPJMKLtaxuTPqXUo0N0vraDMwZXFQDmy0qO+Cy7h0P
iUzeh3hYsZWhW8Wx7QJXA0tdfeKnbcPJBZrQfYXvMPyeE2R1iJckRF0R/TSRs6ueBY9Z06AV2CXk
DGR7XeExYCpmHaBMn++TJMxkMy0H8XnaG5HOZPtmATQLkuucqmTuZeThDLwzsFo7jkY+RiJb96JS
ZA+1fwsLJP3jZrTxnVjWyBFgSnJMEECH3SsmfV9XjJCDqhUIauCu0R8Akil147rt+cicCf7areqy
oAHuHjExamG32KY372iazbX2ERj+5Z2BF0c4WoO+hA16Z4hN6DokKZqilLhGbPaah/Gl1LN/WMe2
2TpYA9JfAwxuwwOglFWnFG+orAL8xCk0hrRDm1IwN2rDY5LgfMrqQnED10osu/lQgr3ZpF9GxH1F
pY9vygj6YfDgs8AWENV82z6pFfLYiBLJEP+r14hz7TJDtRHWVYTZCKzNVJhEv44joGwQvKpIEmSS
kME6AOxw8osnf/NjP9fiEuMReQoQs8k05bf5rUNLuj1EtrA4eScTEDXeyYV+rrfbAjPsBUaGD8O0
5aWterxFEgeu0Y1VACbxRWh5LYFiBxY+9z2kvslQEu1fTRyL8RhZSvbf5NUvxuvLjDTKSnCQu2SG
agGpQEeM6+jQUcg3ukwJ3lbkyC8+d8vonuzBznqcqqLK2mqnzils2bfhwsBAErkCblFg9RhUpFz1
G0VfH3WNt+fPteUfIxR3NYuj5AID6+tf9De10eYABuFRAGL03GXivb39DS91HgvRz9SDcWkFjD3X
c1Kca1pG2Z+0IGYLBlVRgKzphtGXQnyGrwyw+TUtENU1axCuvcUZqtHJ6gJOX4huaJcb1tPquknx
6lLselj0eWoL/9629UHf/a4mkflGgOg1hmMw9h6P+XUiM25cnelHmQ0wtS2hxip66W+YVeJWRbQ0
nnzUH2FUA8nRBeFx3mXXjPWjLnYciXEPWa5H7CQlvgPOnxi07Nnljo4MAnqLAYv6Z8LpdT2e0pYw
ZVANnmEjNmiTPX8cB0ltWTeZTfw4DvOkVn3z/ekKPBFdFK4QFuLlwDVmXupSEI9aZ7q+TqHcFK09
Ozlw3YNcCS+6Od6P5BpNwRAM680qy4bAeyH4CuWVQgwNCS0sfNkryPoAdTcQmfhuhQM2iZuTqLKt
f1ycv5/tsuikZDayofL+y3JOV0gDAyvkITPLmSyS0XApfafNbxZebQMrLJyaNnOA5KqlPwTUqH2h
VciPxT8EpDFpXSBOuatsCvdAWrvaNxmV4QvOsRgA6HhJKdfXM1Q4N8bdoxRT3yHbFY9eYitfI5jL
xjkVVu6XAlWEzbzHcIkHSZmE1D9fp3TWuBmwTmWKHmfN8qOywqv4L/G2aOsuCHrRNUuGCwjw2bdY
+7HQkVZLaOYCbUj4FSQ/QKvEbVqORcRL7kWlj46d5TGWiiUyACRqgYSn68HZRUeGLqalCXBPfnWL
ygfA8sH01sO4hPzP34OfewEJ+Zmru8KHHJ2VhAeLVgtGpr4BiTCqHUzVDVYsfinwaOzufu5dWC66
g3+1W43f2GT4NHFk4s2XCXZfhPFfBBKP2u2FtLuQDMm+6ZRAO1356PYHBqxBbauAvR8vgphn7tmU
Q8TlBB6YLZsjkLG7oSma14mPjwPi4rOvMuUjlejKq2qC0bJ1ZRz8vgIQSL+TCzWjQvI0Gx2bDmLE
VkMctJwkZe9BB10W6jbwCcTS3zP3nUNEFfjP34gYuqb7nmUKjhdR2E3NC7f0JwMMkIbdmKA4SABE
a8aZ4PptH4cmBPE6jzxPQ5JUkh6uPjCvhZZR7Fh81ImOyeHUe4yFrReqBozw42DGEu1AjRaDPaIk
Kt7DxmLwhaRPSTHZfLxr8FTTE+L6G7628XtaBQe/0TGve6mVJJ5c3ND+G2ys2y0IkH2uH40f6kH5
BBsaHtbfclGSLvA6Xcr+ZlguVvzhXa/tXXo9WR5nGdY1+jfaKddULMIQ7Cf2hGxj+5AUUDptyw05
dkE7vwvaNUi5QU0SrOBzSTFewTRx0UqOqzt/wCQTAQNpSgUJDp85rgs6X8Ne+fRbeAZ8R7y5i7EE
8GZu6GYlMHAAf1y6veeqglmYoSBhL14+5djpfmx1WVHbnbGTegMYp6V1syLX2sCGu0CXJGMBNEHF
Rsxqim9F6DPXCPaj16q0SiFZ/gZ2vu2GR4ZxfKC85rv0EK1Cr5mMQqc13OoxkdR0q1JC+My/jFMx
0zbGRIG07Uz153RKr5v6CATQ4+1+TvK9UgSXao2xbvEPFU0ZLossayQ5RQoOa5R/Gq6pRq2BFlKg
JQPby/qXt59dEBE/0AhQA5mYdIAetUVLev7hNB8nK7vdMvAXdzfwM1aIqrncx6YyioWbNbe9wyF8
Q6uvGZn4nKgzjlDClIOhqi7ywGUaDT/05mV3RypOmrvg5KMvwJ+Bo2A2mbjGe5jn3jXh6Bzrnuc/
35o1ztKAXpB8+pL8lnsyF4H24kn7voP2NW+H18Mv2/kk9MvwaWM5WR/eRH32A8f8asPIbpwEi7aS
ZH86sob3Fn0a1ERGu4KxHNXBunphdr2LtARcHKqpIOvAJURHRDkHwOLkfVPBIe+MreVFlLRUvgHu
FeKoJSltYjql4Qe53mv+aMGzkl5Le6DvX3E68I7jU+uR50iKfV718VIThp9zBCMZXfLdoAefZu8X
hC079IP6u3S4gF1nOoaWtiCeWe6JALfJToDgMtm/JfVSww3/x1jqr7N/4l4y02T64d8KtcuNzRI8
kwHf7WQvTToiZn6kcDXb/6Cfwulp8wVYus6rO0MZj1YUB5MkNo38AO4iAclEWuRjZW+yKLJA9zal
fTkCE4nphcxZr7D0kr6FROxmizfhDzRb4mAenBGMUXMx2RJIfVgimdOaEw5JJxNgzxfSwhM4z3Au
hl5Wqaxwagn7OsIrFmtO41p00Y0/TUazn+sNI6Z93ocz2oNOmCEKSQEHY8IMmY75+lZPGZX86yGP
gkgZTAteIPWVONLBXbC4QbgQKIGzS2WYSl232JibC40p6mRygW1//NWBsSBmo0LIs3nl6PnP9A89
ekSaubzS9wclHb8QQ9/s5iPfj5vdU/h56KiheAWcbxr9KJ5Xt7GWsoBRv2fhLmAED0ZGZYuhvtGt
7Aw5FBN/BGAzBxmn9EKnG5WGuy8BNRGWtsLTr8H8Q0jHxNrMd5iHAchg5k+eX/hBp+CdyLyjZ96Y
ZsrcAylVP0ldDnAtJiSUGo52PD/16FwdiGs0FnJigqTJtE58zr3KbaQk/GtsM9ZYn/h2gvxrVab9
FvW1Rnlx3YhOJuhjWFZR3lOIqCTJvTmYKblPU0tgIYQsSgSvBvB44ynBo33aHwjldnDSoWKqYzjY
moFfX7gTR2jO8hoSDBLt+sCwcuKf9PpsNg5/smnpU8CdjpZe0Ok9SW/I+UspuqNHxpMGsiRSxXoK
rlrTfG1uwfPc0OwLzgDulyquc/ncNN349Me8tvhoanYG0wnoPOgiXrMwjS0js+L6IpesHOIMFUKM
aCy5ZhcWI63JD4cXPINDhZcW6h7QFuOsfhhK1iBVNfIYnmGTnyYZ2/EgC/KNv+67MLq8ExlujcA9
D+dUQFYltL0t8VO52V0dSPFwOvzaABnIsFlWrUtUEr0pnlrvbCfpIBTU5ONhRt4I2jQLYfnkZJIL
frm8LgqsOp9aBS0qI73Iz+ChbVpN4GjSs6AmNQh9gAKQOKncKJaL+qqjYsj2/yXhjKrruiN6iHrG
s2mXsXZAy6pUD/SsW9QmzL53MVMCEr5DtDcvbIG2V3AX2pVzI2QbuxVO2Vszh7dF2YMnt4tOIfMq
9hiVc/Jx/qSu2nhv7pb3NAg/lMPFDkQrUqbNwY6Z6dttv5bdpcbfvrRKmFsUaKHG0khswubp+IVn
q2LGXB84ucV+Xf9atiyDAhxFu4c6B0HU7fymX35Vh0jjF2dSwNvrk2OrEb/6InNk0J0iCyV1aHCo
kCfA8vwTRRyrlX7QVvKWQDH0LyidvBzt/zLpSOHXL6Uwpa9HR7lb8+N4iTGVD0I9L81RLK9tYSkx
Rrdv/jFqLq8v02Sv7sLK54/52R5cNzaG9/MJT0aPyh/xc08FIyIaoOo5SMv9uxh3BsCS7cD1bwj7
E98gYhOWUbLaSgLwsVGk05KESk5qSlq900RaXTRdSmnyJ/2+vS0QEVkcs3boP3KGrhg/BbfpoJVx
hDfeUuVnLAssPpobd4+I7CCC1K06VLOSnxmEtiib6Mz3VdHFaX6tj23eboetB3wVCj1lT2Vqt0/e
z/+rE/SHCPWob4ne/X7BQ1+41XYC4/nCIrJYjLooYvwKrNuhy4VheGATQq1SqjV/6WetsqaRMyFS
4MFpMLVe8AgaBVo1F0ywXBf4hiGZ3Z47ozAj8LVMiVZpPBOO0mRI17wUt75LCbZ/kWzSXZU9iG6r
OgEOz+x1gR8pmtBfQRdAeKfPssrR6hEae57RO+13LFIbD6VPfWFUque0cIhbihnuLDboZWLrnMok
7bPm5t5wB8RPQv93CcFwB1yFmjvwySRqBKzun9GVDnG56uGJdFJ3WJT9Ci655X4xkH1dntNsxLcz
5eIvogy0Nws6da4/47JdDJ06kegwvFfTlcHUtbBwsOGe0ewQoTo+GPAgjT1oHATUBmSEBQMODc5c
amQyyDn+2orac4SXmONKmSN3PmWXUQzcbqT+zfCDWbSjXevW2sgcjR+7SMY2AjFjgf1JKuXIu+hh
sunjM/thuO9gbr+Zsxle8qclHEhzMyrSeacbhfdQTybY+U6cZTkZRIg8819YVA+4H2KSC+f5K1VP
KTaTfobyRDSktrAksS4MUQTGpDJMNznGiKWrtdnVwKf6eRU1DX0Hb8xKOZcToxQr0HVxgC9J6B7C
W0UpmodOtoKXvFLEgIscfFVNmBhv5ltmSVgpXlEMRhGYhgbYTAxMitxm+h5wS8f5aob/O4lXsHHq
r7p47Hkz032F0CTRx+UYJDu92JYEqeu9FYqLa6my3CP91xtAf7JmgsnSTciJHojqGrFxffkitNKC
AUlYWhSw5cwLYO3rI4J1j2uMv9kcqKev3lq1oJlwVtRUU+orf96DXQxHQn15lvoUxr3JaVJGc4zf
k7yLpAXDBk9/twO/j4bnUv8tTKYrKtpgO53YQ2dXbwOuZwBjXtl3J+MpI8IkJN5PGYttFbd5PXMn
SDrKJ3BkMvdRVIS4ZHQNypKIoxdfIiHCptN5VAOe7MWhpHdE3dquJeDUb4EIZ/y+9uADjEM3+FgH
zC4uZonuK8ygVGRtnG3c3sIfBbwp/82UiSi9CHRmmK9r/Nsv0Zp3UAvaXbl7Tw+WzYtxH4MO8WNa
C63y+FrvOUeIndTi8rmYVIklv8dP1slNKpf1D4d45OqYY8nOTZAf0iyZcLwYJjM4d6Aiv8RhRtJp
RMd7SAPvq/ZzZpKt469ycLcXKdv13KX2kPMbeXi1vPJP8v1zrlY48ZE3mHA/sBkGPFhtFHXI+ssv
/VZkfj7dJWm9dl0oHnHrXXaotfE1NuNRBUXzp+NDmyBCuhuYQGYKu5aRojwezE16SjsoQyB4s/pn
44x0NQ9S0Zb/woTGhrB1LE9uEbHjHTvzFM4+0QH1BlLrXFMTZBrNV2+JGQBa6pxJoLsN2pnkDLWF
+4QNjAikRmf/yAcpDLldFIjiAs5TkWEXecSNqdF9xhTN4XzPLWJzQUl4d68gzWVXqqqawwYM+YP/
WKtMUjDrcigdyGEIDWJnVog9kUQjT6ThW5jGqbglGM+Fn0nFENu9dKzMNu7EcoJXuLb1OEZHWXN3
mz9nrfSv5N/iU0DxF0Alw9Kjy9Hxdse/B0j+urLwSWf6O9Tf43kULTdx0r7T2bRdYh+6aryR4ar0
b4M4ex4Nq0jfFVkksDgpYdjinhjLLXeqbVFiDpMcEa4zR8V+gej4fTrZIpz9y+mHDsd6bJj61gvq
xJZwT5/b5NMy7g2n6VYWpdKyxZncv1LdUoX1yIyMdwkXhS+s/NKKBuXbeQHlWDCVziCSS2JcvUvn
0t5NxTt13ukn0btMcSUxk0OnQzLOzVCwO93F9f9txTvwashmYpZeA3atYRUNncDFYVaxYwJbtvP4
OikTisMWIf3nyECcNd21qDlX1VBSINquvo7mPskO5Sdt6VDBziuFERw54Anu/fU7ceaPG4kx4KUl
yk+BoFn4xos2DTXOynZpt4uVmGKaw2FACF7hNUQjCFqdN0JrWu5um1u+vvB3yHVhtKXcgVc+xBpI
TNY/pWG4eXWSp4aod0KQ/+RDUP+rCuAceSAAWQ2KyZStleeyux1w+TXDaQ3kbxSLpPOK17lCr+/F
o/o7ccW/NpeO1q/pFzt6mdzJ1g53qxVBEl8cz6lAulOZ8dnXKWjOPNnGBgctDTLZY0mxO9cpg1sF
CrmRQJgvn8Bn9LQ3qyWa9kDHR+8jdlu/906bxMDu5We/FchWYVDU8U40gifSiROIXCJ4i8VHo3vf
DYkkZraPJRlZsz2a5zJeXxXgaDLdbUncfM/PnMTBsWLO2MFDElhP5eNfq4NT/irc3fnfp0IWPypn
mXcHATq4WexDSYvPWYT6yG0CfACY7h8P1ygJGiZnhbskJOygXgSz1T76isLcPfnEfHW+xD/UySrt
TXTT7BqAvf32b+YqmzbnKVdW88PNn5X5BZB2t4VJFBDGJQuLEUDp8LsJbgiZPBXxdcrwCeCKhZsf
OHRE8CbDd1UoQz6uS0VeHc+KIWrxOA20gwiBnnngblq9y1niUgFsKr6NUp90XHWgPqtyp2nfPLXR
WV31hNXQ+Q9/QLlIgQdLBWNci3dtNyGylO89JSxAKB1wSMW30v6hg9dVcY++zwEPTGS8vMoQQehb
hikcmN8+YdiuI/nyCJ11SvnJje2JH9uGNHBjynL9z8jr4vhSXRRLqRt/saJ7NwfTySIxrpsbYFYn
WCyU4ajy6xG7H23peP5qgMmjib60q9CAkmy6V31eY3k8R3VscngbiN1kU5RhCN57UPmeN6jWdVru
tJHCK4pHHHjYr+H85JTDWeBm22Y6TqrVFxwLMsDOedZHp7/soCP9VXivDndl3m84gW4pbdTeDxpA
DPVfJsJXztSLJbVoZxpSrWr2GStEjNn/meOEQdqc7nNT7SO7EvIFFfC6P5IdOJoyix0XynqdIRLK
DanIZ9qiasSKFjo8Rb8C4G0uwnrsSvHjSyMutun26qG63MJO+2xFh2Ei2UkwbwrUEufWgtoHb0go
KQEyafmmPcfzvdwUMvfYGb/0tMTxc/Z6BIocEXtHg55ZYkWGEg9TQvFeTcCiaoZ5rCmfR6JpOt5E
bK1z7HZf3Z8n3ylYNs0qDqDKQ6oq+D85bsvKppHdzsmeJiwEEe66EP3GkxIDUSzKTg3d+nf+ZucA
HekImA54E4xox7vDTXO6un6WbCdaJzqOUI4Wf9Z1qxjzatRAcfx09a8Drh48uyfqkH1eFtY/O/GF
UcsnPrUafDXxQ6zQwsraM42Wt0v7z9l5SMvW5/BzUSgvGP8+pJ7f0cp1W6CefY4O0V9kJif+VrD6
RtqHssK9unJ8NPeOUfg/NeIH3z0QH8Ucvs8H3JN6bOEDPRoLTz5CAIdagLHig6WoXqTCOM7eCHVM
E0SySNmMw4NSFUOPW3atCgbdEbpg0gvKERUoCLurUmaO+5jelDz7fM1ifntVMgnvw22rIYWwVYBp
5YaadvVkl0kFVTvSJGPHDU42BrIZLSjPUIMqGGM8lZtlutrPP7K8UbKZqbdG1BRZT0xU7B8ygLdE
M3eeGPeZj7Mgpid5eOg1VMI893RJnQYx7WpTnNh6Xg9aTtQtnVB80eC6+sk3ysj9FIgIZAYr6GRJ
7FIJxyOf9OmiQHVnHfV1HHbteoRqZ60VWWRJnbiNpTbDylskCe8ylRUDGgrRSC9r6OvkzN70/UDw
7fqIlM6/csO/gDiwb4vA5VJ+MOhT8M7SD/jKH24PoYlBlS6dCMA2geZ3pbDgTLQfPd4UfpXk/aag
pVuHwchqyKftCG6fI/1MJ+EiZ24B0vTXkSXqRJfeaEm82eX1wTV4rMiSvMMp1RoWe1OhdQfYbM+L
YAKw8a7Z0y8ztJspweujNoquAn2ujaNPiB3xFPd6ONRb/nteqLEeUm9pwz8KseTA58oKvuYXoZ+t
7/SweI/f+/+2SxdTiw38oqTWbxUEmiyKfg3lnzBfe8Sv4D1TeRQJE4s1L0r4Mu7F6pcfozw0SAnX
/2zpd/SznKOtyjqlAPcl25MgEz/xQOD/sFmUNigL/DpuqyXtci5HWyEvdj4v+zTtiHnWIr63Upa6
aRQ3GAYXMKu7AY4sDG+WmW6yqzAs69TpvwSGz1Q7KbN574p/1xWccNilRHljijYknr+7UhrKM9C0
kgtCe9mYLQBxGyryNjjF58TD7fBf3yDePl8CYE/c1sTdSd+1WbZqWkAngXDhfmudk42yTqF9KWsH
xOwGyGTJ8YumspuAwXz67Izplm92xNSh/YqjjuXaN73LKB8iEyIb7Z+8dkJfjcs/M0vb3wtstnhl
mcJhQ4/kviYc95vJh5EalVXce9wtBK9dXvehf07voZMho318DLJ1pdySCpldzDc4n10sEr/WOhTu
gNd/GceZasD/0Hz0g4nkzrSoiHJcEhvLndKg/JRFBETIG9FK9KNK35qgHwL4I8uPPclLJ3yNUhs6
OMJGjYo+wsiDC0pK/fWCDxRdqc0/PHAWLLxu0yWi/AITY4P4Gr4pNsU3l6zNjzlCpOjJVGAkx0mt
i4a2tZQaAdRdG6EYIVSRSYR713xIEP0V5M/tu0n6GPF4jVwGFZqeXywdCP5KwgFRtzBJMPnLEX/x
KgfO2idLhmHIVC6LOILfyiauPHYi1VHe+DKD5QrsZC6AQJPMkU1jLa+e/2L+EYhxJQvH3fBERjuh
gPI/hjL1I5dTW2F1uA/o/lfAB9cFYIr7mgOXXt2wD2XqcamqGnMoHZ2yKO9z9iUXvhDVGJ06+pdI
x9rArCnByuPGOmdtXOSYVGFRh2mTT3Cwk9ANG4YVTwg/qDbPsPUNxHfpOc0n9QAZ8/tpidIGhSik
wBRg3f96YQSym05ehPhyadNbKOiXWk5Ycppen6Z4C23ZYje3VcP9YdNGSb4dtxWBbtcJAgaW22Bm
WbdqShcq/t1Z+TyBa3I13c8lUD5I3vs8en1vJeA5228Q3yM2D0YLrstp8OU5ZuVO2CBkaa/nkL9Y
umEhX8tO2X5rgRc1eikvQtiRbfeXinFFTU+SG80Kk8kTvwn6UA8FS59u+tnYm+K98a5io6z653EO
aNfvCKd9YqteRznd72Vdp+7/qY4Zr9P2iWXccLSWqMkGcloHKZ7lR/e66d7DrQFS3H5lH6lzO9HH
t+X3uasjsbC4boHtnbahHjobir45a7f5DP4kDYbucUue6YohYpJkHeGIQTudVO2yrR8jwKYXmLzR
Lut7rKGkduM2UWj6Zhf8NybeYwp7a07R1josNDEbl8519hGWuV+CaPXBKcDada9csQ6sSCXC/uFq
thHblwNdYum0puJCDMgd2sMA8UCwSReLcW561wZtYDpy4Qau6RhnrSL9YSuhGpdLcjy0dgasBtoh
84un1yFhfYZbnET/L3E063ZYx4NpiGFYrgubFwshrungedvTl8KPbEueDKpzdNffDRSA/mwa7dQ0
qB2WF7dTWEJWZBt7Tk07xBKxe4XnyGDcPChL7V4u6lviAHkwOzxTq5ksPFDVX35TSxv0QGcFpCwd
Y/6u5jQW1pcHVZTJlhRu0yKp0ThaM333JP4V4wkvjjCkQmAUEHM8A6aIAspDUyMgbr1hkooVj9OZ
oGQ/tpIn2dDQzVyQ6zuOKMSNYOAjrAq2FOQLxSxicoROeuAPvY8HfVQwUYML4OBMq/v9oWMoSBJA
EIrmkq+4LzH9Hh0NZvfIh8X/2L+ykbAsFEvrkZaMePDheh9Iva04vSxaSIJXPqpgU8iWedHMoIdg
bbKgcxFJt0jdAMJFkIzeybuLNa0DXMB5EMwNzsNoaRknO9Pl25y8/fOj+/zDrtPdskBIijFkWws2
ICgkCSrqbuvH5TzFs742xjv2kM3Numzs1bclwSclHOUaWa4qSPFkXhD9ieeOKKNk3qUoUL7ym4Ho
QBHAuFcpi7B+0Tv3xciMbjC8TFkQZ5mIdXFIVFKtXs0mar2xTWZofZzQJ1ZG9bB/onYwUjFoK1Yb
DZ0mDV4AW/DLMoL9ak9akA2SvO8f7CSXjSuGWA4gw+viGKva8MeUEaV40xuQYAvz96n3NkaA+pUz
bPdTx8f15UxZTOlaKu71CemJO17/Z7vJpKQhNjs5SaMdYkiUGWFaxwhXVk/56h8R7mVeMgXkY3Bo
sBql8zcf1Y3wg01cQKaarvevT9gPoyRBt6ER7wj+4K8I0UTKx6tksPuNYsZq3t+eumY5yScfAOiz
xby1XbBatQDPbZGya1Ji+U21J/SB5mVaDC1HNf7/cwy3gjxNq3OU0VHL1JG5mPrTbSEy6Iz/Z8Ty
m3afX0vLnca0Eua6PJPEVollJyDAWfTUfTQ1Y2G5+l8tSqiUeNOUvxa8d+tdnV6OY6mEmWj2CGqX
ioXMk/l4q8wWjXXdW7Tgd+7OJ5yts85gpKWLAoGBz77Ad0cSfz7wEbsw5NpwyTCaPnyXD5x+eCdO
/Hhvk5A7/lU2pfx+BK1fMAuRWrw4U1pWxRa/61FyNppXeWinPFNn3W/MRFvUhaTYDDpJq156VgDU
LxzUOai3rAd7Ow0+96lCx2Jj2bVqHG0Y1bPwPY+a9pTtyfTyFjbBbT+1GK/z3RaCiXDiE/LxXXfd
giE6mwG6KA26/eCEc/7nsEIcl2DMKvGbsdDwBErctyeiGzHeFZKtzyl97p6KAq85EgZu/hr2ACqt
5BEwHVvnxFdEWxQgn2DCDcblGIAs1WhM9ipwQ0kObb2Ts2qoEv6bvytFoftGbJZPCgFXYKOafZS0
b1eZhREwgLyVCA1HaNHJfgdBqdPSIb7udYT+6a3PknWwPSlpPzXC1NlAeHqDTWj/GV9c3UjAvu3z
6kGUgjh99XH3Jdmy5/YP9TxI/GkUtxh20Boszudl4pCUjRTD/Yec6md/GL+2jvNq2VZTce1kkw8R
PSDF/YBKmUGPd7BXgknyZjcg60WCEKgEHBMr9/1KTa9MqGQluqcq2kJ3Aztsb2qvtI/MpA35egxm
mDAsj6FCarBU1RGAQW83tBpY4S75GC1RZV8I5b92MNf9ewouL0RddF5qeeNTJMs2Wx1GAn99YCFJ
L7Gzl9zM0ALj7ZhFmU89P10TKReETQv8JvOCl1kgMvgBLPSOY08jSW6JMf/ahd5YSiyaV5z8oXz3
4TGpdB1ACQF/eTBo5o4n49MTC2DB1mEyn+Y/3TdNupDdExJnG3jZfCx2cQG6ZLF76cZh6KjFeRsD
qlR1coP6ZC21A88A2B0gai9ZebzqDn615tXhl0/ha1fiEYGA5Ng1YDPxju7w0e6WVjlmbc4BOeQ+
GOzcdNsVipnYwCMCGGwrV7VHRVo3GaLMqtbMTfUMvWQhlm16FtdFYVt1KytbjgT3AecR83fqbAkg
CWwLFg5EUMixdSenNL+pxMq44IPCKP9yJagrbtrM4AAQHqZcJmxIs6QgUGPJP2lby+Lt4Y2N1/zk
3Hgo8RbDlAGZBNwD8kReFw46r6iKPHWHcPHlKAhmK7NQMO5E3O3n9H0RrivDKgfewgblAPFtO3tg
0mqIUqkJ4DLG9lwUb4uMux35B4HiyZ9+VftFzNbJjJ1MoN7s8iQpDo57IZibkkMMHAqjcKkuUe3F
nHIL5qdd40dhdcgu4ALJuXb8ITlW0OuS4KGKblY3nJyGl+AP0+nOxvl2wYS6Z2gC6ZPhjHBtmxju
eHlb+TsaO5Hezgh2KAGbtoU5vvd9446r3S1r+oFKvl2pqRhCqwbHl/asim0VtGirQloArDhpjJgN
ZKYyj/WM8K43XHUtcgmmsf03pvTxsduYtdGmOzexlg2+nMKVyOjIdwh6gbpLxec9SluAUa6W/Jip
/mkWwXqBJGYGjXjSXMQna/f6aJn2ogWRpP9mJhf6T23uVYQxHyCi+DHYOv/+8g+qSTqOvbPOLKno
7Zu+NLHGbzC3fad9SSeWdSCkRO+Mwh9jS24UeBDe7U98C2Vu/ijaCwLT+gLwj8PGW1DK0nuYSLxS
ODJMlz1ruDifVEUV+G3roS3UhkjR7SzNhirS7R+I2yNxH6AZm92WdoqcwQ4soo5z1Ph/8lyB2QyU
wStVX/v61BnRE/97a8YMS0CwWUXqtnb/WQhs58+jY7DGjH9ow5vW4XFLG/iNHQTR5gn8ngeWaLhL
Q3PvVnw1X7TL69v7Fy70oCp7/FZM5h8wnwCa9oEPUeJHNwAUZDa6qVQv2af/JU4t2KVxrnxMTMo1
OnhDsehXwhI8NaoBITxa/ujJafFD2WFx05qzbaSyZg+Ae8IcxgFVhJSTbae4kZiJcqEL6SXOcLjB
UPp0kRMzkXfHmfBGThbTUEhJvfxIB0WedQwOF8i0706Y+GGlutAb++iIMbidtvM4/shMvcUUTSmm
ECytG5xiRieA3grs128kFsLewuoHZoDuLjEvbhxLhDMNAJYKd9iKQqWUAqMhC9QlFE5VSFS/mDO3
DW6Ran7iukh/Gnr6BX2m4+5//mcf+8gd4JiIe2hOWUG7Y+OAd+cLhmlYde3dLSiJjLyeCE0w7UKx
yNpsVG8ERj8Kz+1sPCZ1uppDFGJlgemEtNsi8yJ65qGon0VIy0FLDcW/qMCt+o+T2IN7bhklyjvh
rO+bm97yb0EWCto3UOhN3JbsNQyn/JH5qJ4OCEAT8D/U0KG8m+UXT+p26C50Lyz4PU1YfFV0frIP
7e92ev0KiS1AMgE55ShGLvOQe7p2t1/TzXKN1BfGtKRbcvk+y7JwHDclHD1rDnXZreJCqqMQ+rL3
A5dSH9WU1AoAQ81g0gQxc58ry6lJXUBmKqycl5zq//jIUlXafgwHgA1ZjXvZ6LsBLLAYPs770hiM
n7I+e9Th5Nxb1L6KTdg0f3CAyDQ7BzlE2+5xd7wJMFWCEuHifar4Ks0CRResnJuLqIzcqSmNSRjl
S0D2p12n/RKoE8CACn5uIZWHxPCR9MsfJt+7c8jzSKmUjIJhMQH7Jf00Q7byMJXlWBEXj/mWY4Tz
0zTX9U0PRtjbg9rw7WvXkq0soJB2LFybDaavzXrZGkQKzA8nhRyO3YVlyACs05A2E587NC/xVEBW
jSPOk3kOOEOWMGf0WZZdCHDtfi+BNeIwLoeGy4DsvA0t9lPMXEXReer7yMPQLZKJcFKvrz8fz1Im
DgXNOfXayuYVuMxedbA6tbLUNTRT1riWYBvyPjKXuxDCSRGB+QHCw/LTklwQ4d83OIjuS1PirfaO
7m8bUM5jRMBctPmRRY3a89I3gW0UJapqUkzfKryGCOP6ttjcworK7vtyYZ5qN4xjR2pUyZg7m5gm
usaCGKXw1xRE2KIwof1E98uPYM401ntCfezHM44rgma76F92pX7zj7wrYx3lDHbep3cm40plh4kO
wKcUGZYLjDY93rAb8C9rOO7T+/CJW/0Z+P7s2AzuZjNbFAViUA1RHRI87L/XUFlv8A2lpljBViQK
uM64nmwAaM+NXbcyPgRs00iQEMT0GpG5p4AAoHzTghdDM1LwknAfT+FZkwrMKWU2DjIaq6c2/IWi
lwW+zVfEi8Rg9lmlkrbDlvhQR/cNboWA8IiVtII6o5CIQz3h8fXRmxCke1vojBU1Ftw6Bqd0u8Tq
nPbLPWPuw2+m2PR73gfaCzXuwbpSP7tnaLUncZomfGDhFKZhVLgny9fV62Aw7PtGlOVprqFW0mTP
NaHKJ0cxsQeaRP8jt9BUr6nvJfStspRvqZu1HtUi69KrKXUhdmdKkxQBZfz4YZJtDDBJTdFTBeeb
WXcA5P7Hop0OImAGBUYfmGvUz2BbIolxuTetRrPGE/VPhqDFEJciyAy/QPxWO7fMExfO7ZCgMeXS
O6XbPsFLGCdARwGMjkDhDNqFK5LyxZEz8wLFINDKU6bd9FM6pmLgVe5daGhR/ZjDbFIdL5HQFK1M
Omy5tkHpz7FhmhSD21ppqK0vHINcU43xKFCL2jOQTo/gT4nU+xDb3v1v4rQow7MRNwKFjUg7xUAe
8SENS4Ko3pJCF/z7lP2Qb9ZW4oe1iOJDImlWbXNnCcnoTPbdk6w0I4XFN7DtoY7w2ZgNKwMZe02g
CEOc46R7YX3bYPNmRDzBd0A7Jxpj4s1iYUuZkL4I5AS6TQltrQ2Lc8bT7u4fgYCW88iAbqYA20kn
g8jvrYU5b74Pn6fi+bS0xGYzrelLt17AzoBB0d2fmjxFRRsGz/yOwGY1vY5aN/IGxDwKs6RzIaiu
n6MORiwHAL0U41EbAaZIWhVw9UHblmDXu38BHWEbjTBpM7CCfPYd4RcxivjeaGSwy5+eklzmx0Wh
/dqQhCAKffFykpRXqn1PpL2hWXC+SwJv/HDNu20XuUFscxn78ESUxYnf/jEXxaqPshnnSSOg0qpQ
dQHi5WvUo2Ha7NlAXieA1cWQlJonmoe3SjxqjQqSjaPt6vfAeZahq8qmFz2x3g4g5C3XJ5jwPIwd
DhiNZxGaPmc/SdnNmg45ezkWQrBNYB51wSU5KsrGlTdfK8hKnJXD4dNAwpXvYSVSdy+7ThiiyppV
VDbywgcyQXQYRkqEE6R8r5aClawCKpztX61GBzjcAYJCchREpngWQsemOJbbX8T+X18pZ1cuVkNd
pJpiCLG5yOWafjInLqL7j3fKBE5Pqr8nXrJTuRn3jLf4hI3m58vsg9fX7hQzP8OQtkTNPVLLmrne
s0sjyxNWE/7Dxu/944VQuvN+RFouMiKASLBwYPELPL0vYJmJHP9gcziRITgoGtvklfVBjtoeemxH
EM6Vmdn+Wxc++wB2yPX7uPOeZ2lFgtTsZl8JiqhlAFSIwN/mNi3Qr9+psHA38+ZH0BiFwre+xplS
DdCDMvKyKsx9YnQ3Ya9+M+eQLmL/SnmDFQpipb7YVXq6wERNLU8c+ngkbdM12Ar0yAySDVEFy/uY
j5ZJTMp+IDpFEiZdIrdbzPM/EmEzniZLC+pQHYemiLxP1udm4MT/KtZjZ996l2TjPKOeXd5kWY1S
DTh5Fukk45S+zW38zYX6pATEghXvVMZ92X9gOXwhgRObcUudI1esBAcmiFLWQoezA+FJ8AbR/J5m
FRJJqT4mYsTpFuxiXVCVFg9idbicslpsv27dm37ajFcbRK31/vA0R7L1rOCviZx56W6cIhCF7+ap
QknuEEJ0wKn2uFiCnur7ngTEDA51SXYD/onT6izMpVItzEu3FtziH+3MZ0ZZ8db0rDnIkrelZWi+
2e+VWqegBb0mMtIVkedavJUsOqHmGh2zyV9bdoAjd9mhCC4mgNU+gyqLGMu7T40hohvTPYaquD8R
KfvhTETtwiJNDO+GNTR4elcuxfvhMVSymX+Nm+8A7dWcxCywPu4qC5tmKenlieubbNnwLIe9WQB8
rOcbRu7kptIngq4MSlPzrsWNXgodErYFlbs8FDDToJDWzHyMhCwVbht7Ku8es2v10PiHC5h+twK3
eY3YQmpW3MCdFppTAiNYkU98qcsZZ8ilm6QWFV9djqKdPNpCReLKT12Cyl7JCY7XIHvZyXgMvf1O
IDKf/nhdWb0zWY28zkn5m7/XFEcRfQ5bluG+hoUcof27yWTJiygwZKZkIbXCVWiXgeSOZ7MUSf25
G+H1CqC/y6osGS2qTBQZIB2z8fNiDJKuyggpw4oXpm2DvT172ai21/skyq80rM4t8PoMrX95dJRS
01eD8mhwqxLnNvTqJAOoRAeeerJZSyc/qFjoF+1Kp2i3erUmN+IwgQmVjSwc/RKsz8zR0X1Ewfnd
2yH5Qb+ceJqTNJYREA/+iWuSqzVqO0Kyh5phm4AjqpQIOgCozMkZ6Mkhn32/kSsyCKcHXAIjSlJ8
hE0amHh+riyzfF+Abas2O0epOyN+1qpZutg+/F14xjTrjPK8pkaWtNwBxaVZNvSHWibzfJ+tVUN3
23LaBntazD9rqFL0F8IpFapMyFBY6wBlGDmZcGl5GouicByuSAE1sKw5yyx/KsvPy7rB62rCi97a
K7W5+CwW30VXtl3w80gEfnfAvOvQ18bvpt+fbO/juj8I3YTOgJcwVdKfuaZdafC0ekUMHJCAesYO
gIPrY2y0NYtDfolUIlyacH/mfenCMpTdyiS6JeTd0XQAU2ex5cdd3bsMWa9RDN5IbxLJZjuP9vAD
5hdVmIclwu7lVOJYW8BBlW5lmxK4UxvgfyiKYpg8w+lRYqpJmTsEn3hRD/kkOO93ZU142HSW+wIQ
0XeS+ByRDlFLKIqstH2vFZd50MsCiNer/cK6jKDFP3MzovWBxbCsmqoxDLb9hX/nkV3/uZEwULq5
d+hWyD8yYwnquJA5Tarx15G4uS6Cr2oyNXa6sBlCILOp7KaKIOSZDkM5wHt/pG/rwPpBrg10yk9H
yK71S9qxhPy2kFeSIlSKnS8H/T4/wQz9VYJmjbjXclA5Tjv8tzEgcW2lQU2ug1YoXrynQvl5Xq+P
1FJbneai/Xl2S6vnx+jv0pRLYdm5C3Vrhv40jlYhWKDSZmuPurF4N682zPVxgV1yxP2t7GR+vXQW
PqDOE7QxpB3edfKD3ERdHBm95aW5VeQNo/4MAEIdoSr/P6r3hv5Pqf2bQLolKCr6ToXBquuUJqb0
8sLdYLkMXzFhSlt9ZS73IbWglj19Xsgm02mBCcto6eCH1zHkChbSuZe0yfyiNLjiQyf4NAf1xA5A
fopx5ajzwbL7e4ZuV3XjFCaJcb7iwv89REs456qPpZIsmSsSZYEtnGXFTovC9zImrKYG7pahtf/K
JzitaWF/zHmM+WtEOHzDhw0J942DWD2ufJLaOgUE2BAf+WDpbTD6ovm4L3U1FXUMHS/8tg+tCVKz
sbVMTi9F7aLNiHz6xF270XPYdk/yke9nxFceHqrf0VpiNoIUtAcXe01InEgPp9njBnuvamSVhfam
EqaxcHmjl1ti6MKJT6i4QKhVQvRMsCnVG4+RZlspJlGrHjaBMccqwBOuYu4JyOgFoVDBn2AMl8Pk
tBeIaxzuBfPHys9an9JcyHxtW6O2EVSTakGYYBH4Ju1GloE3BZgev64j6K9LDlQV31NfUBPhqA8T
6gxZthfRpwrnkrzqDgaJL2GC7QLj1wbF+jNG8GMXdMQ1jSl3s1FQ0hOrUYfwEOaU2tbY5l09JXpS
7SEpqD+kY0HLjGySKB+qzAgOJbi0DTVlAmfe1qVqhjJZvcagugCe5o7LO+dwRaz6L8UPJq7SfRdF
E7BBGeenSkFafVdiz0EJP1GmJYWWvHkKyt59egi4EJeucvUBG7TI4KEQUD3/D2TC0RfweYg8yEZZ
fV5Z+k2t0IzbJ+CPCSiKpkG0/4DtKAVq0GTrbD191c6NbblHKN2M51WgJ9pH+aPYDoNBbiGC85JE
KR/6dsr7q4M+i0CPQ8TwgvAg3uKPA30nFXlSSdOIoLFqu4TSVaI6AbLkBgN8lJ45IV3yp1zqU1cs
bh2hvGTZ0DkhWWKXkr6v23f05RSNipfeW1bM4PFMy08jJg1YArLmXnRxzVPxNQeUo0IEviCdxadR
kpB6GdjM4Yrzv6nvpdJ5mQNxRxzbIi30TfwpPxx15k1m/t2ttEam1wnVz1KKCwp29dVdlHOMAsRQ
yB2XjejZ/pkbuVZjY0W9HGUf520UWLvOD3iVYdfGZcgtAgedUo9x70UQIpux64c1YiY93Y7d7o8b
6n2Bz0pOmmBU+Vs4IFUvbwuYKnyCc3bNz2v3zpPbZ+jPeBY2p9c4eNSNLPpkUOgQmrvM7r4in2/F
/CZdFLzWtuzDCnnjK8LGIMSrxcEdH1bm4W/7a9VDhuMCPax4hKdoVzEvSpSZt7h/VZaoNqVc80y6
Zi90T+qEzSjOOrHCXfLl+5/WTOdh1X4Q7aDER5p2t99XKyGV3wMcUS9oOq0zzUiLQS5wOjNInLYX
LThl3Z+uhDl4lcmTeguCJWq5AVdKhhd97eXCwI4/f0Ye56VBBmjkAUgYtCNjCKNbi2XOkSJWN8eI
HWf8QnsCIG2DtYYX6jMTzUbglxHGudD8wQWNz5tEGtAEUYcXCBiBAfTFVy9Tq8RqDvlW8OdyvX3A
eO3CibMhEGylnnaluN7gvgD0zYv3vstJIYshAeSxm6siYFWfgC99fjk6NuvnNuZLKGvyvnHpxey5
9UqIxatAoKzOaHTesnj5b3+xOwo4GVaZD73ykSeH6HQGBMiQA8DUPEpPXYa+fB8gBH5nD6kg6zj4
lJvhBH6EZVJhmSlvqTYVqnhljsuRWz+6k18eNPgoVHMjdU4toeUWBeSrELJnLdXq0OSIbEP0DiQs
oWGcvzXEmlw4ywjxlaUyAbEB/HDa/5qG5W6NpWEMkdxrt6BMe4vKucWEf3bteh8nxJhjooxf9uYs
z5X9R3+04gJeqWVfMJ4FxeC5ysmyeyXC+YsAMGiQJu21Nhn42bFUz+jfRmR6eJcbQaOf0qe1xTej
Z9YbuulbScZDGPi0BVGBIE7r+J0ety5epnyO56BxM0WyQWVb6A9kLW7wOriCjHWGwhptbdcEell/
YbLiSa9x0p+36+IVCxj0OUU9M8RX5BTqn+sxLZjbDFlJNeckua1BO9WwTtpNczP1BtfniYaNKt8l
TzGfzEmkpEcIcFUP+SurmpZELmXk5kn7gMadBVU6uimbQ1snvbYT/2Ia91sipgNf533IdUrRTIlt
/yG8I1w/ZIgcxs0oWyLlgBMYHUNnchmFCIBvw0QRXC+F8LxilVOgllsB3jcYVO6jmpV3B1dMa+gh
GiOCZOKEhD6epoBj2OeGUc6/zpaUy1dErM3WHnmFTi6URaGQoY/++vomE3EoLSfxUozNm+fWqB3x
3q5+7O3+2uvCAwnT6dHF5BtWdslbU0ODRXQMdtMuEms3mBAlWy1i27ESk4455jbub8W7A0xVsuoc
/s3WYgFKANu5l7FpUhaqNq8n+gnhK3ljzKoeKtyQx+IMZeNXXajUxDwLiOr9NRV8Z7D8flOj1cMW
hGw/w9XvJ5ihw012yuf/emPyAXyDxpfikB6qasIlILF1QnvMwmrDhT8t+T3r9o/Hdj2oxmo0AdiU
yyZCYv0QSXlIN+8D4WFA5m8as9m4qXNR5/scUCJpTu4oWTdpMiqEjZawLXDsFAzqkWJP3W988Bp+
pUQbn/VUadJN5KBcLqw1leAj3UMl6EB7Fng+/v0QeHMvIDYQq9baADFH0e6feDFFrjYMjwOSNV5E
KHBr7VTZ2KuSCaOufyu7kYCkP01XHCeRTAX/ioMVPIfiboK1FxqlUxGMZjR5ZpX6ugb9LdN25hI1
Xd14QBwQw2nLgPg9PLh1oQZSHfcrDo28kz4wChg+0auWa7V1nV61K69Rj6w5xs6SusbUZ9H/tJTE
mFyK/F0n4ii9/+IIe3TTlOoxOF6xFNcgyp5Vo1sEpQARZvynMSi1n8iKnDpiUGR2P7w28dMi53Ik
8CSrJDRcsuOnMmtdkhTqAfNm/z4wZ0oNVrfOOcbSRQOhRLRWmnI/I8z8rsp73zDwILCrWe4fgG9u
DIIg9YUsgFzJ6aznKGwjSeSM7RVwh1IRadb29ZoYlGFwvJ0b3bDi/GbSgCOeSeLm68IM1eSyD3i4
BxSqV7xkKNNGlGEyxGsMzDhbxx07dpT2tMLsg44qV1oWVUexCjfvEp+hZcMq/JSTmeTLIMhW1fnZ
wI+EUGr/metDjreMyvK4bn1ptYiYTDip9raOG92g/Kffs7VUqmKX/bphsGEORHmdwXdK1FaX4iTo
AXzqZS8JHn7QCMqykQTLVefT69FUXhHINsuwkF8+Y8sXwnDnuOaDQed2rlpLXti/acroy9xFr6l3
sHcSVSrAmDsgwxGOJ8HcxCTyw3FZi/uNKUUeqeoVRfkGZAkdas3UCHbn9b0kLF86vBQ0/pVo9tdj
TGcEu8d2Q0IL7KKwDGgFWoqIreVRrlYbeZs8Z1ojDB3loSPJ+BUFNc66pkHyFd8lYt/su65u2DVb
jFrilUYqls8mhVvScurHMbTiAYaSKoZjTH0VdKF3w2ghquXHkE6SZ1J7AILxQ0ereVQmvuy2r0R9
cQ9xsBPDAJ2ufRpeJaPa1Mljw8L6SajiWRTb8p8kO/Nbrq74tcLHinog2Txzf/K5dj1WHiyG3eut
i2c0HRQHP5yvB+9/4m6jun7vM9QrgN5uNRMZITNo+O143/nkivVewHWvEWPWYg8jfi26RMXoKFd4
k86+6YZuTHAKv9abWpxnEGjc3qiLqlv7uBlwO0QNQFHJObO8TeFYHBVIKoWVobFr5YWjgd1Z4Cvb
ca2sBi8L8TmYsKbshpy5GaOEd+ShMZBpHExJ+hNszYUnS0ZiYGgwVuHN6ENU6yZxXVzFiqIuAwc2
eUm0JZ1OO0lMV0DxxUssEGQiGWRrPbWDq2kyojT5sr01oDyhpXjwx1dSFJXjgsUQ/fj+XJeiMZmE
cwBDMwZ8NGBTs4xUkf0ura5N0NOgT4QfKmTpL1f4NsZUsLqLXQQ844vQvjvtsZifR1LUyrQT9oRt
Hb7tFdvqrPo33pnrjITrgIUl+valW02UrqNThH28peN5kaDn1hUpm2JyK0S0Y85AvbHzQgCqneH/
NPKYUuQdDtaMReY8c/oJw9/+J2K6jUZ6LqPdAxZNYPJPOgRn0MnXH5yB7X/afGjUn63FH/OOw8O/
a3rwxF7SjfxClHq46rI5K++p42Ef7D4AgWZvqU2HZMyZ7RZkwqkSZCYXIHnkZW2Uw2cQ8r4IRUqJ
UIS3hRTfbuXSG2gwaXZAb2HkRI2hYlSTCUjxvN2LeckQB/5fMtjWj4Gf8FU3irkds9C+P89idv5y
iFILj8CYuI7UJ5qWVbs3DQV9F6+XawLP2oOs8GPOfmZPB+gg7nzCjKujYcLbHCQKqMgLD/lns8gu
+nmmGUe4FeFntr/hw/Ic1mZTzWs+yvQzRinhV/9AP3hZ/ximUetWLFRmlWyghMisnP1mlg2oazeW
8mKLpJt20ZB+Ud5RIWPIaW9Des1OJ39VEXpwaWZYlxiEv8HWI8kxdhLoI8fxbxSk8RVETtxrqP1S
444X9kHb0pSq6uiTQVnqtEwTYWx68ghTugXtyOwoxmLHVwNzk5BDAaEKv7MfeXbbmowBgjJkyydQ
lIMXAs7UfC2FApJWQZpall9+yZRrjvGJkHHxiWqbJOVstRE94Q+kR9GFQwFmIvsoBi/8k01eykvh
8fA6n7MUErAQir+Rh4b81I3XrQzqb3wsieB+KlIjN46va9Wv8Zr11jj714XDh7QnJ0CY+whCXM1y
38hV3BTZV0wmci+usdyZLhDfWIGugcqu9UWIbgSYn793pXnlCzbbt2GexRz4WR//wah8cxgaJhHV
Hj6uc+5/RhQKJqRMT7II/clv3P/LbrgRpS4GHpbwKpB8ljDNh2hGqMECKoJQ7xsMrynvaxwF+Kxy
cnuooSSveEX3AQspyDOMOjfHpvC4iDNFA7bW54bt/YTEDGEd9BKEdUrzLer24F4lH9oy0oHvHzbw
CcyXMZo7X3rQXcylshGk60p2vZyvfoeoPIgpgM5ypmQSSpJIqMbaqMPnW9+U6Qvg7JuRxHbyzu/V
7yJEdZ9QN9V1RmYVhLxS9oAFzcQXllXofZDT0XFoPy3OMq33yVIEihVKUDqSjkxoWFqZCIAhL/UX
FmwgflvDgvLfS5krH34JZ5E5ysLCac0JqTorRVxTn8iRDwBsuX9OOfsFHGlib0mWuMXEEPQ5JcXj
uszB7JVl6tPWfGXQpBm1Jrd4KmASwAiaMfOndg6AubhA5ARLFy5HsNx/suKtyUrmcGr7Cz1e9hwu
E1+8AH1mE0SImI8lnbTvOcO9bqJGGQVKbTl7CBEuigs5qguiPeNxCw4+zZHUOdsI9oQUXCn/5skx
PkSjTWQebRAHfPaTfboOHMtD0xrpsKgrv4IyQDysQoZxMQfza7ROxovtWAN51BbdV40Vpj4nDLbL
TZC69rGdGseubnQ95Iox5cNJFNb0X4t1xnoTfGogJnBBh0yytRSs3qNhYe31cAxjL9qiUbbwMiQ3
HQ2Fls2djW3DLFtWL2XbMJCXtpQVly8SQmzX79ml4z+AJNpV4B1bB6QROUypJOVJjqrvESDwj2et
92oA5NcKjWuYczu298DZvCrB+qXUhtwBb4U+/m3nXVtIIDRb/hEnO5RY9KU64r22qybifeaDvZlG
ZVCUxmN5PVcd719xBXk5lT0y/umvTjYSmh4/w9UYkUuclWQvCCxhIVxfT6CwWthU5YJgRl/hTA8y
8RtshSQuhBBwDkP2j9bQqaeBn5eOp4mt9LsYW/8XiKYyAMHbZtlzrdcmA3ln8O0MSS8GzZnqCKCn
09K4k9DJpiuQZWNjquqf5ib9HRao3ChpMNGleoIbVddHrbekmDNDH1yzZKUWb0XyBbz7tP3Cg3PM
+RSjN+NtpI26rW7YN03xJK/FiLapU9sWmyOdY3lSzNmvqFb+kCYjZBCp8f1jcMVK0bmu61GsRXl7
hf+PA4EIt01YoQ46SFdy3RiQIhCt2rQtq5+/i5FFpJ/7Ca+bFPPSZIKcQxPy2wI/P6O0jP+D4/yN
ba8UwGYDrVAlJTlOyFUPpey5Or7Kb/rCaX3oFLwLQWI7m0+fmyORuJMUclDUBHkdo7uQvunnxM01
RmQEs4kF27VaIqSZfBVWO8pts9qcFvUmSPziPEKmn5yv6QTIKuZ6BDc5qrtghkMCWOp7KjOLoXc5
6b/3yFY91FrHVlVJzoB6Wfb6mtt8/faPeDBgzvvhxKpMkmy3orT+F6WPnO+kRp3FmVeIwEZWE4oB
raCh6YePJ1TnQ6LPRN559/LyW1pRZzEjy76eF6K7W3a3m2+LqFrkGvHFOkDj9IqYReQoQA1ky7HZ
kciCSriMVlt2QVRwQug2JbeaZfcJbpD9rP+TcmKJper+js0mBVALl3kM5Oh6O2wLYerbwav+n+Dd
u5C33BZpBoSQG0WuihvFpzlZ7pLvj4AuXLx4X9MH6fqnX5coloS7nhOzYCOshu/nUwAdSX1cEFx9
eQ13pdveAL7bIlD5lqQLa3y0tLFlsZ3Omc74WljbsJMfcb1gE3pLpuagHoO1qjdow+Adn8dzbaV3
fAuUOtIywTHUsCEamsc2iUH7whgq9BX3/2xperCQalDdzf4uRSA30zxjH2aqWzvRiE32ZUXI/u1l
3AzDBBlUGCAigwEttEJJ6G93s88PdoIJkIbX7bzc+GuOfs27YUupbmAMn7DHN1b9Gb6kx+EIkTru
sN9sjTQN77gdf/Ph8pQTfg5X8zPBoY958bk49TBZiNh0cSzPozteBNIkIz9Ax2l/RpL+0WntllRG
BKk3llMrozbaQtVkG3/yiK+1y/AWuXq9tFTsHNymeRRh55lUFC8dtHHL5S85i7VZcGtvB8O4/+9y
R+9rY7OFaj4DzADMZC2cVSaiVMqovooijJcslAMTe5JZFO5xTpTBe3ozQ3A24t4F6YX4MSTt5gZz
aKMyw4dPqkhPgS0puis9+Hv7ZlGlx+a0ZbqsrSO9StxKTMuEeneNzUpUDFNi2BUbyzBKRnBzTH91
QQPFxHxZfF1hpmoac4d41ZAzBd1j/gNIH9LmpRuhOTL42zTlZgk8nDh9Tr3CbFYPcnamUM230DO4
SXhCZhzdl9jOdadB19q/ue8V7NNYoY299eL3YANn/aFq0lAWVW6+VqienMtZLiOQHNiEBQI+1y4g
dYJ6vOW/WPm3RNUqBGu0zSb7UTKliUZolMEmPb3IW21E8G2KI8ak12aM3ING96z8XdemmQW3cw99
avL+akNfF9FuLvWQqGOkVsEvdI5DTmXm8YfX/PU6Gh5K7w0klmPp6tptSNFvTbFqciiWCarss1Dj
Y/MRbzOFucqeV7/fqF5IyhZ7xMwQqhh9Z0fsxkpBsuy7altYw1tvsnyMQJlq71niYf7AKAnalxvt
1s/5JvLdzFfw6uswQqAaWJs2mV1XcZbuaJTUSkYRxe3c4yQKua09mJmRoDjnDcaOK2f7Okn5Jjze
UpY3abXdbJjylPpsQHVjS9F2pWtscx6xd5lVBTjwoCoHxxAzlMTVAnW/m0xOmO0y11J/RZyIM3VW
ErKRmbXwthpAQz1d2GX5kosYhzWI1UsV9B0/yKJ5pKWvtO5W4J83TuzRb8DVQmCSOISshYVbQsla
T9JspBzZLAYw0wx3qbCRHeSeN1I9gj8jAliuCWLU+H7q25tz9Gc9YuX3JwF2gjSwKMNlz4NBxAkN
yKLygpLzA1Q8WgS2K2LhpLJphqHcbTzNAOzarxeRdPy5ZILuUKhiHGSqhMa1SxYwpVU7XEjruY7l
9WP9JQg5qE6bCfo5+EN3qjlopJh65lX6/DFUZLiZc/Lwk4dcnqtNrR7cSB4OjDt6S/fqGQyl0qNF
YE4tsi6lJJAPtyA51xrVZ1G67G3ej7frNbUjcumPw97K/PfRe3GR84dF7HWxrVDYdWIWpBRE0Rdq
/SIogp3DsO7RsAUJ/7nUjbcs6DJdDQKzEn10fviFg1I4RSRGYhZ4WJrLOZuAswHzGnJC3jjIeUAr
oAaE4mgjrUzI9RzpbDVliCebXQBON0EKFSu2LLB7HokcA+tKXGlmtHTkTbvBo4alKm+ivcXQcNy3
px1y/o0CQUP6sddIf+XMK4wZGqSuMxwpahTdS9E8wV8T2RWGNxE25Yk9mLeoe/960TZ/nnIGxqO8
MCbEhRd/dziu8QpIaMsvl8VSIcv4U0AC9UCpoxZ8KLx8Qbzkr6ridOjcGfhU7RWIjgsoUhLmSFpq
P+8Y5XSz26O0ChgqHNvKS47YRhuizLy7FAFlaa5LQWWdqpMzESyigtj+sB6JZNgu3JH2MTJKvbt6
fjAG+GLUmxWsC0+BYH6zyihivWCuQd0hkDKx3kwwuvaY15ZJGBtyqd2UcsFZ2/mqeWovLh9BZZ3F
MK+iPmALGysj17I6mqEzThUJhuLefA5zt5u7XQPR6697IK+mq8kA51AhJFahOi7N15yZv59pf0u/
AapGy2GyIrovB1whjiryX4DKyXutaVGARYaPqUXG16J7SG+KeVhamDCJtH9dypGLi7VveQCaZDLD
+WvtJ9q/1v98wQSFfByT88Hh9TJfxdhXx78NH4fPgeWbh9iWYip21lBX0QM4IAwxZio7JU463cFP
v3iW4KXuV8CKQoQffUfnnpEj13u3k461O0VvRNvduf4Mn2OLaEAeb+7ikVIj0DOUUTrk6LDedege
OmbA7AWJYJLDixDRv2f2TKzAkOPptDUXM5DNcvhzU6aAE7aDm6PtCaqCOijm38hDK52ZPi2M1JJs
AB39zf8Zj4n9yGwjXL7jAGV0mh2Ol/HvIbC1XAAIwBk9FcmljAZSJd2OnUBqVRY3vrGO7M07qajh
JJnz96y/TVHtfGHTbLxS5kTPzRQNdpfVuNYJ6a+kQZFZqhjmc8KNNrK0jSmQhi2mpW3893hJrAPK
VhqNzfsMaO+dhnFtmLfDVRbL0nEzUdEIxerUZ6MeyMrKd8XlBT+VRb+3eCzYyyQEIpgSId16aC4f
X0guS7N0vGm7YGNaPoVZDGTEkbFs3wzt8C8tct7DK8FulbjU4Rv33kybgnnJElON+w6zqQ/jZcSb
AbuIwDBo2Qn9MITKOrj7MT/ceqRsF5/tkNhvMLpFktgo/pHEh4Y122I8rxQDZ4HOy7R4dObeLKSS
DSjcl+W/SQnIdX7LcWV9K9uRlNPcls1gZgqt68rRxY3MIi5jmUOThU1ZvK5HsiSFr6FP2JIQvRHR
utRP+zlpgGFnI5SBqDeaJIdjwVt2IpmWK6Dq4yWxLwOS2iORemoPIFJgMG+zvhsKu/j7DEeEJ0tp
12jwidSEcHIHMoNTbZguqbDYkQH0COi7LbkRKFwYO1/uMWNWWo+NtR1L3ou8JRT2H6sTS9irX9C+
x9HnKOzo7Y7wRm3HnHyNvCraRPi3tIm9Ym+x7OGNhcY3B2ZoZx/Yg5QAApvimU7sdLFxmhq9sNlJ
SfpMeEOAxaA5eQR69heom++oapw7hT84+xurhRqTZIuMS/idp45YH9xstk9uVJGsKERBsXfLV9bs
fZttc2PrbwGals/N1odRiIz5iq6fgKdIAF9nHUbb4B7afT6whxTo7LECHO2z5Wlmnkd9RQcXpQoU
ADnFoaeSU+itF6SYV6Jz//j3G2c0dY/eu2/reIG9tMEcZna/BpagDjX1sNfsL0KpMIgFk2pyWnvK
6HcTR1boT71K9Coh0+bWmeEncEKEqs+B8NVVJm99v24witA4GQiZ/cRaBXoxryqBmGXZXxJhFNfp
YtdSM2mpKvbB8v8sFkUV7zL8pxz0i4lAyF/cp2mkmOcE8EJl0Hew0eiAuV1UOQ7uCvROCRpBgM1i
hgmOHOBxA0igtSDFKkMVfLX4Lsz6BOAyOBMlX9SHkxBeRSKO6B0oHYqme+0hd7jRiWA59DuS006G
nrlmc/3uDpdJowYjWn16JVIxBWkmRIGgcx3UnMtzMsZZIuBoKHR2iIUdX7k9i8g87zuLiU9IlazH
sFRCQY/uSiKM5ExlyHmxS/lSicuSb70E5eqluQyomnNcb5XJDksA6Um0RF/+ActIBQUvvboibW2D
v7XIGobC3FVMz01l9Z66P5r5pJNqu4iSOJT8dn2iIf6w2sjm0DovzBKilsxwljmrw8YeN2P59a+n
0tCCAN5Nd2QCLB42JBCRadPHrb4Psth9YfOobgJtJiySQ6qvUflRH8jzWM/mwDb6kLMM1KsMr0Nl
Fbg3K1bU6q5gp+nu9f34TgkzasmHdyAAoPFPrnGDGDQYu9rWFsqWIrWwGuJTbOdtzO0td3PTcZ0k
Ih/X6fOWZGOYjqYMpH8yc/8d2fMD/xz0jMCbDnLyNY/ksVQYZnO/EaeigB8nGKbG/hX8Mma747G0
ebGOGWWxYZx1r0pTRfFfPouUSyZ0fukMw1FVl87KkHjfILfR9i/BEA/w2NErxo01S4FfvGx48Iai
xhqaaBtpnVR9f8p31VNXPfiRMGAbhSNXEUUDqD0Ol5ut6jKxUy+jUrtUHQKEOzjCWpHgdE9kyYTh
qqwxEvYUrMsJLXZhhGFydmC3QNMV2Rp2owbCHS8pQTVsFbtEGuMS7eaYbnnTQPz6GqiwaU0Qfwek
Ru6gtil9k/TZXbanwfDybCsJ2U5nrDOIouP7U5+kjVKFP602ob3EQvVb6mMgXrfkoZfM5EaW7iL2
uJ44XHNiEQAhu+NKP9if7LKEp43xABFKy83GLGZ1s2szP/NseVAq/5q8Yz1ZOi84rSatzutlVMZb
0eFLI21bmt9GcJezSQE97s1BPitMHkCoWfcxeQWa3e6t7P4VXWpTcXhea6kh334jRV98AmI4HpN/
7sW4wnLQ5hO/M2VdWY56oq+/Uz2RxACJxF10fTSc+Gf8yA6acs5KIkmKdEF9xDc0X9Y828q32lo2
nRXyAf/3S35UGaUrx+15aPkLN5td2OoANvspgLmSEYo3VI58XEWn+xsCSmArQV9hJvQau0YrO06X
8An1ALjAomX8Dmbr0Pd5Gn9hjWCDP6GH2x0xFbDFnlpPd5wwOY2SN4t7Ml8f9QBV/zEkA+nKMrS/
ShMoFwfvLNw/94EF7RSRL5N7gVk0MEgnktY8p7WlBa4WKpdHBzy+lXh7CRf1236QJFUgn6Uv3nE6
/OO2mpblsZpuPN9+eDG7KzgI3tza2BHAsdDQUVNfIoXCEReKXxvaLitA0tUONCDKAZCa5erZopaA
n8sTvsHoue5JbqbDFYSASCEMCMyNvKYTDne+WdjXZ8bt9JRFZSblQH8en+ZKz/92yvhjVXn8IKwm
2cFv5dCUcPOKytgGcVHHgn7BB+rr9m2NNnDX8BqhQVXRWJAFFQOwFlIxydgS/RSlF0B/CzzNmLC4
uqyfi7s3n6q68sBjYAI0ZFXy4n2F2mcfyull4AN9PWUk7N/MTVcUkCnf+IUs61bxhawVXrsZZLKd
2PG1KnTZdyvXl4sV335sxW/GuE9MAAehPPABIyBl1L4IQ+PGBpeNSh/Anmh1PumaKRgadNqW63I9
DWsb88hagSCbgk8u5P42K8x1Hsx6sgKpXA3b8Yt+LWECOqrCDiI6AbOrSnubPTBA6zSSiFmWnA3i
BWUzsAWkdSyeDUfzR+UlH/cyBLOJz+t67elNPjR6e3ced6Y/e1zU8S+LppzxIdN2eU+xigPJeWPD
hNnZLVxRs2MIY0VBgcHm23DrR/psaanFQwwH+24Gid+IuqLe8kYr3xndxVqHXBFci3oG8NyFWXQy
JyUDfsF+qLjirdI3e/wvAu/R82n5nuHCsMeiv6aXklzeMBEgQYpRnvrEUxNXuAesNgMr3sc+b2bl
9WFvCpl/eFKXPWJFxsBTuSP1Z/bkDHaKTZZA/wS1pxKNn83rR52efTb+eHxlB3SO8sFV7QQIVRxt
3RkVN7PBV0jBDEG6LiHicStd1Il746eks3B/mGBoRNmrRJn/oO43HMyMPHUWtNNBpGE6FzUzBNs2
sw+xgqhyzY/L9LBiqJvMCfNiw/NokKudUbe1BNKeh27XcGtvORQhKed5x19MrZdmFpiHBGL3We+E
XEfhuD9E33pH9PjsI7MPqZ/DA8peCU1hLz2uEtZo7X73BMTHyOaEBStgyXObbMqPcLObn5GVUKEt
iM0UugjYOggE95zVikdf1NDokvd13QkAPQmweeTzs8lItLlNZYTlnPv/enzzqqqVaPmE6sbJV5Av
i5vmzWD4ZmQNY8UjxT2aw7uhu6GrmEbN6dbiQrzvuwGAiRShOkiB8BFFSNen5/I1uH3KoLdohQxH
MnCWOS+C4slFBUctOD6/U2FJbTFY+4PSCBTMcC/0m//Ngr5X0jU970EC2qGI7rjPZCEYjWjxqjpT
M91Dxa5ENWnViGhxk7FC6AU5s5Xn5PXJTI2X//+Ul2Uz99QNID6vjqLv2Unx2e1zS1+A1K8tqos+
DCqVxfvijDvk8CJpix/MM8IK3mdYxKio1KSaVg9QcCvSACDNINrlcsAlRE2Jy2mzqcIX6/IqhoNV
9IbyG4yPqCDZDK66AY5c3GXQuypNXSVgYiAyMssfEmGOu0wij99ftw6n84pIBT/GEqX6Gu2KSY4g
wpkfv50LxcJgIOxnNp6lARp5Cpl8Z9tScPKH6iN7PtiIUVxtiUkXmSSi59vEnjyKIxovB84J/EdQ
UcJh/Gn0L8Ua4ZywHjdkZ34zHnzb01irEQok60DOfxi2bMwr0aB4ynJDQhAGHhPSxxzmTmZynWMj
kOvS+MPpa2LJr770B77J82YVp3y1a8Mb19wnGbggbmPfZ7DW6WTn+LQUTLviKRe3aaqdgvXmouWq
LHNeJSU3j8HtHjVGR0irZq5GbDUnTRsdho3+pzMcS8fPWPo3yS8V0qL+dCUmTHf3XvnYZYyiUHaq
kkB3osteY9lyB2QM4RK3qGBM9knxarZCqvPCEun298p3ly5bJwlF02abF+dxxVnzUOeawuKo60Gh
4PeW3mUbz+ebCCr95yJ4VB1PMqyZ2rTBNO0qtXwI3Oq8ThVV21W0gK76DA++U5DeMR/OVGry/A0P
13pggETQ001ULWca49Xwk4HvJpFXStoEOE6w2tWT28iH08HNbaUN1iY0LLqB8wnKGXlZEv8rReVa
6FVX2uaG+pp8CJXtU9MtZ6xEb+RyyXYmkNFtnTdPwW7BH37kBJrPKl+zkHEwDmmjq40SStA1CQaE
zQAc0WM6q0T0PdBTEx15IIgBri9TNWSSeuZMfFsT8CFIByXXh3wHXHBoVtrpw8dDPGu263IvnMZ4
qzsUep3ufXE6Vn4/d/ack1cno1jkvtXZYPAStf0zLepUJIIH7QPFg8KmdJVd45BUfFHGk6y+3miC
p5DGLJ996PRoxTcZIuZpqCFkCXSJU6cErMGePNFqu5yMckRABja7VG3rJwQP3jWB4EtECAVVhq/g
O0y1PKsUjsVRwBrCpdGdt44pBppJHe2o/f3aRepabidSjCquV6DUjMGiXsYGI/VKfswDikev9P0I
eXXgE4703Yewa3z+eV7V7Oxu5J2o1s+C/VOIjhF4riQdW9MkrNFN0NSeA4K6D4QKOf11MuRZPQJl
mTt6eaaOAKviV0+1wIxoL1txcCxBrEtHhC7BPAgWocx0RjjfT59otocwE7IPEC7ydjj7d3WzForg
dXeXu0Vem6nEOVKOOCXJxF8c3kpTSo9lRf91xX0m3QvQKkoudF6qhNREA4ai+EBZpIdNw6ZLCNr5
gw3Y8kUEmuDySpb8kD9p71FWtq14ojUHxZQPBuB9Z4FhiEpykRjGp0LUeympI9FRncMUo2KekB/U
ySGw2KOHAAFCB1B5HF13UzpAQaL6ciTfp3udiRjIlyiKcG0Tml0Q7gVpYawn0tm1cRmKP9lMTWLL
FCp+4fB4k0D/cJ4SjCvmenAUR8ubSf1EMy0AXRZfyXHc19fuMG/viLxzIczPIYCxO5c5vUDMwVhL
W4oNMHkZCd4q7LSKzxaxquu7+aJfb/D1a8UDIfFBA5lymiHnXIi8i5HYNVOgkQw+DZ5Dki/rTmT4
AuZv4zHpzobBorJEyghQAoMNWdF2bfeN/fcBVJ9DuW28egyFR9Ko1+NTOrlcIL3AmE82O0KH9FgZ
K9ITo+MPuzM9jJnUrkBRQiaFgb3B2j/A2D8zinhasLVSHo5LnBPv2zyR5JWtpLlYcffkfZ6GYJrg
buhJ52l3DD1mbPl4GwqAkQ/bJqM8mromLzgH8epdF0hO4jjEUh0aIJ0hkH9tBYAJ+miyYQZqChiH
lnWKZXkm1dvxqTuTj80OKGD7KGPGmcuWOiwb8enjtjMXKvtDc+xST3SH6ZMcQ4r2gUnZzamxNZ2r
BEOhyJt7g7GkAS0sFUY784RjgYewcYmu/euuQqPruud61fxDnK4u/2D7oMfYed+gkcI9yHOP6hkV
FkXpUE3AT7zMTnzS+RGG5ZQdRRn9+9iHuJZts55Pc/46iCPzC5eiU+yEvvicFrZpOsDk7HPysCiN
vD6VfHh/D0lNTR6LGRh/BSkFOct5vuq6OWCJHQqSBi7u4ouCZDsOrOsWGt8SEmyRNFZ14T8gqIIR
1vv98YPUd6XM8/0CSt9z8zqAMj/zxIrobJRJatNrLLVIdlsfoCfHEVbqbCJhJTsRKIUiSyfs9hLg
vw/Wz4RSeeWRbZdkE1nj1l0b16OeY3mtMoj5gLSh8bUJbEh6vD95e9TACI6ZJRa6TL8pL7FqTsND
HlJm5SPR/FNstxXZCdKEOoiR8YRjHELB5Sre3/ZWRboJKzXGyALwlDSzUOnm3y0nnu4KmESYHI7t
b3gyI3Texp6Nmo3X8LLyQh1mpajPgYkrXWztMywawCafbLHspDi0Wpj7CM/RN850VRsiL2AkA8tI
TUtC57bh7dJI19/a5abpW9WeR3oMRfnmKHFfwGSWvj/aIGxm7gp+nHN12f5slNQuh86Bfneszo3X
eWJz1vkSQYzv+PU0Uhd56HyIvp8ixCUCApIBkZX0eLF5mjBQxPc5Bnx28tdzk3kt3fAAwRB0QDgm
kHhbCaFxWMJ+GqGian4tV9LqYCk01Ptf4lvfIB6LbWLYFRKSD86PkOKEUMbeXjYtrXq9bxGTnAae
a9m1I33kJZfFPRNdtvy/dQ0hrSIjCwgY84H7Oxr16QjfVuTSUqUBUMc7N+rNweheG6zqCVWQd519
5tll5seYHsj/YSDUQU6xHlMEAPkqippV+7wVr9w5/IoJzqhirtMdcCfTEUWhC2SOcoQ6hQfNoS4p
vSxoEjZdvAW+4Tzqs3qLi+yxjCU6Y+hIR7qZWSDVIFkArz5eUfKxWcuOIoBmEwZz3rMYcSn+yq7O
flksk4CPQ98pPYjtH1DeakW0Kwy0OO4UAXktypRPYmy7edT9N8qYJUSC3c4ilNK37GrhOcnlU268
CsraipRgWbQVlCLxTAFS3NALWEc7PYZpKkH9T9bGDh9mZmFHFaM1qp4hWUaEDnXowHql9lwbKcVO
yw6alwooegd1YgU4Nq/L1q5+C3uuODpy7jLZAvAuK1x4WFKb3vqqrl0hS3MXZp2N+wYaSsAAN4O8
5LYEt8FrZOSJdLTR/PZfvhOID4U12jJd3IGwhqw2S7dOyQx9JIBdrgO7cv444Tfub2YBiLkekbsU
euJMppgG7sXb+9zAjkLNf9K5kTG7SKQ/ClPNSr0RMeJ8NCJkGc01gGF6SldwB5IY/p6QkOFBelHh
yXrCoGenAmOEAfldr+tcXaJrAPUgZomTqbibtJaBJ+s/sErQsm5ClUcKt625T2xTtswcJezAM+WJ
ccfJ4WGx6XgvRoTv19d5EKV/OyA4ZKvzCr/F7EWyQBuCZ5dQhf+teW69l2va6Jo89Q90sO3GO/6D
phb04Z+NmD+uCPbhJfgRa+oVdXGqQHrXhOVQA6IW5q7dK6ukiVc2cqMJvPUmzHP0G1riA+sWvBDg
IVf55af9yp1DtVEoUMzv7CcAipiZOMIlGibsKa9ovLndo1Y4zn5scF19nFt0iJW4Npl49GkyU35T
DE+1wU18t6d64/9XR2gqlbtWn+jv8ugKrEQO7QynxVs4Sc4cIySjmZEXhGVtp2258PDYKtVBvO0w
L1xEBWDioQ/2pdX/fVB3gxgivCTijMcDo5tsPu7lhtonNZ8N2ldOY6deAA3G10GdAme6gR984sOe
m/NsmkYt1rq0DEQ2v9++9UrfVxsQqqRKrcxaP352gsV0nmzWlDypwV5AIDOr0PWw+K9WZmeuuviF
ssH9B09+r7hMWCc5crew27ttQhm1uSVYRwuhxJJIvhtJqWW08rlJfjqGHoxm9UHxGir+uCWQzVgF
5qxKi2FAazl0outZPtoc+DKX9N6FzWLuIU+0QNGMPQWHQgC1xNoK5EBHV0nvsMLjlZzs0dk+CISe
sl6KDSgONW3Ih+/+cnPVq5wjcYRfAn5EMqs/GADIVaikJx/tjQJWWnKwz6N//CPbsRvtAaIuWhbU
xSqAKtTt9G86VGechr3ilyoxAWJsS5EGtZpX2ufQZDp6SvWhhXXggcLMsH0X1TiUHoRgZDxTo/LK
3Pl/2IBu03sGkR19oIePr04kwTaW2RmpW2z3nup55EZ+PKl0F+sOGfoLjCr7/yqZmhEfv45dihDq
skxXG69gAPU85cATMnyCaByW5hlJBFiC7K2cwjJKat5SqJUqP4TV7BnmwRv9u8YXC3XLFhy1sMTK
IYlMCm3WzTahNOsKX2tVihsYmzIlDY6kPvVHHYJAKAe0p9O1UNAcYbRPZzsgKBxwTb9zHMkhpuBE
KgCVqmpYdKk+VDBLGSIrcvU+EfsPfvefU1q7G1QP2tkfIi2jml6RWN45jDdTbBmBbx2fBpFf9HXD
LR/SU6k8SlBVqbxVHoxEnGNO3pGlgJFrz3Te/8Xmccw3fhCZRfWDx4S8UkDKeKbPjKaIgerrYHdM
pmZA+EKLlYOX1j2uBowAC7Uf5kxBX956ZMmcNJqee5U+liHrsaBJghigDYWFzGTEGOw4MqW1rojt
dJlIcDYrZsMf57vQs9Jzlgxb8lsrYv4reP4JhS720t0ffq/DGrmZUeCIyP/MeVb2SZZKLqdF26CT
737sQ2BiA46rTYO3F2Q0U//kTSuoCHCULoQyiFDH1khjF4NoyYa4VGjmKWiZ5aHtNj6QxMYUaEOp
uAtPa2Skrju1zah3l3SmjnDTTVBCWcstgRsqdlY8weRpbkjpbBggmK4lPAogQEOOaQIGxSRjJBvq
ToU4SZaLoP06N9bhwA7wYi1m/JOOHS/SeyGwD7O80bgZrkLT5/wnl53lZeQKqGeGOmllfDKAd7H6
x9vDdNA1CS1ZQi+spkfViS00E4j7ayV7LQcTz21kW2ZXj+rNAFKX7rNSdJGbhLJjeRHDrxYbz1mG
q06Bm7y2KZeQcGsiCbIG+cnLx8tByd03V7KQxeU1NyMlNad4pQ895bzU1Rp2fE2YL7Pfwl2SoJN8
Ik8ZR8CVHS6x+warlRRjP9BbGHqED0iGmI4inpg1F5TL88tyVJfzBZnHd00zsokDQIASmzqDV72B
qa/n5IM2y3XaVIEwj51v9TuM6z41EjanrP2g1fJlkPm8u0ZGCuyDN8iEuOAivw1z74RfQB1UWyMh
Uac8zuTUnPicLgufJvKBlk03UT1vWAV+ydN+8dtX76q5z5+AWvrbJi4U2qAguWCmnlyDBMd8g43c
n9ss2DsPmlU4XqizQuxOHcBtUKxWc0WzF5ln4tC4r8lh9DfZS8Dy3rLONDLSObnRB3v8QcBMAzIB
ggIMtpUWpHdP7Osy3K1gKbO6XO0sTqLyXKHwC2sZb7Mz/vAXN9h+jeSQyLebihSgfFj0J5n4wEYp
Bl51IroMJh2pLQXcSZvQK0/qw5abIYDXfwt81XugLshwWm1pHSQdhKN1FbyiV2CoUbmEpA7b0JqL
sWyAs6M9D8ZH30VT2fR8xHOTy8qIM6cLWmHwiSekRtfkswc8Vsp2+7YtMhSCNPN5r/FHO+6FDUfW
HWUwLyUn6Yf3riZHt0wuw+PDFOp8bQu6TkL6OiAH1a96O+FMcjKBjsirs4N2RlNkNYs70/fWPuEZ
Uh6Cf2KfpuKis+uNwh/X8bAP/zLdHbpChJ3kPDiwlvA2c8h7Mvhcu7iEaTIb7X60FQQ2JwC9ZZl3
Nz2ng3UN0MmkJ6+sWg3/hHhmElWxOzNCaMe01Sxln3zFxgIXfZQfjmEb5BzBkMiBdfe3X5cv8iul
uQxAysZBg+wxxPslGSJCJ7OldTYRMR6QHTVnZgAhFP9KsqCG8/O8/fDOQVPfhjpicJsaj6ej6w8V
Zew8ZxA1lD58Lt0jwcndfVuMr76lll7/+5IoA/gcJwQ0uxTeUHkFGRkAyMKT6TCbu65koK0Ku8Pe
f4hwCjBEQ0U48tlNg7ob8Oqar78aphdLcTpnBUTBXQtqx+wThQHJGbJsODhmGYNEcde/Cn2uEf5a
svm1XQxc80gtGYa0SjCckgmjMHVTi6UUS/xIrUK703aeATzTCYRX1nZgBDAtyPT6D7isOhVt4Ob5
5dJkbXiePpTMiHvtevjiLrUzWMH+HfHTBBmwIyz9J6ptosA9NYY1tEnt8xj+osYEYkOSlEIC6XSZ
r3h8ApiL8oIQKCTv3F9o2ewzNILnU6NnrjuE5ODUQRa7RnfqaY2i20ugvFXCGOYm8Qd700DSGPSA
j8w7VTssFYNQzhTBCtvvE7N2u5+vxuBwBYFxEO68XqbdnVj52NfqGeQtI7+UuSne34aKAE5Rz6pe
5Bj4FrTD/cIjGVpXW05XWbrCbru7LoFMsQh20INKYGsCrUu+nqHNShzi0t/7eEIVbwxNzRTw2Fxg
Qt/Y9OMFM/dkrpBrqYrMABUvf5PB8i0hNLKk/WHhsnoltKCJhXVeGlB2b+n2wLIdjhAVu8x5pW+T
g/rsrkLofQkoVlqSjcljTlSfsGR6U1/t78wA0fiZFnkggywV6vvUaqzHSehrx2ODC3U2IR510tCJ
fEU/jr6HXm8aAa8vi6BU1J4T5pdMo7d0yPS0zpfjWkBddSTof0Inqy7toNpWsMvSsdNtfYOLHALV
NFySHZg76WlP+OQ8uV+uUtkIa1myepIpUHaGc0E4m3BeJEnI4q+IjMv9j6Bf9zFW75ZjaI+6kc+B
l/psYxsNADKJ8JSw759G6JzpqbBlVkpE3Adn9LhFxuE2hEhz9KfS13zHbtlaHaDCx0+m/qhbq4xx
PfboBO9s0ZynWecbZqalE1UEngUIGPJcxKfl1+Q1VM4QoKEYsVufK7Pd8uS7zHVd72KQcjTzX3HY
CIY8adrov5BP/p/zlF65mGCi5HpGX3ghnGE0Wu6rE27CUyhTDNLQ2OcATCZKNq82ACTtPej4NYnM
vuM7KGeVIH/qy5sXkj+e1X3uQYR8EYtXLIceEDFx9KucPA3BpzI8CVZJ9TAO84CmAFRU2CYAMb7I
AL5MIasfWSEStBBUomQA68dz1TiMoXSVGDkCu0g5s93i1uLQRgmw5ncp3RMUXJm/36dhKHhGy0nj
YDNTeUaHxMZ69OgoQZkj2CVNZNyeuIznYkPLSxy2fAfwdk+x5I8F8vdapW4cRnKTCwBfx3x10vNh
KwG2uECDM5FQKTWbyZzkpEvIkXWizuKttIttGLkFMhwvceI05skIvQsQjiuXPo+xaENVAAu48vwd
4TpQPyDVjmDxZ/mnVNeYIO0n3aq+1XnSucM+mii9AaWZbNLCphcZpgkwQU62iok5982ZO88lucUR
V4VGmtOJwARmFqo2B5B3jd4V8rgeIO1lOPeE8qxJXuTY+ErhXdbk0N2lShpzWXNl4OzEp+HV0kba
UGYjemUsam70Mpar37cvDdPBftZz9YYfwpzpdycAn15aqAlXeYDnKphvLnnr1QSaY9Vho+KRWaLh
qKZ3bUGcfQxG5RU2zGhoW0f+sIm6vV5+RnlL9ATZK0sjtevleWfNQCeG+qBpgU05qDm5yhHBqIPC
70p5KRHHWyZzYB0rySYIBmGAgq2BvaeAVeYbkwQLHSiXf42dtXy/nYPfb8vG59Yf5bDYISRL7fhs
+sXUaY/9BaU3ZytRjVn/tvNddWbBnjeayqUZrPaPhmUM616O9IHJBTVEM7PO/w+nvJrh8yHSg/MV
qJTifgXIHZ6Ud3/gbMhR4dtlxL4TL6+7CVj64cZXzM/AmsDZ2QKgv6yqFTARYS8+C9AdN3+ueYn0
uzfY5YFXt8yqTrSxZmwIHTBefExGQnuAVbxPGaVux0QES1pmNmIiwELu4h11YdelAAN/AOx2oPxd
eULo+J0ap58H5OxqxjPctbCaXi/1zmSNpqPHVcbIgsij54KQ1DtW4wsovdy+c12zQ5vTQvblnySh
9EtuS4DzQ7tRIfuR3ewG+H3qgiXCG9eDVXywwDOZK07rhyAwZbKm6v1lDASojnvHFwYQ/+We45Y3
f1DMt4Urct7en7uk8BRQ8xvqGJTG02O2zefmukFhQNidlMMQMfaAV6es6sppHJZcDSuwuC+omo6u
aBO9VNlA8Yn9NfaUF871T1aX+M0KUqrm6WFrYY//dDyF6YJ7y3S5jkR883GPeA4yh2rlULhECNQr
AjSvlGyYUDGQnA951vGbv4L/rpKJ+eIXcb/ALvQFR3S+I8f5Q9hn0xRfAyRa9kqwuvo8qnrPOUUT
PAct9LQIjdlGsbycYQHRm8cFVychlbrvPdS8evNa8dQQtUehpOz5BqfWrLa+8i5D042lV7IUyKrf
HDa+Y1HXvculOJ9bK+V2XRTI5QhOnfR090cH1meiHaVtEfXaE/8N+rHIdzS8zQB/+ko62+czfLBE
TLNxvZN9LeCyNayXEVTwHC9Jm/p6jumN6foBDaUl9Hk0ZWyYZltvRHgFHrL3eGIOKkL0Iszp4uBp
cE9lJ1Hy/Wfo6PAFKW0dAMcauaqdk567UbZU1sjjcA7PFIQpEBGRX3xYwna6i7gssWhniY6DlzFH
U5Z+4L66ghLenAuKRLGsVtR0Ci8B7ywMFthjdM7CvUQMA3ajWeE/vfxsphiuQRw483jLXGvcUnAR
bL98gLuXpNfYq3oNGLBJJIFlC2VB4rjwimII+OEEgeY8UFjg8wGBZHh7SbqwSjm3A6EyIdk2mwa3
6bcdTQh2GyXn25C1VpgzU4zz2VHiF8tGWhIqdXLSFOa5yYtziJqJx8DhHtGfvvWn1tc8I0fsGq3a
pUDxf1v/cdXhWPYbpF2niyVmVu/xu/RXlzYnc6tM4r1G5qfg2XNQhNHufLnV+fS/gXDzJx1ZNVtm
DYmPiLCY5EOW0cg+c2/ekpbEyVTeJgWMTAWPYnVUifQicweQV6hQBii2p4s4oQkQe5ozhI23NfWH
a4aptN6S98qGi4xpyQZ1K834WSMiZCeuWbG4RTqpPYWCBd2WNdKojU6k0FDU/OR+E18+EYBz9Vbc
lU/OKROMded2vNvamRTvLJka/+ul+xOMdW4uj4g2QFFkoqaHTrtD1fgQW1p99WHf+vkShlfUvmmm
o90wHjcmcC4gdfad3w6yeJ8blMVwSgGQL/8wjBEEz6SWjBAmnj0JfcpKGFGkPAz4D+Q9im232tHO
06uGMPdIc3zckjZm89cqAqyAR3qv7mpfWPe506knEaBZ5iP+OOO5Ahh0h7y3TWVDUaz7m6ud0hAQ
rvg6xurC6SxiMgcQOaJbKig08l9J/lkZBppLf3a0Gz+4DcN8v9jYg5V/kQwhmy23pvmXw4R/pQcl
j6giZYn1mMgNVuYIRUecu3ic5QLltAatGJOqwZ97QasaXPail3JXqe4aIV/+BdiSg2pyNSaCB5zb
aAPMO9rHeMbq/yE1VUzAO4eK2D8T7wjaYt4zpcuRjjIm53nWJftZZNXhVUWXsjI5Wx7PraRKBqw4
RbvC2BgpNdv4QgfohF6VZqARZ9Og+gWwJflJX1C3HmtSRuQem2EfOyzw64CU0EWv2/mjc/wluJYo
CF4o0Y2Ldkow+lcFm+GTocFilvFeeqQWc17qNmOfQhq03P5QTGrvPuYHpLsFv91uCIYDR9V8xX9W
vAWA7C8ce5E8s8D7zSeh7MHmp5h89atgvj60qy8jPDmhYvHuAQTgMyWdOMo323Fwao7iVmyBTIiQ
TKElaJbP3tCeHLYsl7qrvYXoGd5ijDZVEzkP9n+Dl7lMMrE79OBhIvIxaZMmDtMLWV10CPl8rZEw
+jV8oh+TN/OsSBw1xRGLp6UexZMB6q71Tu5VYhDW2iHD7jpIZofTLFVM+EtO9iGBwRaXZo8n7m6p
8FocoUAunogDVSter4iAJkUYiVs5yXR2RJEBiKAW/vxRgUxamAQcpOmmf/TKi5Q6htn6ODvbZp79
Nnia/VjfHIHAb5jxnh7fEu5y+Yi/kM2jgorD/+rTZQpk0lbbvxncAduzjO7ua+EdsZWLoQEc2vr4
Si7rZ7MNFI3GKQUZYzUklDCQam6AybNbrm8G/pJUFwQ74pq7V2nKBSxpVK9IiO1eHRfKfw8r/Rzf
N4u35mguEEvTho/SOL8Vp6W9l+o7OwaSD1LUeOGuxaL3tDH3GVS+5As8mKAHko7LtRQL8HoI48Vt
dCtmrSP6Fsl9Pp7bthPkPzgQdzt3T21HSZ5O+HNzzvuiXR1RVZfGSljX5BT0BQ1Ga6i86pAi/v6X
QiGRwcXogl9PRL8NQuiSYEAub3JHigI/CcpBSQsiH2oRSTxyiucoglNzm/7MRR5dVbSJZpZ1+0+a
4T82pW1I6H2PD/s5ZPAL7Itda535zDls+5JgltNS1IhfOWtl56FoXhcI8Z7Rww4QQZx35fCrpL31
AWA1yA16NLaPnR7h6L3B3GbQ1BenXtUMuafUS8leSCu32oDe/GUdrakfgMQqS5FSE1Tsot96ld/q
X4qK38eKMus0eTqj7J1wQR/zSk4sB5O6L2BW1rrcmUr1fX/5inp5mHrrp5eb2qWcTklFZ4pYKeCZ
yOwW15EveGYSM/CQuxGe4M0hMpGWUFpuqpZculYBX56SjMKjiJPocL4b4NC2BIBd1cFZYlvqJC9+
63kNnsRY7W+6nXJ4uptHABqiAPaU/vmKj3vA97Y3d97i/2RbHpvSSQeg2T0SU8VOisUz6s9vfkPI
phaVVPUpiyhASjQeGKx2u2fIUokZU/QoF7LAViqBqIAYu9i5iWv39YDoZM9Vqa3kFjSS8rXf0TV3
dyR2ov2zQsU6y8zsjba8FgHl8TcXFHCxAtpbBEJSr4CaJ23MmGoBPb8l++5bCLWBYyrYYYJVFzp6
Ov0VRrk8PgtB5kF0M4ftf5bgVkhUzFn+GX5dYyLphzbYUAmIj5SvxU9bvrhhcupeZZP96nS2K2e0
wslhtJxwFAEDYcTc7B6Bfsa5M6Kv003pgu8SyFIF7z2PE9FhYiFnkYcCvW5/Qk3L8RYAX5OURjq7
34Nocf3iSdekwo7WMh76/NNZjDZSDrfzuhgG2v0P61VgjypkooO8PV90bzXh+pFh9FQbFtmsG1ag
CzWpW/EmiJ7opMfdAuCnLtROtj+N3LJkJMcoH1dS5cB5epnKZUhlU6/TrsPJ+FQoqbX+r7IqFrkY
wf/Q5K3eWNpmzs4mfeJJE1boVazbJJ1Cs0aSXMopB//tDtUiPQ/iOFugiZqGmzIy+qjLnS7A96Dc
XH91na4CvKuvM/ljfCfvXIPXFK2tTIXAWZqHg2lzn7gR2tbg623wmZCRoelLfDgeYdr1MPp5KHl7
ZjujwSOdQ/FIfwTtqMkEHzpDL15hp2Ttoiiit5Lfx2UBipQqqxXxE3i10kWZhA4dJdes676Flnf1
L7Y7Mf9jbIP2cvYiXkArAFT6JPdqPfbBJUZXme++cyhtoHVK0o4mO1UwoEwAuzEtUnk3aZBhO3rb
wTNd5k2rQv2L2t1f1sH+K3YAKj8WFhzg4AzmR6Q8f+QGGfavYC62kWRwO2YF7ybMqAaVxxUrHJTl
mr5x7HenLYSV5Yp4IYBoNpsrb8TGgXJThoFjY033H5TgIJNaKfA8scl7c3/L91WVDLTKH5nHk32G
sOpLNoiCCMjtXv6PxgN5OvzflDf/u29SAEwPdPPyohxxKXXncoAuth6kVqWJXik+l0uEmjuf1F67
w1nUu0bpApwOSp2gWPr0afDunSSp4ZUXNPFWEO42gw4Av6Y4XRTiwPJISURnZ25SforqQuS4GAoL
NVspEhRFvIvysS0S9OTiLED+opYz8Df2t/+wJ0WzJUkqaqKFQKQuM+5ZCf9s9B0zkH49gVf3YE09
fxurLzxEHHINud1ndSMKbVQ8jhDqUPJVx4azUuUS7U2kajvZfpy3jMFIwyGi+TWCeil/7j984+tv
vHI/VgqWl7c/BfN5AnBpf7YfR/1CkstiWnBCBVK6f/JgUBYdpQFuegE1dp7EsHTymT1CaimbIp4R
JeW4XUkC3VrfebOUu+q9peeempzJUAqeWVG4zrVGdFI92suSuSZWPW3TvzKRfLZ+Qaov8fFzNcRy
A/xOwQzRgfdPWGNG2MhQfpZc4V9zpLi2Sl6CI/4aZpZ+q4uODeBlyaZnDesfzyH4W70GbufTQ3Hn
URpa5biyjLjTYfT+m6PFjiZZcjFc0J5Qje39IgoDe7sbHAnyN+ycY7gY2RBaeI0EPTrnrjYRX7SJ
XBP1ErZ56d2q3RXNPOqzvma9UdecLcBHxPwy6dcsB8VDx91Wj8Na3uc4lR2oSyGF1wChCvo2f3Sl
TZmc/0p5snJnYkWhkCt02Lz+3P+mHfnqFJ1cxbpoRinlsvN5I3EGCpxHQwKoZd01UHYLytZ94dOm
mSICvD+7lfAjVf9YUasoYyeOvX1WgjXWZc3VPVACpIBDU33dnwFVtUNn7mjfir3AkMyG52FvjgP7
KBA7QYNU9dxXAtTGcRPiGUtb6WL1zbXys6eX5CvSJNTCY4yCPPSQ1vAHj3ymIvebuaDYZcrPeCL/
UAHRN9G0MNZQy1JptJIAuEqhHiIaaMzo3+PoXXndR4ezIffXSlQjNmg5Lx3PlfFvK8VGxyFDvOxk
RtdD3+fX63ZqdUbHifclu0Khs+pDwKnmDGiFTR7qszeKNPhQnp10KTPgxKjTSSFpdeS2BGVK9V5e
hRRDDP1Mq+osus7OLrdxQSg7VCKN1Gyul0sKgar3guU4Lje1v75qKC5GTI5Jin3yPbvG7XPD6la5
d6SuTamk6kUAX1jIy8DUWw2JJXq3bX/yOjusvhlYXCWnJkOlmudg2pHTa4DGlwjPHEniuu+x6EGG
LgEyFqQ4UdNDcFtr5VXO1VV+dzfw0vVxYG5YDovRe6CiGozTrLwWsDth+SAgjZO0W7ZNVHNaSIEr
ZR8LgCmnDouy6VXq9m4f+cOiBuc6qvMmfjX+KA1llvzjcow4nB81Zv5MD4+k5zGZBLVsSoeTw5+h
fb5QLHnLJ7n0wEQzBvb8YlYR1znWbZKBPX0zmHEFPwC+QPJEhZpCyPPoa4kOpRLCva1IICKrueB8
r6EDw65EEQkGxY2kM8/o5zGYSQUN/KwNZOTPA757uAILz50LvHLl4qg41kkY6Ilt3Y25AY6lzVdp
36lFX3KDVyrqzHI3NGckaL/k9QhKJoO/KLSgRboQgvP9vVHnbWyB7a4nTkZvTEYz7a+MNJPDQ9nJ
cYDOO78Qm09klWfsmFuUkUEacZ4dPcUwGB30qNop5VqT+24FX1O0QbdXTtOrhoevh+YLTnIJsVUy
Y4bPg4f5yU7UupnGmWh7/GeCq6/yx1cv04bUxymwlwAVhUemHFT/eyrOSWpEC6TMPdfzEgAQPM7A
L7tYXZ0HYCe8vE8k61nQGJBr+TmbeyNlEdgQ6pUR2yr0RcOVs5V6iB+p9JqiUcc690kNVGshmH+F
LYICvkDz9GYemNUKnCpERbZlGbUIb8ieIqWHcv+scVKx5LHIR8bHNVEoaCSvHo7nmlkZlsnJ2G/X
RuIzZEKvvfWtrc9N7MR+rSCuxOHd6zN2b/4e1nUxFZTKLy7c8JJ39nLEB2q5fvjjYwVjAbKLOYwv
x+S0NmZ+yGzVKOSUMFbEo2+qGcj5kHvs5aZ6KqyLaKImosSsNH1prcZruQ+EDLVEy6YWm2jwFmXp
1JujTApxYbk1uoAYL9nkY6xbnKRsudIJZnU/YsDpMhvOhkL6XK6MWk//BlutJBUj4MjNRLJuWRhb
0e07m8+k9Sutwl6OEPB/sHoTfak1QcT5BTYN91rtQIjSbGqSQAs7o08YU1cszEjFVpHVaMecxNiT
inx7MaCs/JY+ciAjeE9aXKDgqfX1A0+KVePtJ/Vtkqja50uXbTEcTCH880ASTl2rmRzZvpVHMmt8
a6SKdnL2f1FFgrxx0yTCjeZ3cOEjzXLabZVq0HEYOrdoHULvV3zVg/KK5t6tGDRT5zgVjkSPnJHn
6z1oRN9PbKd3L43lvPxkFxGO+6yXtOKwwPVSM0Tyy7CpESjjym/QA/9b9dJD6S9nNFz3VaFLCUpt
hf5yJNmDt3sXY5M7vkClDZf4pymDqT1Ag9r7olxdh6utXGabuNu2Zd9ZDxB5P0s88mzWfhdbZbtS
OVIlk0/Wv0Y0469AjWygKC9xW4ySZhJwTbVaujCfRhK9neb4QLHUNMd4UVTRKGDZrxXtAe8SUDSK
T4zmZVKcjQvjuQwGt/oQqDaFBR/TEZMLJJTwmVz1tLotnmHyOH80Q5xql4V9RVBdUk8uHx/Dr5S4
QY3krDbK+Ie3SdgyfGAJcpQQbQaWGHVfRs0EQ3aQUdRRbHSoMrwetcsOh3PynyxJmlemQakNobHi
TRuTqPvKlhgZ7XD13HyIaHeGxhL3frPVwmXD1nQzghIp4NQza1rYHjwqBvgF65zNkUUwsBq9HW4q
vxI6MAwGX3Rn8KXJ9wUcSNKH9GNBVRacJLH6NVE+r7V5yT3vHjxlPMN2Fov5Bv7uO3xq778H/4JG
9Ic3SIkLXVHEqiNVnUBx1lmqOj0QlUcvGRjxI+WizS066lnUDxlJzysfWC6ffrRA0oGy38wsHf6b
lT2EpmSNhEoIq+LnEb3+Q3r2VZ+Ox9XXIM2/RnFt5lB4wrP8BFlvNjmcMWnFwbZpMsWkFW10VkLv
qwCjnnKzcgV/3Q33sF3N2UPP0ICwyAPA/emIU+Dx9nEf92mdB+/iPt5OjBT8AYb9lOBzSJSM6pXL
AtlyBoSsjIjTC7ue0h5Y4MYSMmOkDlroWQO0Lh7t242GG1g/Z/s7wzWyAbMkpgvbK4zTc8Dktcu6
xM99PXl48V4ee1bzyS6amBV6xScZEjza2YmtIVR+TBCjD2Xsar6lCS1N5sU7E100eoXarALF3QIa
UejDEmACYYs3UMXUpEbqTsq9w9DnfrPh2ohssKWa5Zx8sshabSmoXB8eTULafKj5p7UTW45XQx0p
j7CqlrP7tAbut5a79CWnJs+0PTjgTjagId5CCPK2Ul+a/Ibn32ysTAlsq5rQzBjq5RKpp4STrCeD
+X0sMaULGKesmX+kNxUGupo19P+ALBsay796Sl/IKD7MIc4iUj2sKEjDhV9ThDNHTcb1qj+Fz2QW
V/wHqy9BfYm3xtff8dWQZ2f3pJWVIWJvYaTxvhxcY3WqoFyIIxLMyyV86g/k7u34YM8nphjU6JXd
N54zOroxFemybafu7g/B5EpKJPUhAj4RajePtx+wNpOZXsBv+EOjCEK135yWAd4LWT6HJU8X0A3t
Hw1KPo3YarB+bJTJkW2th4LKGbpRH0fK1uhGWfPAzjE3kimVtxjjSXSq0g1HHC5gU4xL+8KVs1ix
xFZoWeFqDC8CVCJviC/WidCdIWwVVUd7TEOM9KaZ8sZTgxRtguqIlBm3anZ1mMSbQh3y2U9+Z8hQ
WWv3or29o6Hh/hpfnxajtoBrWTbMK03Wy1novbkYcOFaBDdslnGpXjt+BAQjLdvlLchJuTAy52CO
A1ZvfVlMv2WB7VBWARIhfTc6c17DqFFGsQSA8MEURSo2J1omwqp/bIwIWE7DNSjXgP1p42K0hyjt
L85rVQ3ij78+shsKHFDLY4lY4Kyo4ZzllkZ8hJ18MKQcAYXXF2U5tgv+71S578mhP7frLP5CxjHr
hw4wLbSHJgoru5xNgH1FRS483l4duGVwFQW1tpN30+hj0BHKomfat8XWTBOWeXOeVKNgN5cyQEQk
qvse4FDNcCp0ra3M/CfuvUQI25RGeKSyhVnSyxCHUbDBQ+pc64aRTg4/3JTZiXLnbvXKlxjwfF24
NEBLMQsuv6xDrjFOjSlRK1i75mk8yFIdlkBhQxtSdvRBrPyk0iZfVFEjxd04JlibEV1YFAbejvTB
ijXkjNgFx+SNYxQ26Vx2Lb1indwtSZ7cfiYPf1xFqs5Vrqpi13F/SFrP8No4CZnDpnhHAlwf6XOC
DolbAedsS2Snot3xAgmeVb88aQ39RS2y3MiBaQs/rAyCTNZGBVlGmwH59rGLU3Qc9Cdj5MfoL6Ix
ayxBy8rqaOV3p0xwj2JeT16oD+466bW6JiZGYgPowfxlLngwyjfrK2pAInOZWm9rV/Q04Vrygau1
m5Rd0fIilvK0of3QWODfWVnGc0RV1WjPJKtdaEy4gsg6PybYsIVEmbqQNZvX59aS9XNI86eShQYz
bzE46Q1kKhh+mlb0jlN+Alz0fbeBQdlsvmKqhL6CFzU6AF29WoXjQlVIacgGMnowB2r5q7E0EmY0
da7etgj44MGCKENK/Ktz9R/+CPk5X4Qn7LA1dWqTDqTJxx3lOm+TwxzISB5P93VBFI226m1nID1c
FudU8o+3wSWd6epAaxTPFrFLXnsxnwdwFvzvwrhwp8rn5Y2wCwk5Xy0+3NftG7xP6upKUwMqc4lq
HmcDuOw+NkVuAGOLeUMxBEtSLRx+jUuOiop0y8YuCL/hmwOHkdZ/MG05cxRjifaP9KfAzNTXajNQ
Q78mhWC/YjxkzEOrIVz0usmVORqrS0OS/r+VtV98n6vygQvTp+by07ATMsf0eCxif+bFBfL5wVg4
IBTGly6jt//if+sQjD9UsjwwaUCeIwGf41a//bVAWvByCRUwMO+/SW7q1qXifImvE/dYvWtf8Pqx
FPBqRENnrMALAM+iKigpOe2OwAo9w5apDZiN62cDmPA7FbVeZZYDEGtOra8ApFKfeJ79bM8aWYdK
LnKy6WgYyNeXTTeZJnucl1d3PFzVztkzPARYyr6AFIq6AGzfLrUQx67ocup3G9yvl9bJqxPGZUNg
9SMkiaZZwh5vFfU1m6vGHvp7jPUVOlMtd5D2Ri37IY/jVJOHYvRz2nka02HMMgBKw/8xtm9/kswa
FubY6c61mzdVblfH5/Wwau4YAVauvECG40omfBg1AcneV+TfV2Wf7tzeoDiVObLQY/SE6fkqBCPS
QHf2lQVZF8XzVzTFHKwKoXlge+QQn4fX9HQ/HDsikE7ivBInrv90niraEauysRvE09FUCYwvzk6z
P9B7UBbt33K4i8vV9SMVu5y/LwkgEezGAvMm05IBpNYRw3nwmG7ieEyNyoz9lISmgXS6anLnnfH4
9nw5hyZ7DIwB8ThQhfZCmVZI/Ndxkan0z5aZMFiZSQFLMYZvLn+DVB74LStt4OTo+MNZWrtBQSWo
2worYJPOhslsUkC4yXvRE+3Tx0jZ6wwJdy3vmh2qLj58b/+dj8erPOP4m98c/+GQ5jqSrhnuUYNt
zpiE9rHYJi8UDvPbXCHdRvFzp55BfMc6fItDdVKp9jmYzVec+R/joPgE2uWt4ka41/QFRPNx9wOc
VPhkJEMN4pW54o36T0nUoobj0J4u+gfMjzzO6ExBAm/xpFa/upcxaQdhQarNSZeTP5UCInEFBEMH
MnFeTOeMnQ1vDLm8qxLHicMRWS7iw+pbGXB6jGB65Y4gmuacHEyYzmxuGQNgDktBseZYI7S1DOv8
+NATPbqpnEWU1VgqfJSyMuDwKqV9bQO3xm7U1Xunhxo8KbmHS725Ifb66hsNEIrFAhf4J7XTw7Ps
/oRAEoz2qxyObKvzLiwLKJGutg3tUlsf18HMUpl0UakpVwygODaZUs75WdmoCj8Joiz1FFA+w6Sf
HsfydYYxzNhCHV20D6F+aafM9DKk3PK1298IR3kCTsSiJN0gURAbFGCYlZBN8zVstXSjosScrAIb
Jyf+TS9QLzHzaoMiww6ZJTTwhggVqjh2lCWdlS78AJid1aPOVLl21E+aHRDY/khQF4zC7FA5CjEA
g7S+vesnuqpzBlrf+YlrW6b6OcC3h93xM7U4oi1Y75D3cD7v2JQd3UpfYSbMJN11u2iWhIsiaehU
3eRTC2uJYp5Ryxi+MGqDRbfEoc0Wno/fJxS9OCurbuosU06xrfHb25ZxJqKlhRCRcHqADMlH4bbI
Bw07oHCB32Nik1UHr4mSlh3FYt9aBiRJW8Nn4S4IeCMQwbQTtJUEcQwfHExxR+iMcRXStcaNSRmp
sHk32fpeSn+mbqO+vfXD2qVlW0xUU4T366gAw40dlsmBPFfZDDZrHB5wcw0yukb1zoQaV9ZCi0J1
tmD7KhOOSCnvqdO7CykrKOq0PsaPWI5sBtFN4nXmWFK2pOWBjC3YtNj/g9TLdUtATp8Gu9aKQ/ks
as4vynZo5pFfgifeZox7Aajh6P6wudMQeQ67U79gKoXdEHmD4ZXOYhlX4IVx3FUVCKCy2zskhsy4
9v9Z2RMPlAAxWG57yn3zeM7iX8Z76Im2QrjpBLFybKjsdkL0i77S0VWvjCGwEFdDNjoMZ4+APMbL
Eytt9UpTy1tbvJ3PF1+fiRlrqbdw8Gz/42ngqf/AhWJVIn9UR9bRwzrQvYR8cQulAnP+ieKVTXTO
QDBSGZdBkBWeLyrpIpFrwZLzNM36Lzi8sjmQLrI2SDSheNbAAnwonKTFNCH+UHN2TAFdVPKSE2eH
It2GAZprGkQXdLN5rq0htAWOFzmZVRvptOj9tzPQsE71K/zId3RZgKDJG/qnSCmzIjvsa2Yl9Iu1
TM03OebulOCneCR4iYpothQDSnUHE44BuY2pRzt7pHO6F9qI8edYdy7uvgO8xpfpY2yPkvjMhFHn
UtmRmaDiSHpf1Vfz+7huSXGd7xdq0vaYte6DXXmtUFvAD8jQIvW1GSt7d4jt6Ke7oLUloSy6O7mm
LwezzZI0n+Q8rCCZBSagsxgaLDi9SEuHacoe2Om9D2cU92fjczd1Yg2EGjAYPhbqFU8jTp3Xq5Gh
aQfrflm1NJivDmLvGc1M3KcoTatYV39jN8eDw6gcWRecze5EYHuGOhS6uazImM/UctIJF+pnuTSj
bNv81dR0DSWF5Fsi+s0/MYIR3tvr8+s+dyFYreAnr+Mo+TR7gAaVxMe/cgMtGY4edC5i0eYQwFJs
Etw86P179yQx4g8Juhz+exkAqXG2lcJxsgAxWoGbnjEC5D1BCDf4KNKhPD1kApbNPZ0UywERNubn
bz9HT0+G3vrIxKZB3Jyo5InGbd4quk/F7Q2TZSin53t139PXVTSH9oBvKbc6uAzij1IpX/+Yfm5J
IUnRp1mtUkw5SX1I5KQW+a9qUTq/9IW/l+mqIbWA5z/j4K0fdGsSnHaaLTib8ozDc68azBaon9B1
9mw76jB2hHnPF+4nFSYyX43BweEwYeh+bVB3HyLp0BMiizuIO2CjeNHhVn/GIurSSw1I48rP2ZU4
vaYZfEhXqGrwXQ+/aFeBafORfl6q4d6PLLpGfvvTtHFjrbC5CpG1Lvsv7Ch7olkugZZw2ejcjplw
Z2j5Cl0lUp+t5xJZfC4260f4z6zM9sFBzWTlEjVXDis/xa+Nb5qDmjNpp7XGU3d67VrcNhO5zlWY
VjYJnmZmwmDx7MXfAClhVT++vFfYkJPE/kDDKCbV8+jaFDU6b+xjTER8w/YgqWgPnHRXlWbzp4zA
DIzZ/+T8a1SdO82Cz0dkWAeJZ8kQ3MlAlTJ3eQgwl8wYgrDvasGc1WJSEoseAEojJKBG5I7CPUpi
sjxFrP7Pg1TIamJesjgclA3S9VPtDofj+r4FcruXVCmX43M1hXGt7JRIT5LE3dxOArd4DL+9spcU
32lib+BFC38uD7l024OG7CEhBexIqEY119ClVRZU0KnDcTZfwEVEdDELZUHeAMu9PaO2tTzTUjO9
ADedDUhM9hGCXAI/6HoVJObmK8bpvwSTKnsa5qobMUMPoEHaEneMtA6OFsK6HSq8issDsjWh7hDg
P4UaPt2vtzSCvm6VKzLYEz6ZZIKU6fES/qhfqX/FrO6dr4nXyd+pQajQc/G/10c/ga0RK9WOdbpm
mz30f8n2iQjuT/jQ49NT6nwKz2kTg0pX/fvmWOrFUwaCxKE2Rf85Ex0Lo3pNNmDDwWiKF3NOQsBM
7HmwbYpYWyUSQDemAjJ59s91C5BQ6r62oKDhH++Sz1t7disMTUAm1o4KI0b7fptnbgFkBtCot+A4
gGVTnLLTW+j+eDwr+iZFq9umZiMQ1yUSBR49jkS7w3q8eBVkvQko5K81yzkTstH1ooViWnLwwiSQ
nPzLq/iNVEWNr5xgUtni+sXrtxw/qcdbOzuJXrX+oNmVylqNvkBv7p8pWicKtRGs6otYFkgusDVM
XrIWaOreMWaI+hL29CKYdswKQ3aDDIAY+x2umspeRSOVk8vtYaAfdsdDl1UpEqGw+KeI5BGHUKYt
CMSBApR8W3SIzxqxiqnysWHNMbQQ8tdLujQOzVKe1GUO2IDplTnd3q5MyzPcpL2W0B7qnfkeLzrN
fOnVzgOnmUrDupkvNq3xKSW7GTzRUaxUxW9+u7Qp5DS7NyzLOoPZDaHzOu7IefDEmAZrvyXIvwL6
7ed0HVZdE7h9Q4x+MwOp+KdwoUQ4Fs7+JTfSGq1joZFaVkmXkjJrdCliinw8yzfXw5grIqfMl1qD
jTsFVD8Tp2Kl75F/2Bgy/gxU2rHaRJD8ga3BUIb244QA2S86AkAwqidk7uN1UofteYEn4ay2Wd86
4BjqpZgybE8H0bOLVyifDwNXWyECxBrQpFJuTjCnf3g82RVBkz+Cb94HWYdjr7x0E4+9F2XWFhbN
VCq13TTxyp6mmkvSVo4GusOXxP8zpMy/jQNFSzu0Bo6BKYZWsrtf+Pbep8nBR00IYjw5KXJ2SsjA
+Q0fHm13JzZhSBp0g2xY7vPs4fDlIVgUpBiT6aA0PT5dACFaqQ6uiKWG0DN6Qr7fzIYO/eVZ0Jdf
eDMS6JjQHqkPL71QZdYVc/D+2khYi6lKYNai5r7baHamurd7zYOCpo0qQc62em91s6PF1k1P+n7I
BObSOkaZ22r1K+g0Lid7Oc9ZfcVqPMCel8f8eHNhT7wydHPUVxckhjA29YmElQ6GWqYFa47IeArh
AwQ2h2QAcVAPf3xBEvJqzcKOWzzZ8lC0xrgH5JW/uibtwgSaN+j9GRehoZ/XUwYjFGC2ZXFek3St
ItWrLrbqskxsTXRQcXO+GDz6Uj/Nnr8CrE7WKREY5AcedVl8ODfP2SH9v2sxiIXpUIUkrvYqhSWv
6czT1ExnVmpcBWP34Im11sX6PrjVTv4nOcXAqfzkesMhYBmIwOMYS50IiweeLWm0htQkA1hbeb5c
PI8NRmWldYlMiRrAEfpefreBFa5W1DMlYCMuTpDEe7EZBbb6BSR1Zpuh1GzqnR7E1vcstnggVyyv
/f7kdQp5YX2GJPqQxIUIFE+u2YxbGGYzMgeYnaZyi6uAjkXijgmeMFgNhR8zU7ejSG3h/RAOWYVP
FPVmOPTbmroexcn5LGoXO/2bQ3qSsVrow7q6R0XULJ0axRfJNkfTI+h9lZZfoi9thTDzDDmYh0IB
C0l/xU/4VA3Dcjq1SjM4kXmiv/OX3Uyqo+v44I3chZuuXY15F9YXyfF6jpAj+z6Jg4N4FvwMh3y0
YLtdWfwZx3CRo3lap4VQmeozA1IFUQhNI4r9eYrStJ0PPSvR42ifnPyCyTojh1NdA947dRd7/3wZ
PN1WtqpY7jNVhJ+Vm5/7BASUp41hUw83UsnNtc7BzJ6Pe30WE7ocmlCVPsHEtNNVRwQgAVLituiI
bQIo/4937KStl2zuUHudsi0uFmIKB6SCdovYlUj0wMBKw9frCGxBPI7FtxHOHLJZ5wiS+wR5+naf
W1LG6jMEzl+dQG5g+kL9fhCNkowLqbYTnIf8LAJDrj5IkQozB1Rbzzga2NpINtuHVd9D1e/0Vkl6
f7M2UcseT/H8vz9Q34XfbbXZC3S/7SZ6VkSG9fTjT+C1IKYY46MzVWq/gU1iwt5JUz4C54QZrioy
YsInpFCTa4/CZW781qYVoOTwHPt483ovt8lPk5SfOsB021L5ZwBY5NbYDVr0N6S3+KMazAKm0Ggz
sLbfOnK4SRHhYLPzRcgoCVMrOfqUSU/S5P1Evtptp01A+urCxg2QSuNHf3wyGNmBkU1VLLraT387
mQxx8UWzDc1gKjhF/h6GgxdPAn+Knagp1+1CYQFvcWe2V2VusdH6n3os8qKRcotD/vl/hxdNiBAA
fMnNBx45+SmHmagwtctkF14yz55rYD0jbb69JZk7wQTN3I6emCipmDt3jfuqbFV0+ZqQbNQPoLq/
OR31N91QEjqyfufdXND/AoExqLftF2Lg77AXvw998RFN/n22LcSv0eYlbnvT+MwgN464KQpkEFCu
WzzHYfGGwHRCbkvEWsfB4+XKy81f5D7bGYlKUU/8aBsVRVAp3quFUVmw+ESUBZwjAvn2bIGMa2Uf
UvmaBMMpTfokA5OvuID1GlHqNK8ka83B2TULZdFVBtZh/zmt1yxkzD83ftECmA1pXzbjUkr8Iugj
ib5ckdt1CPr9oonsi2tFXh4neF4oIA/pgB0e635ER9vHHXqn44D7FHUjXbcI/wE5Fv4jdaPvFc2Z
2qKosJWFglLFXIJeOmG6M0frbTKqn98dljSoL4xrVlGaLWXJvsxDCSevVZsNyi322VSqcXnLNvbm
Fmq59dg9rWCHFigwW9tGBz+/IYNkoJ31qYtKjfIDylGWh40COeIw3yMxIwEcCki0A4GLj2CsDxQi
Utz17YYc8pXPi0tC6yiRyTo/ArxbkzBAoIAV30pXRfuMq4JKdq0rH8JShSJOIR12UF10yeI7aCL3
IZTW/XkvZVNqGeyhmKoWBMzS9fwQvdo9iPqBU1SK+VBRRe+uCnxXaF6gRXSUu4Yyxuh0C4Unfsdj
GUdwBBaGYgdued6czj8/iecrUSYipHzLOd2Lo6/Hvf0cGXVIrqiRcEWqGOcNUQndCsgBVHCtVggn
LgkA+E1ZAGfGwPihJ6JAo+bXrqLq8gHmavhqtQQesQ0qMzA9EH178aurvWWJ+G1hoUqz+P0KCZrt
yJXcNlD0ElsG8DFi+k0Id06o9rmntdL8Sd2TwK1NIffNFEtL3fzgwUHgC3vOyWHda0ndd63hFFrZ
3ZXB48ujeCBBssmuQDpF1MPRpbRyZwabnrnxbi9G0HFfANH5AHXlHwjuLUaXhgNtp0zgGSmeFxkw
SHqn1mbsDs0Zxe4Lg22+Eqq+QX8OE/hquEqWjbKnPGvGiQa84qI0Ib5cSK+EnQlQuGNeV/Sncip6
gyN9c3b3OWAHkGBGh7M0dE1vhFsKH1k2wGlluYXIsPRVURy/MgMUIcF7fn719Gw9qV9CEpxHGNnz
tChsWyRjj64WM7WmbiytUcfaB1PG2HQchfpV0MewnrqD9ahNuNp6DsCxi7Ii1R9G288SOv7V7LOT
MlJljFRbxOayxnKGh/jxw7cNY7RWQOL0vgmfJ830bKJ7o5zKvBfS92a5BJa2PHRLL0ZfGZut+mDt
84KzGQ369A1q1KU1SFERPDgkzJiVqQ4Qm7aw6I6m5czteUwPkKvkBchNpEXPrQmgS9qG9cexeH2K
nWJYfMynigfeqe7IyV+cl0OgTYomWir2f8bw8SuGwkjMfTprWCU65Q1ON9gR7OmGYpKgsO2P9xOr
T0/UXjYUaJi8iyzK1/GKQ/wTj+sF/FVhDWtHjWRKeAYXEX11+v+Ua9KrswEJh9p8IFKs0QeshHf+
QAYq03oK5BpwTy2r5Ctefba7ThkwVWWib8QYdHLLZ4rl+LTR537UHARJ8DS6N4+1frw8hp50qaUa
0GeB21/3Tt4ES8BVJd3TG3M6+AHVuBRXDL4kZWF+2falJfNcAIhh+OVfu3nnXYHe1qD0OuM5NYlU
M6DByMwDKCi3s401Sn181oR3YCgfPB1IxF6Y9sce0BhtyJbtIBgdKQnUietlZt4tJ9a8q/YKypCv
aSiZwQASouwYr7zeOGe6qFIeHYHxmvY3EonJJQk0mGQho5XPy1pWGM5r+WXew13o1uB3QVKUwLcZ
rNf7AlckrH+DP9vH+9i6Kf+QTYEXChRvQgLrSJNlKJKrRCDwPiS18kndc6YkA9jq0UP/WP92mbWy
VSGSMoNuEZP9nWMETgO628jDPJmhIZMs8QNdPWulx4AA/PWDAk401j595GUnQMRyfr4E1c6FXRmT
fvihqq/5U9VlmPLqL6tBB0aOJezadaaA3l1rfz4MY+gQKaioqOswXMV+VSJCrdYqUo/02G/Di0IP
TGdAi9Msgs8O53eQW8tdBgRR9+31tccScNyyHkDvzjo/OJEIkYa3DHB3ANvPT/PzHaol+RAHJ6/V
x2FLdZhuN8kUSjpuiHsFXpLTWMK7A83nHh9sTKH4V1ukvzEtGF/Y7zE926xn9fFTOurK1ADpMJW9
thXDLwkbsQ3uCEJihXOGkmlfAJcC6inYlfVllSWAVrpdJZfJZ4a2zABFi0r7+PDzAIYqY/x5/6/X
HiIKJmcWDfZlRw/KCP6Jo92COZ+sGMiIBb3i6I+C/Df/c7KKc2BgI0d63fQor2v1DfzUaNPEXP8z
CFpwuAI0q0S4Iq1zKwG/ZisXnIpqYDV11l48DQoW+f0j9iRYB++ZMnsGZEIwyDydWgPSiaSDJsEl
IPtVNeSUqwCpqBBTQXtGgZS/pHqT6eHfMxygb3sPSi4wKsSdopwP9h9m2i+LO520Jlw4RgC8d/UK
JFSrZUQDnCnYSG7jhoGRzK6DGEMY2S6ZUTAV+mGP+C9pOw9Q9VOHaDpapmj2I77XX37zk/2uj0YM
Fc+GBd+cUeNitNCiHjTYCrMllZmRV64KGZ0jWXoB/7xNRo0mgHyKzN8Q98gqXBExHS5jdWwwBkPr
fgaB1DNWz4RXjPjIvqAw2tKm6AiWwTfZdMS6i1i8FFhlOTIdVUqvIrbgPIi6CYNfF+f7AyKp5knv
E2Eqy27rQ7QxzBjtQzrubU7Rjr5PEGKiCuUDnVstoxXfoJGf0oYpIQ1tn+auJygANo7I+Nr5SY3p
o/d+Sjswv1pkZfWWbFN3gQidlLpiR/5Wd0GWC5ajRtKdbKy5mq6VuVcATFG5uDTwXRwh/bzZhgLz
xZqRSftPwjM/R5M6RFyhgkj7MpVBmO8ARbuck1/AfN/dKcIf7DGzas2nOThX0QAacG3TLbUz7jKM
uaZSIWaWNwR66ks33cGrZefBEd6htbUYXNWKL39FPhJQA3PFaxbBZOpinfCsJZmyAM66btyBFOsf
hyq1ThoOYsd+sd/mWGq8Oyt7oAey7ifa8xK3uLLojHEb7VlZtCo6P3wOETDJW0MXZSheIcj2byaj
H5A0TisyUB8GN55ymTeE8cYaLfdMNldhMalHjF7PS5LXQDZzEmjaO3ZYFmZy7zy5Qo+30H87fjJB
nl++BKuue0iu4DaFsG654I2ROJOwDPMsDLWHdDkSY8gPTQFu5rZ3DUVXCVbT3YqrJkRiUlk8fZ7/
nKt+Puz7+q/OScEHTJ+EAJ0EtJzz3yGMhTYpJs59OIJdE76kOcS+naPahl+BzgHAYd40EH45X+2K
dKsyR63nGqwq9/XW7I24a2U/xSBydNbX20FHBccVS2j0ktd4IftiP9OjyV2dbvu+24TwmgKjghXB
RpORs/MPhHZ5CUyxf3lq0QM+r+sNux/odTazlGzp1bwCD7RdmhYyKWeyH3HZos+vQIOyfQZ2tVbK
FMJCr7IiU+eEgoiBuHoVjidV3xMboDoT9LnO2S3rXPisC1quwO0v7iJizMiTcrz6obr8N0iPtINq
QuoHWrJE3AMlt5P/IeTjaMvJtRAr/zz5qhnzNl+YMQXlQHP8gNqdrflZDG278SJImPDU5J2pvZUW
BW6ZQqRF9xn3BgGTD7LIld/ijPAX9XJmUDzmKIOQHH1vspJof6WiYuWPFA07IpG3V688iJCVtesW
PYRZHXtDM1OcipuvatIju+G/GWeceLj52KTyuwwM/KEYnfjx4LZrCfQf60ZOnF0TnsPfk+1t207Z
5GPSTCr6VVbEOcWH7Sya4W2XJxKu/5wdvZp0ngxv2p19IBXaUA+hgmbFTJIv7/pISL/qgp3hTe4x
isCn6QeJZJ+ZvJbgrqwQtc+AME5t/thE01JzAD6eQEHdjJtnA/xWPv7qtvhIoqT5lURSEouqzbox
zFbXQzHMznth9jDnxL6Y5wFpWWxT9aXVocaMAJlRp5VXYZJPXdcuUQDmoPm4B+22JgGreNOdy5fL
yvRHbNNZRfcO/R76WVjSJGkv7NYM+KnFLltQu0rIeSltMnQTr0Z8CjEYWxpUjIYeZigdLeZdUCVf
7X12CqWmNPAzsPveTS3FtLK9U8h54PBh+rw9LkGfie+pINAX/FLtiAZdyEi5m36fCoXaOrZR296P
jUM5xeHppiGHws7A1tnzFIQJ9xqla1DUSeVFBbcXGeGG1T+GaUiPWu2RZYnDf/STMFIjvWwLhGe4
XFKayNWpijRDiVeCX/D95UzJKAAd76MZUm6j40/vKPx3R96o+b7HCJ9hahzE2+wjRTfxDmel5KYc
9c8HmIkWYavdUa9tC254kJyPPu0FywLxQ2k1C3h2iGLgk6A3aDqDoXUD9c1LSMPk0N1RpLB3rAbC
FG5iMoMKztYZjp4zTeQThwaL4rJ8dXDgD6l6SHRX++aUMVcd5pgH6vtTTeFTF0RVuA9cLabDirKU
PL86NbQYb1YmBtKe7CmMZkT108csmeGTnRS+xC7yXu3ZEWm76EogwVruWbX40qw4wudQCuiz/512
CQBrOT/Exp+H3Rt/fyZfEH8y5OVsARwMoynhB/KoorzKej3hOoFWzCYdZWxzdoyf9MzzwAKoVTj7
RgEfWu+JsFf8PpeAU1ZmlB58JTnP3eX9OR4HoZoejAJ0sPez1YgC6bkSg1gIS/5q7IcnKceHe5HD
HPtiWrVtgSmcbm93I5PEo4OJ/H1BsI2tuMndXn1c2paUtAm3/66wk/2oLAISFTmkXC0AfHmDA5mu
PajzXng4j62sbAKZZ28QkPi0E3QGAqr8YwcYaKIsSH/XEfibDzPeiLGpoR1wLD9u0MYoi3xdmZox
8sU3qwexKk6qkHSImElsfrhhxjNvc3mnB40sE+2EtGqBIeL/kAe2qMhS7uWXOd+cD7MWkzp1Mf9E
ViLa12Aq1pj5D55V4I32k2nKNJctFagjX93Mo024PX5pTGtdJjAIrQhj+CJJ0yEqK633Bs44cEEn
w5wTqSRQHUS6Yo5UkVUjHk8007CFNTFqVkEgjOxASyUsvOYnBOI5ESNgbHRsJUbUjIMt77N/GI7W
YYFP8J7ONPv4+yb8TFfv/DKll4qoGtlUWb+dl4fwsjJYbTSnC9aHVnooC9UP0y54OV73sQlo9TBF
S9pWZYzRxni6/j9Tf1hWLVBHfGjsqMys9wOdtpDHAbku6Lw+dqAjzHuwRJ9id3PQEmeFA9p7I3xZ
OI4Q/hlUsNJ1nqqoxgdr62kvGmCicYTAX07x0rT2Y9ZQrTcTAcIS7uC2zJx0YM6BCTxdHEm89CcU
79EpQQSTV3j75lxLlgXXP+iFpq5uJfvItiBKP9FH1LnzgRkccPnRGELIX4BLcikz+VtEKfdR++aB
mYIYLtsYSb4AH0PYW4Vixl8XnAULgHJSXvok4yQd1EZNUJHYls5Rl6ueNblJfLE4q+6/N1e7usoX
WRypFPiNLTvPwmS0HnvT7wUwscS60AMT+kw4o2pLiSp8Q0D0U5ej4veHjpm/WxQcQyBdA1eIXsAv
ReoYjGJ01ExV0C4LA99tuOIUc8yJ3w1BKQmqAiJ/RWOJqTtS5LwOEbvQvdYkWkKbUSpnBR3bKYfs
jBJa5RXNq0IaZDB0cPkA4zZsG5LxoWF3OkGmTTpcrfRQV341/gVk8ENRH1V+lvNPNXmgTTfreD7v
L3NaYjgtOAzoDh7fP6O93P+u6g5xpGwNUoNqz6m+DSSliA0JWbfmnay/jCYLDVB3wV3sxCaz+JX7
4dFOGO0mmAZRw8PsOJxD/k7kRBg67SSApUkrXQ4sD1ZWIZjHdT9uVlHimtQkYmnQPXJeY9skbJ3Z
xtM1w82X/FnQ0tDcSHLDq2E4yPb23/a+T3yvshwnHgmK8P1nXhdqhIt8V/v3sHCrA5b6A2fjNouS
U1aphqXaykMoXBra1hYFO3JXroxQIICUAqb7G3MvxYrZjT4vcRVFz8Hc6IBozxHtQ6GkIOfpI8lA
VNrHwoXz96JNYfNRjUEkNNbR/FcAfyU63aoHPRTudgq6rl6JHyHvhcqKVWBU1tIBqRtrP9SP890u
Vh7h27qdMB/pqWldJMjVXv2jGFkCb8cxlmPpeOq5gha24i804fG2XWMfhsIedNEKGjkrkv1AMioo
Xgfx+fa7LlPvQ9ec1YKwy/rAJyvtZtLG4l3m4SObziJp9hjwPh/SdbwvrJKOuFMuUzECL7jguuee
L4MAtrw8wsoTuWs9vwX9X6DdDZwryMGtGz6Uwi4OfRgFrrzZ21sIK9Z8smjO9k1746LgNIv0Gma4
HOh7ZkPGeFQOw+ZyiYi9E9tWkneAEEzOLSucYR4tnoUIO0NnU5Jr4TKLD56tvsdrC/EQZncTlVpA
mBtShwT0VGagZiw/509vy7tP6gHI21yjum0QQXnoptMlTPZTZ52QKBXp4XeO/I06khWxMTjTmKn3
7tQxR9QtuLszBPMDS76AktCw5jDdcUgp9pUxUtqUxNpGAMCuY1HsjFFgdNlhYp5sdpN51s/KDJkc
7oAU6KsMHpHfh2s6XvzJn5GhgcDPLC8FQ9x8yW7Pxl0Pzun71WZatBBBxI3sL/Xx0GdrUqUOrGPy
ahYRYw9qirmnYLPS6rXx6VJB97274jzkMZU1s2ObVBK+KlqTVu7hNUUHc19x7UinuMh4Zio72Yp+
HMbf53AfZYp171tYRDDF9v3Gjx3BwC1uGHZDS0FyyQvAaEugsJzJsaBNR5bBwVrgyJ0jUVgDZoWL
xaOWkIazHjA7CD9PtGgqKzwVps0FX803h/rR60R9xwoSdoHbOm0DOaRvZ0hJXU1ZdKSS6SpyAet9
HquMvjvBZ7K3NjpqtY7g8w9TcjGXQcuRSKwPjT0WALg+nn9fhb4ucf2cwMcCJQI/oElmhMT5Hgoi
SDGHrGQmmwECXKX1rUxyi8UjZB0zPCwP4kTML3jYc+DwJzBGUOrHjXL+1JpyuUPwOzql1FxoyMmr
haMglGrCDqnJQNivOFv0033TJh57pp0aTA6oc6UOh3WHg5tLCT8pO+FhcSCaX9eG1YAlm/0AkeHl
YHpR1pl725ylVO8RaeVupoewiVGuiFMWMQj3+y+BtYWmfDCTl2FByfLhW2TDWHpYG2CnT1YM7RGj
jG5I97EbTcMSoGu0Wg6XBtsiKhqUlwvAylDKuYe8WmcTaxS7tlrGL0wSGDzZGu1yKNeP6XXbXU76
UWpaJ1yg/wg6ltWyxnMo2dvTF+0pAncpozj39vYAUxTGM/rb5uC6/zH0WTlR15025HAbCuJU6Qgr
7OhpeaZ5obqnDCZN5bNe7Shcj8lrKin9kbS0oxoyIMH90kUVWw0I7c4RSD4pywKD+Z2FRpfoR7Dr
nAb2wLSTBOvHe62twzDwwg7ap/hDoFE6wqoQCe9+iEZq/KyM7YIZrZRZ1tEDiGME2bXs9cLxThqe
8YrUhI5eKmb8LYOd5H5CWtvQDAXxT3smlZnGyS1gtF2ej9lgWYoZ1XihBmTQd/9o7z8hZeAqqRte
8xXnSt0uj/I21ywpM2L4yygCa3HsZVe4O/MDxgsmfaNLZr57MCH/AoxFL948wFtoKzDSx5ODn/64
7+/KjAgNQTRNpd4wxU/lcNtHvhmlAXWUuPbPJ2wuaChieaiAwUooKCMP7zc4nwizI/epEj3PC2Vg
E49SR/c2hc46Rp+i4/yfX9umbpL3P/HOnlUXjORQWr863hJH0rmnmcAriXxnx8E7rt5Wofjuk0le
IoAgwrz4pYskYE3IPVXPkHhSHMSwtduX6bOz6CY05zcSI06ntkVW/b5r7sU0oBYFWwyZR8D/LpCV
fB30pHO18eJ1PZp97+tf/t/q4tSweyY2THH3/s694HIk1Au4nOBA/6r8Awg72CDNiwXuA8nE8+w1
IUeixIUSx3IgiYMqkmkUa8YcDjV24B2kj+I0x0PGioNsGvYjzN91N2Oenxk3fLFJH3GHtGRUY9tc
gyCGkIlWEs9U/brk1a0fhmK6g7n8sPUWuBnBM6iyQwdLlM7Sryqc47np35XwhuqL1lVW6QnZVtfW
cOpWrXsysDH8jrI2jVDWNgJ3TGBXTkugied/7FRyggH5j7G75/dZGej/7M/XT3Tp/BJ7DLlfWanS
SDx2/7N2xy9nYVqTa2873+COILnfufuF3W7BQTAH0alzg2C01ty71EWEj40gAJS5M4u9cZTWzt9Q
pCALJw7fhD8s4dbzI2WSjzXBHF/sWeuYxiapOovEQyPOkj5quMohIW+TzPBUDkn0WFiD+aeetJKx
GC/RQVRw0w9LY65HILydNSK5qlviTXxhtycY5qZUa+WvGVxtZQ+qsOGaNG67mp1Bf2KqiWBcI0Wa
3TqQlChckCbpizcf+lO2UI4zWy/hFHKUVyVlnGLH/XomQBXtV8b8aKK7zPaeXEuvzr2cw9RIlo0x
8K5r22K7lm68ciQ7jweL5AgloaEDJZmI9y860KI+Nl1FxyCx2+dn9uf30hcFpDSIq5Gb5dQqBisT
x8PstEKPD7946JBm515LyD6agx31S/YUmKiPUCRMQy4T1AUWKpOj/KQarmMWPlENHg5Ywm425t3S
WHqxBz1iqbKfCmN7sN9XNAfcLjvlWXdmp48eZ6nSZOg5SkQ3rdsCbXqXSvtCNw7jAWESpVBm3Xmg
JS8xGqh0QXS/oCY+uwpxfheu1ix77J6cXfHBcJ0FHd9CwMD19tN5eKOVGDmEQC/oHoFV19fTZzAB
ifZV2xSR8L19jx0kjcCwPDH8cLdeC6EqclfMPd9Pzn8ks6lWNigDdCJ73+vtpP8k9RtfgTpww7ij
Y+uULIc1AEJxgVigG+Z+qFdPxIjZGg28g2cxlN5BRxPU0pxN6C1EXzUhx3taKNcbG4avgOWKGvYQ
BCLKRwtOdZJThaxXLNceIAbebKSrdsbtQtIxg9UOzar6NIaanSoGAoHSyX8vST4xRJr5PDg5lJJf
24feuu7J0SeUdIolyki6uQhG8bzFp6oYvdkMQhTLuYzX2VI4p8LqT9Hopn5D8OatIqtBlz2KCZEv
EUc1o/+YDdYmn8jlmRxmOKmwQZXsHWP3pq4O1XVX0gmF0QsKYq+mnYChjB13Jm8K/p9Md5UISMYA
GbjbVbncUezltKN2opNVCRzWFtm23y1mvvlUcwVcN54Zw4Yk9WxbYjbJjX/1ksB8aYz2xtyZm0Yl
OCLJLpwa8+suTJeK77vkrxAmCERz6T6hpp7GKha1cij//cJoKqlWasPrsMqpuVjI2ucyCL2ieyD3
diqMQAS8C10u0hyB4TArirEWN5T05MkLV+iFtKoYvGEJvU6i9a/1OQHYqZvwOrMvsxySMYoL1Oe2
hLUi8X0CFqvfPV/iZ+R3fimz3uqbUk08o5tgiTebOtR9AMwZFiDY8jXdJjOUObmlRvND0g6BxHts
sZt+4yjSY4ZzB+T4THm4yo/q1yyxOAvWe0KcvNx7rGZ1PjV3Os4uPiQmcZRtlcAhLoyoYKxHTkZ0
ungdRI+5majeAHXONkQwQ5iFPvkr7Q3kt1QqoS0eoOB90zkvi5Ue981tlGn6y47LmQA4DB9LVXnC
0HWr58viEkvPOnAf6sTDQtlPmBkcq7rbtjgpyH7rx+9gzWLHdJwxk7J9suq+2ZH4XFHT3C7ilaNn
jLvyEdUESxKulUxxQa8Dbfp8B+IbDT0C0mO80y4wat+a4Gkc2MRhocvBUPbKMFGNiD49YlK2Tv/n
vPW8aeN/MIW368K8RbPaDu4S782tfq9c1FLhXRZJOS4fBZfgy63GFOMy22c1hBEJe5pzMbFc5kpt
GuCTgfTtrc5mmQ1+uQBIxRzVTHEuMyoP+YeYtvuEtXK4+XkKeAOJjnXgDY+EOTiSEFEX7Vyv928Q
H8MkqJBEzW4n3w0hj/Nyb6RNZ1JNI7orZx8sy+TXj0jsmfYTKfUdeWzqJvX4rpqpNIJ/p2IaRTQp
89Lro5vNkbQ/CqNDrejaDGCmgDHXiebqpL9Tv1wOneVUqSwGEm7GlsvKAuenoOmI9sl+lXWijKcf
jqE/vrtzTh+cIUnjLHMpu2KzOPuIz6Ly/lX4ToRcbM/si0Ot1a+PBOG1cqUoBIP1A9BDJFo4JsDU
MFhdr1Vh6dU1eGS/p11QhvcqoZbvwG2m8teHNJBEJUYkLyrRvQq0HWCwsiSkTtKwW9h8oYexrpL0
H8rIU8rJMH8UBvsPiGoOUrK0naIp4xn4tdNzCRfBHcrpU5W58dOTQ25CAkZsYH2zsHlDkxm6BBJ2
fRogXp+I9qvWCR61V/+4rIFhJ3eVITFKI1cHLvPmXrS1UOjeHXMQuH4kwiKp8e8/aR021Bq8/LtW
4ZUJ1v54ounfUHolv3Mel1t2zudndVgTu6KJ6hCKdJ+ZHAw4K1+g7lzPDJdTUbP+YgIyXTVyV7HX
E9WyIjZXawPFzs1QdifrkJ1a1UgqYblxe97TisUxvl5Dl0IaFM666zTXvt9fkrjPYGmtD1Vs1PnT
W2SHE/Kkn4jtcMkcZuXkphVAXajejzAwqi8XKfu+VJ9SN9KTaS8raHLI2e4ABAHiujp7ZnwtK3f6
2cr5+STmD5PNX7dklQW0dtHY0U/dMe/R3SAWIOcCSZXbNlRDhJ8YOdRjtQwtCGeExcXjm/0PRsz3
oA9lEQuAicUYCN1tPfDF7+oEn4a2UpUA8EqHWuh/8Q3tN/CiKuw0HnTU8I7K6tXT+tVFewJmGLuh
bZ1JnLR6kQdp4F27vzEHQrU5mBES5sC4I2+KCGxJPG2qawD6Z27lu/n8PxqYYEpoEXKaeqgmMz0e
+9S8K9bJemVp+zNSjfvwpQA6meZh1/psE7LWhqDYibDt8frrDF9a/+qnjNOwZhX2x/Rl3a6w3Hwz
FM9rzar554zSYxW8nfEh4BNBqpXQrAQBxF9HOVoX079Jftr1KLo9wimcseKSLQXKe3GGTNAmqY+f
PBJV7DyDY+Q5TfFBp2HQeu1IGS47jHVPT2IRogUI4dzJSEa14kir3162xRIkfjD9Uk7D04MsWcJh
Iv1plGwQVpf+eBCCzUMyizZ/v3xA+xdYJKfcmxOxHZkjxrqYQfWSIQWKIGCmzCCFy9592D0AnamL
fKfuvSmd1NraqUIT6EY56fdzJ5ga0YiWBjUDUbdqBm7PVmy3yf3oPk8ViR3/q+L0e86DTiE4DScR
VIlRI5iS525+V3aqLsij7etRtb83m9NddpLzkgPA9naS5+KcrvWtenzYFTkgyw/qUIBzfTs1tiCO
0E41s0/KlaLLbcenHGN3FD7ErzneeQM/mKP4vFhyVTNvnjeip9EihcUENf3iLWnu9Jgl4313hgWm
eBg2yk7YxQ/KO3fjI3ggZZ0JLVDzQBivjXLF7nwzKymrlY3OHzSWPbFBL/GlEYoqJ/hINYIWGjXc
qWxNW6CHAP/UJ0s9J9OuN6eSEaaJPpdfIYw1etY7mbuV/aGmuTVEsFmlOm9U/2od9pomMThUKAgu
vsrPg6GMkFZiv5aiElXkYpDAOBAFZSyzYkv9UYDDEDs0/YBL4JKffnw1DRPd8zhHyLthzXwAJoQm
H5wlEW84GkUhzBiHyCiredsWYbN12hbxPAaMJgB4Tcn5+ktHh/mn/U119qnT/T+ih3HjsZZh8SEh
HK9lM6VJMQaLupnxEuoeXEjlR9lTcVUbV+eRZ7gMJgqrUT/WLk/Hij5SmHmCBvAVLCnGoVqa5gm6
UjeCoMvW7zZ5p9i/W1nF90UAbO6y8E5h8/Fee56rG5ShKqbMI2dAGo1Xnd1rO2UqwvJ9XPNhGg2Q
4spCgSGnT8aoybVLmvgmbtgA0IB0RpgiMvTtVa7vIctPpC3WW7o4FSKfu3FeZCRSwuQAVLPoQiM3
ulVJpczvJdt4QId92ukj4D2Icg4fZYqAE8kc2ak3PHOQ6FOU8O/Ox2bkaBOdzmzSUgjyETU0pYYw
ZO4VRpkcqd/5yjmG0tlq4Cmmh7qIFI7p5j3FkVFcuToDBxtyGdcCXtNKTA6k/KLHdIcu7S7Igaxo
9tJxggpOR71k9TmopCbL4FVrLB/lqa+jMPSYssdPtio9wnGBk6W/Xu3sXjOXU8jDBK96Nr7TBATI
m0lEJSk4xOPQnmYiW6YfHZ1+mqD9U8OCJATBYKhAkyzlWXDCzT6/yXybxzMhhqk101Boy/qtNaKV
mwJCZDdAfPBHRnFtOTzRcRRNHrgUNch2jttTuDXGlJJQ9yxMuJEToRqb69CLCpEDMNvlfzvk1Yxk
0bqms+1AZwyCrtagauyJI1c6Hzw60vq1ws03uqfYjiyxryggfgRCNVXmW8fDn1uOUfncGM+FkwZ1
MNJd1NF/JidrvLCVPKOZf9HRvn2J6lPEeOOeCfnNqSU1yGwe5U7xhz9GhLHxbt6R0r/W7yEOAGks
HygymwYrjL3BAec4InTKAoIK7F6m095Pv0qust7el20hhCO+bSvVn9r6PH4z3Gzl5dFIMH3OEHIh
yeE+nh5rMviR/LNy+fxMgp7FtYHGk/gEUxR0WYUpv+8runOSQ2y5QsGqSngVKbt6sBCvtdcfFZSN
2LWzGbk/GqVxYrpzkeE63L4RbmpyX0SR3UV6ssl0w4cFxPpLmw1xU7/HDt5cspFcPEqKdVZeujQi
4NOfesjcgY6b8rq4LjqkCf+0GhW2+t/u4qbUTwXVgabr4KChG27sDf1JVG7lgAlD2fYjODRD6/n0
X/Dd/abu37BoUDY0HLgJJYaVT5T7bdxzgUCIP0yOYObTVm/v+UnvunNEB11emEIsNEflcVCZAj+O
2mz86hwq5pMaNZfL9bJ7ZcPrQvOYeOosv8Je1/DKsV6qtMjS490sQrHJeE1T4GEecZNkvw2gkn89
6VDSHDRy2e/tiGBetbLdEeIXBhyZOjusBXeBa60K2Dz4Z06bfV/EAodmcy7C2T+gEYTTPwBcf/c7
hTx3X4agpg/Xz8YG00xEk1UPvaRVLU4QT9Id8qMy0rvmZkAQGMf39fwuqVlwvEQpmn6sAusyZiJz
qEgMtpuxrXoAZX1mFgQE3M0hfhT3vac8uxZoXp7C/Am+dRjypdColX9MkpsbUjLmOnz7CTCPgg4v
RHviNLScNDGrNRHTENt4v2Rz8adqUVjJzN1EVxUkouDFd0kWqJmk9CJNmy3kBNrmVwxL130Lza4f
rohNgpxu+pXePs3FeNh7C+gOakhDQ9AG7ZriyRn8poUYEDnY8vGOe28JGC8Ml3sVuc6dLEnVex4m
i5HB819+iXZkG6+t8Kb8gmCJMeDmujkjE6m4t4PdNRImGLKd9xMNfOYrp3PM4UUxhKDmoU0nW/6X
BCminz4Bm9BC9ZFSInn7U8iRKUxsCdv7xoCBdEl5fp3Zrh/h8KWmhA2On06mWx13MjlZ8sPFMkxZ
+fHhHYcaqe0+73K8ygh9XyeM1Hqmkmj4xb5VuDYpdvhU+VqeGX7DAOgyvJa6weITm5sAdUpFqKu4
FYu4zdrvvoZoIIMIA3eTaz1uBDXePt2s5U9lXPZogQHKlTxtDq502sBO5nNf7Tpd6FI5HEv/R0G/
mI9Ybh75jG/sCI/s5sPjlbbEMLIRJSsIugOcca14kK7amCpYK2IB/QakSSDqPz8sbELLcRUbrZ5C
mknJg8l9hRShI4eSmPBDj9taUAvRiBuvFORGsosaLIFN3DyuLxVTernLDQs+qIylwTfLV3FsGsil
KLjwltooOMKD0acuQsg11mFINPbAdW5S+YXafav50dzsqEdye6Y4eLo2H0AHTDVoDO874j24/0JS
bTKYHOcwK3RcNQ9zsSP7oCMhxdg9cgmAqe1yRbxB5ZZkQgjLiBqawGE7LyVHWGGkZMJLqj4eYy+r
clQA+Oztm9OS3xd9USyV65UzO+JqlUPe9P5hmk0l2QO4VhuTeGBb7TTZxS0EY+ioKDaOqpwo7h3u
CSk6vE/ncrMTnrFtaExe9rBA5rTIzp2xK5TPZG+ygpcmibKynnoF9qYoIze/HIQ2GjVDt10O2idk
EzkHqujE5SELYrlf3g5UL4g2OpvxOGP45hAiu1i0Iz/4gZk+vJPbxUCf7F4pN19Mu7eDCErVHfrE
OagvJURvIXEO8KMVSg0p0AaKgAmG2dpg8rJCH0FAp5PZgoHKKWpGt8s0KZOFVxoz91UuU76Ptdxs
NT6srKHpUmxd7y5IJy/HUOPt5NNTm+gaE1vuYAhSwLIAvZWdUP/J/lDvwT5hzXMcZxl3C3UQPnYS
+UD+nUvmMf3OsQwown8JOmxUUOHw5oejR+N0CjK0BrHRomB6ukFQIDXJKj1Q5cPeeyJkX2/AXQPV
XeeqpU2WAZnP3W6KppuepWYBFfkwZqvwdvMvZktsPYHKIXrHJu1qrAP8vvAxE/QjD0K/rXlzo/RO
60oCou/0UfCJ5kiYWTNcvtqyy85VlofkjxYUEBWDOH4ybBENQ+rdPdd43vmwvl1KApFCIfQYWIy0
SgVe5TkNZKA99HSdrKxQVS+4FmBi6QJxq2erdEuSMRpPQ/tgRBkPCjfeKdXJougGsEl7S4xxYeYM
miYFq/8LtY8SZf5+TiZF960uGvKOsp5VZPVfNrT4UUWRmNXubz1hEmRcVwzcVQl672kXPxQZZmm2
8mLk9vZ8p32N2Dqzdh8JbxfK4HoqU9FedqcOAJdn22VFyclMz9j94yFKLJRbCemFskTjffH3srEg
rvF7+b68/G+FjFlBxHNNezceQndDVjvnycdVfRHXlzWXMQAflvqe54yJ/Xq7QpztNV8WniXFzWKd
o+QQncd3t0Oyj2FddOZfw/m+Lxf452IY9MEpy96119CLeOp3WPGnJYopniKV7ERPybIyahsMvkzf
qKLRplfcKU4U3XTP1d6VVIjNiTFlw9o4/h8O5ZyL73zkfU20kjjzQN+r4K4FgvxLMRLy/ERblPk+
sTRqSiWf+wCA8I1RfqBnp+wppZqe5j9ZHyZjCjsT12OSs67Jgq8HFFbql3qjZVSwVioAgh3yABli
0hqPSvyn2JQXojdor93E8D+160PJHItwTr2Vwlpgz8vu6S24/EWIsFA2wHqS/RXYXE6HNyCNaRP0
TdyitkwcwONVElLnxt+5+34HXgYw7KWUZMW9h98yhmO4CqgYil7p0egwFChybWiRSscvrpWZ3/IV
zif9TA9rEhX+NT6jh8J38BFLrnytiYyex5j41evxksbs4D80gmV3L6934y456LT17O+ix1nlbl+5
xvZWQH+qVbsL06AUXc03RxdClyntU3mKEooMiqKW7efckvSt5Xx9F4OQ+gCaUZtRceS6xwgWpox5
U7ioCMJ0jRiqZDfO1KN/LuAFcxRQprmaUBIXQWpg+DUPCVcBnNQRxP8Jb7it7QnJj8d4EXbG22+l
odYNdRCXeMZbhLwVcAqweLeF8SQGrrT/qUSxDtvpx0GiDPshnWsI39AVuSZwBt/MRvXG6CDtWEAg
7/zAepReMZtGdSgTZK4CvcRjlhuH6+ebmqeFO+dD2bNjXdEwn7dU+qBVzyBiz2sKREkxOOJwdWnF
+ItRscP4vFxCumj3yYw6wU5g72AGgmWrylxWQSc1rygyoXKuBZQZJ+krF1Uph9SFlVa8/rkXFswe
rDyL5lTOjbsxlXw7Liv+yu2Fw7x8GQ/rY2qib+dJPwOLc7slSwNMuAaal+ECGUr17pWHvhexUiFK
BcZZb226VPw9hVS8eBXrlPIqAg9wjNMiBl5KDZUhGFMRC/eYHPnYjlOddSVRDhmS/iZ+m/nWp5hi
xnVAzUn4mYd0+Zu119YmsZ7ErBwhAKuHsUnzDWp+o9Rfw9Ihsv/BG/8rbjnxf25huud7MW0ieesC
7NP7MCcUE5vPqWNtjvBf0kAt7OLoiW1oVuv6OOnsBbYalE5V+Zi4SXoZXkHNYebL3bxAgycJJMHR
z48icqSmckJv2l36hEkxzBX84LfcrEWjIds17EgL1jrsWsE++z9UgslX9wZSK/XQ+F+f0wd3YIS5
T9aKcYxpMOYeQDeSgtFyfeKYPXIBbAM8t+WIN11IwCaOQ1RRDtJP+QWncD/xqzMNkZ3/Uy6GPgZg
/rVAC1U3jZUyPE2sB3a+GQR9ipi7Y/uAWaegjxIkTz6jJDVn40Tqx2/USznbT20hvrcdVrSjggWg
VtbdcaLS4AiJaohWqp36IoiG1K72ghKTYUzFNa6NvyYP/1CWT4EdAjpyuQM6+3paZR07BTKDv/iY
z7qgWfXOrdQobxDwG7lhj9XGIytxntLCOFR4dkIwjL7fkywAAAJWR8HTbiEUR3FFySrwEqBpUzUN
u15ii40HstVmJXE8Ur1SlJm1ZbyuZv83dFQCPFr66xEANaXWo+VpSjCVHzYEtJQP3080eFHw5nlc
SLvoDQFiFtd+Gr0PQXEGZDvdbgMGOefGXZknmqFkQ7LheBVySxQKvpd7LaIdID23sfQNc7FmQABs
5vUuV3Eg+ldMmGjpEe0r0gKsrtZpmugj8brh3Id5t/QThSqm6TEH8+gFRVUYcLvS4x0RqoZEh8IA
Mk8FbXftaQhKYgr7nuPLsH6JCNE1MFI//fhBKV8Rqsz6lJsNumOrsXW6eqE+jIuWlgXtoYqjgAYM
3Aj8g4rKqqlYXTkchTnkMXK74KbqVxXH7wR6FFM/iNcVQfZ/E28aqvc+e66igOJFHZcrPvXlVUJJ
j5dDfaGY+akfp+4wtoYyWMZJz92e6bOXzjAJot3+VV5K9ole3pmh4YuDBoy244eodPRB4xMCdGk6
J/+m+lDi+3xYBAUQph+ao5QvCzU/TOdgFn1MQVCuuOe0J4u+SbVWI8Z+I8Slab31zGtvNXudpzmP
Z0O+2gDgRuSzTrq6WW4VIAFdC4ftdLnFSMt9SGMPeW5232Bxm9AycE0qb2A4WIQ9joXhCqTM/ObK
xXHJBqCeAobEcheKd1Xp+5U/H1S/LsJyAILEJQ0qPlm9+VnTXbxihQmOMf01TzKbWItuXXSjFODh
bqotdIzHxj7v78pr8gRpRbGI7eAgoCxQSHBSAZJNSvtUEoXDDe5mL9hRB+V46a8kD2oHHp8mlmfx
lomBt6Sz7vFGmSCHeA8JVvmKgEKH8VT+9YapkifOgdmvGzlGEu70IZ3CryBljNOwbSwxc//4I/xL
hswd3Lakcg8g4Kmyd+4jg8E+Ph3Znh0bCMBBwX8f9v1enHnLnMj9ho2nDsNyfZ0pBlxvk9zral6W
kl8I5W3fVKEzjKKMu1NymKXtss9Sn0rrqZvs+bmL72fpdXUGaodUUcMsjg4fmMQ4g/CswRpYUzhd
c8aOrQG4EOFhO2JHFjt3sAwXcSahu8wfigZYGmdsU85Q8mFpIXOSx/I/WMRzLZmvp9VUU4iurHY6
meM6oGAt10nH3hmzA7agCXmwA5v6eSYmmiCWRBafegacsqv7XS0ylr4twGssQtYWyAs4mCtwXKnT
GS0uYNVhh5b+1knxZodZtOGtt6kA86h4lg4gkRB0HC9/os/gKemaD8n++RGLkZRvc5rAevxFe0C3
FzpNgYTUMQScbXh68fvRmH8tSAX1OM5GJpYCjbKmZlQ1YajCAoIPhxC3fzOT3cYFw16fYPCWo0cm
bPkZcEFDMj/35lTMFimsX+tyvAmy3NuFbGB0mqt7SH61E0tmsOt/E3xnYjUTziKrXzB4FteySuXY
jEUAaMj7kCANV6UlyBgDO9b1wx03BuIfwgX1VXLtKQT6qDRGDm40QRXJqASgb/Mxd+lkbHzsxnmD
vPxFKF9CDWU6q2OahmmODn5Sd/T2UB6RLovE00kLXwuSLLkyKT2Up8b9+53pZuy9ZVaWPxEhMjgv
z8YH3nZS1sg9FmZQ44lHZ8Pz02wFWOCfa0azAsVdfMqfoncP56RlZBu8PdcnISVL9+P5zpxx6PLH
NQQpJF48pyblR9kMYGJ+EP8H5j/HTJYFet058rJLuEtEBUXI5TX2Yz7bVzftyisN4/ijhfvS429r
kaHJ52LddIdRukU3x8/NLk6N0NdSMwKdVlT4hN3c+4smUhmw/SEwgMYYXRusIdFhCWVmyE888dOw
hGwtibHI4j30Hfc6ocsrc+wpHob/reImVFMwcDA5ogMpuAAZj9vOPIzPfl7QIK5XFjqnwNrArVpm
q2k/goyCErJ9EZqKXea8CoNdXmNB63dXiK8/zybjca+h4fE2rm+Xroq1I6/QQu7RHXiZ3jwjuh6d
fM/KldGH+uEmOmkTc9gBlk3QPwSTQ12qBIqtM2BESRd2MMbag0WXuIKCo1iVHceY80uXy99sDmsL
5a7M+SQMtevGY2UuNazEBLy0MENdM4PI4JqU8xPBcEQxP4xeRHhTRr8aFdUAOa2AiWWoWhH3MYIV
IAGojlSDnvEGwtRDb5aGpx+6eVCNVgghmwn90cUNlhHLhOq1gIoBfo6qd+MQUPZZQC2AZd1e0Qhu
V/kitgRdEzWTQB8ANx/eLgnvrDKmIW6RCTtDAusNQ520aIpgHsTV9TljO2JeHKaOBvOMhHSTqmB7
cP5Yo87F8F80DKsn4KVJMb75Lb0SsZgq4XrirYmuippQL1hG6/pDK/RBDe0y/H9ppfpHr1bWRoZf
OS6nLkTnDgXxfi+Tcg4Us+2jQZJILzTSP28vGA8wW4d8QvXxkIkxWsbMUaMTn/PwwiRI6HoHPiit
aVZ4ViDf7ovd+bWwazPtx+0PPVfpPFoFmRnGzDbDLdP0qhbkq4H16XRNUNSzH8q2L0RMD867uyV2
A33dDNhnMm38TvOGzYaHLJIN3+UOF6buXA4kdVWM/hviSc3OVRWs3TV2tjG8gyirTkb4U/T23ALv
jM4nhoG/p4jEzmmYMZ20qaFefXJCW29dycjjwtIgaB/QSKOhAUfeUjEoEIO8K90wUbNJ3Tqu6jvi
rlBTSk77bRyfFCrhGQQYO1TQN0fJwwzcRENHD7DhNkM1X3X3MNG3Zt6hcxjLeLkgE26GAoubeE4T
Ix3HpjepQiGSQ640oKmrQ/Fui3S66E9QclOjqUpChVjyHGnzcFewYMhCNTK+4csfZs26fjvnTFBo
ZXYF41Doxwj5eXd4OmLeLYLZQ8aH7UvUMRVcgxSBPQI4C8FeV2PJ+1ypt71XbmeRkiBynGTVuWw0
J3y06E1JRsErw06tz5YlC56eC5aN2u8JhOkV9CdELVDfjc1RnhGXpdAbKuo5Jz2SzmIGCe+KaVKS
XHIqDakS+gNT7w008wwIw5aZEFicnGypC/1GYjjAUQ9zqfrJER0YGhhwYSAj6+5Z98kyt98MWXFY
Ljzr49ZXFri5hndkGbeH3ggdYMURI43bHmv0B5Xpu4Nybl8F4xzC4C961xE/Y/F9VmrRQ+8ot3Xl
oL954kVW0DRmzbv4WiOVZ7M2R20PdZ/976BL5xOQDn4nKix4Q0cJVPMmidGYLeHbKu1o98RLyNhs
rpcb1eH54MKcHZhWsSJmnK+9G2+xpssjwXqOLk92yabfif1xnQSqo7wP5RAqIHZutI6wb7954awa
sO667Q/4hEeZ9S81HqO5ZWh+E1TiJO/v/KI82WnwNVjPJ4E811zmSX0tShbmj/9garrwWaERHeIH
y05IR+iKRrN/l0J6hHQp0TEUB6wFMTqxC4hcu6E6L+mH9stRbYQE/g1KLzthz3nfBby2aP2h1QNq
52mFdH2JquzuaktABwlxujj1eTZWGJVU6pkbxZ3HR5RTAU0JfRiASKg4/Ex2CID9sniOGJTNVXPv
dG7O4QOvpyxgJAAVCmMt9DyXvF0gn6t3S7GAmCiDmEI4TAknOUh7BfMNdeZfgSCDoAZeCw6KhP11
S3C8LKs8lxUdmV3ab0+HDV1/mS1c0VyO6nH+iBPV8KlHtw4J1GvFetDHbMK0uu8q3Yoeg88stC5/
rMb/08oH1VkJHlOvAbxHtSshNGLKZmqISme2l/7IZ1GH3R8++YsA6oHVnUmqfngbZ+vS9NzzA1CR
LpdJydc1Dbbe2eBNsHmsZXz5kpBeHLdfLOik3xtNw4NPnEQHhjWrfJBN0wmztMWo6XdFAr3FZgjS
MoMXJgiXOWMdGCh+8qigeDXkXlJ7cnMgoVXpX0hgaKL1psYW2Wa2HrpYwhH1S9GsGZbNLXd1j1tF
qzcNAUfj/IHZmZbY8h7BqOEu/hi7CpJElIZnm/PJE9jCsOnlH83cksQ155rS4oHwx04qZlTYfAkJ
YEyHZi1kXan08hNXEkEQVCbL2vGZhlBkByt6ag+1y9tDdXAjEB79PkKOvAqdmp8G2Z0ewRzkqUWk
BJ7SNZ7TT0G5PjgnNsiOpcvWkYOFpjboUiC2jfoWxLKRxD/zJqzwwNdE0Bv0hHiOKlgw466gDyRu
nxxs/lKKE8iMU0QwaD5BQ03xlAOevdwI7NGJsmp4Gq7e1ZH8VxNl716pWDNeb1vXVbHh6zd8WYLe
98/X/RRBIm/J+GTwfIZS/+LSjnWg2zvc93Z+DipYLirTBje+mCR5HxgNlb0B/av+zQ61Msi60oXB
g92m5DgN1zw87Ad8oVXZFeUw++LZ92q/A7Ah+XCraTqE012+aVUDPpMW3LaZAwbAP6XtIpyAGQ7B
3Im8XKsfDgasDDDkCUtXUAir3Ck1pmSCWda2Ab5kn1fVDVqDStH4IRGP2r9vwB/wolsI9xl/ZuH+
yujiQVoVEWFGXt0JiSWrvLynKSgZCuQsuCqk7FaS7pgu1f/ZxyT2hbUf8jtKwjI/nW1v9kqjWN8Y
gRpO0PP4XNKd3Y/RI2KM3pXNb5MhzGLj2QFfWmhENXXrYEyTnz54KhZM12YM2nDMQpkq8j3UHn/5
53VqWFwP1Wxh3v6V2rBy4/YqrcVYKKM3cegpA+mEOARjPhaNJm10VK7nrlPz7DRV1w/0in3OMxZE
1g2ku/cAmw3zy6d2Ps1LNJGAMpetG1JPFf4/6dXDepy4rjoP9qEzYAl8kOO7W8iETe3RAzzxPpWE
WPOw6jeCPaQ12t1BvxaAUxiGFlj55Ia/TZaKGrtN0Nuw+sGevFghUIyk+D7EO2XjGoR+BKY55TNY
+S3ZfdiBn9FV2jsR79JKaPXf7wx7QaaGcgGaghrmwpTDvRsrEJslDFpBTuhduMP7wxK9Xlwewi94
e7wVtamSdh27HQVTAKAa50bbziFnnoY3Hee9X2TCcxyvNYqVM8J4ui/XKNvkuM8c5VQCZuxBkQlT
sDdma62FEuTWg2+aqgEVtgxTqlhh1K0hUAcU4ra+6+HnNNBtZepojJUzwbyYeU7eLsWPyJ1nKEM0
mgUcmMo+OcODbKkpZaYbTK0KG5IUDv+N2z/grJSLgxP5QrZEJyTOH+uzGKbe9tvjBq6M3oLxvNaN
+ZmwPjX29d3iXiF7KMPrkemKdBnS6AWrIDRh3a48k8XpwNsdA6e/weXMJxYuyablRe8F1wRFlLh2
FitDAL/9T60MJeupoFO8M8rQxom4MZJ5FFE/LkNzGUYO/XF7gp2RBmZwKeMSopPjkZDOa9gucBGc
fLxfPSXT/iiycaZt4BpLoz1S50ukzRNcsLJ/o2fUZRZwR103iEaJyc/yG+C0hW6pGbYpmTnOqcOx
BhZZSeqsXe+Q266k8a1F13q/O8WrU65lRIrTED741QvBxdjiGQ2XUh4/A/PCSUADxaZpDB105Lmq
vxtGZrO8Q+LmJO+W1sn2jBHckuMoiqZIykcljbIOkAy783qEkTE9vsGG81oE47KyJvMqqE4sTL4Q
ZWJ1KHSsh9tVEFphmxhup8UrnqkM+SxIP28EdMQPBFAiebKo1OWzs7ZbCzQv8zt4X99rE2IRXeFa
uQUYC6NE074UGc6lLqbheK6hEZA9IhZsHkDcEH4LsmA37sZud3yumQ7Im727hfMBEzajXnWOc8JR
+Du8ifbcaiqy0Epx3mVjrv3eXmqKH3s8YZBLNoYvT97uaDi9ZlJYJ6qmLrM/DqPZehbWy+ObMqBG
SAxR4LagFz5VNctcCcfwWKYfY6xKPEP4P4eTGuLsfXQAV7XnEMU/z2KRuLke4mkFBi4vyOekj4R5
CeTQWetLIq9vHnUunT5HbGwagy9680EULELV1/0BY9796tdKwKIEaqD3rylayRnJmivqbLdjFx1N
GAWFZA0+aEWUabxAikV4SZNm+KwctdlZ6vTxYXj8ZpWcLXet1VFmx2N8rqYc4JdSDBCwB8DXa7uC
EDD0U2lM5zF9AaSiQdC4KDtgEmOVQvFf5PtmRyv2cIW8OMB0fDCM2+EGbQSVKitwxvvXl243G6ho
/QXliLGhYx+0AHVDt0D/t+tB4JVPzDGl3oRRfoYIp8AVxjS3H4HIp6McwBG41HWzHzXaYWuxgnPY
nITLwvgodSzSzLW2NfdWM4NfhwGVcElODF+eCQ5cVmKRD1XNIh1pheK0cYaps0LlOjbmiGnKBaYg
xUng/P9zvCyCENPlfmhPe9tDUbwsa2+lXsfEere/kq6/YGnHIACdA9A1uXzKzrJlK1wCFhZH41OA
LNW3Tznl3pc/piWuQS2XXDh6JTyOw81b7AdpcBsV3l2i51Qw4aKgVPnxcI4ktRaGldoP2r/NE4fi
sjW2dw9d9IYV32naJjYfU/DjW+1Y4uqWy85uTh1lGajeZhyvWX/d2Xf7u3SrFYqWmveX4Gll+SB8
REMP+ZOeXlO49AX0Cpbq7twHlqso8XhHtV/p/KBjHffSZ6vNRjw6vfmiYe9KiP9YIppnQiD4sCKt
Rfl4C/3GSI8x5NeBwlMdB3/Xl1ymLbnmSQuSguonwl4demssK0VrmuZ6D/CJxbS+EsDq6KsCYCqO
aNQrfmpBP/VszKfDxpzie7tXG/r2+UL2IHi4g1ho4Gwr2QANG8Izrq7zp/q1HCFnuZcKWBcUsyvX
YLRP3/OS/V+xp9HNeXqY34/R5/ouiWX813OwBmnrvX0rT+h+RDo2LUjD37+Df71Ctc+56Mdy5pqf
CxdsXfpQMyJvUISiSpiJCka3zkV9OUAQrA2d8xgN1PSkW+7OZ1S0VKbYwpGn60GqoayRLaeAuFKB
nb2M5xu5v44Kc78WOEFKe5b0GbKiuLKfhMsEarqn/t5NaPsRrOrWQbTbE5zRGnVZoGPFa1vqajLp
dJ2f+5IYJFwb9j+6U6g0t48x4oCghRBp/bYOU3Eliw1+lWhsxyEbzBfoK7XFyBG2x7EC4Ls5amkC
cOVEGtKG7izniy2SGZLXYVNetiEKrtGjWLSOYSS0GU2McPyw4Bg5GggvTbj+zTx82eEk1RB0xTAq
KvKYPbesYNJnYwAmRu+sq79pT9oVZAQMUUUKeN4y+YZVcBLWBqabwm/Zs1GwoJ/SAzAyF6k2JpQ7
lcfKRQv/p1e6Yqm0NsVRFJ2VRfKpiuPKDm498NmrouJM2XOpI+vxQ0skCk9Kpr0LYhcUzlTqYMPN
i6S1BkhJtmOwrTc0WxBU9iwv7c6TMjIFz9UOT3wyF4CqdgFKfOWmtoGlUFTq7GHdg+Q3DM7+UkQo
OBHQBQJ6CACMF+oL8ysCwxU8wqN7JP4/qogHliCVy2Ma0GLVybtvoPBoZQoMtM5rNoSxhryS2VSH
jRzH4L/nmFr2APpmnkLgFjkt+CGAfcnhSxyAH92EpQm5azmnOztp7wunf1WGv1lzwb/5fEioydZb
HfOI3Mo9kgY77fAdVdLCmi/u90d8o/GMuDcknJWWJ6yVwPvvkg/c8gEovjp2fIrRzpJkEft3ZJ/0
s8BD9y++vm/c7px3lUT3EnMRHNLGD7sTgYxW5IqF64HheEZs+c9giromCtJNHkKK7M5aHrU/s+Qp
T5uvAomuBuBgvLBTse9dltHw2pZnaZCWgYb4bDCnECT3dQYBM2lR7NMa1TuLutfqL5li4nV/SqhO
SoQDWsahmkIW/e6uzCaUqtNQrl6KDTHRv4464UU+xgK3vCc4aOlpfge1MjnjZm/5lL7GEnJ3zkuD
gZdMzo3cBkokQ9mBZBdUQzPm+lQCCxJnFWSdUV26vmlfSbJco6/MYOl8GH4D0GXIyTZrarVNkkp0
dBhzvOzneGSsdGuHUhf8vIosOlHpSTc3lCscsyGsm0Vz5uf80+2o8PXZNOjSm0nQ3tsRjGys/PtE
zROVPr6Mi3bhqch58zJ5eafadE+WaxbCpdvMX2MmVhcxjeOeLsF9FQPspQCbG1Q+yj8SlIpLeV8H
8SeKgaKn8cws4mkbpCBtUkGCJQD9pjt+BpKUfWkjAcjMUSmWDItdm5mgsU6FLii1IjuIVHHETlhO
3Y8lHkezRp/JSB8jCoiyQOI9+UVgKigrryzeofKEoLD17m3uIgQfRDXi8k+XYqH8EGA/S4XLeyGn
gcrY6cRNDQYnfu72Uyb1ct+2DunNYv8HV4d62q0LZmLqDlgFCgxVW9WBVrRf5cVwk4/QfrX7sJzH
XZpq/f+Ob/j9d7ohpfnbHAT2r//zqFLmGVjINnhY+5GSFXKC8w/0kUgqOGHwcMTRAryQlLI9Dty/
Kx/IHbtP7nH7CK3OY4EQ9gROXnCcYYicvY16kvVofOOrPO+bH/9v3TTTdWt/esTEirbPA2DsSUnz
pbBgEf59bAMr4QgOlP54xiCWdpppSF6TGqI/7oQBoNCw3GJqH0ZHUevuZYH8GvCdg7MGIDDasJp1
p5cOsMdX1eBs+pV0S9gD9OuyfeqitGsdRqOjGq5VFl4iI3I/enlRBt7txo4/EGo8npfECNfK9/SE
ZsUD/XXFKOA3ityltuENEbzoRmTGaxAF8mZeDZdylERAwxHGTtbKnDn3o4mcEwyvUyyWeKekUFPa
P46bUxCyo1Plia5mVjEHTEC64R2kpQfz2RMjV9caEZlB8XKMlEnbFtMtSJibu8HjCBfgZR1YiXQG
XQ4mV9e4X5UahJf4Lr19LE3xqSNKFGz+rxeaQfVmmm+NApDKXAeCZcyvlFCvITscB6c+bjUiHEjr
zAaVbvwhLFwDq+Tqfbp+zGfPwhuFdJGsc19g3Ab2tMj88agtGEaDV9a+Hx/5Lxebczmbp3EzY8G/
ZqaCrhD5HVnfGvXFLobiIt1h1Cdz4nquXK/Fn2XZdqfiT+BoKQrz/TqTFQuCMJZ2H6NGNx0NdrgP
2xhhOWAyaGGvCtvnazsEBvAiEiLhwHsz4etsSthFZ1vPLHhKFfNPuBSb6fSEh5aYYgHzouyWoc9d
7rA1gPjxigeSu1QQymz7Hz36fP8w8r5ZP0dDUq3L7ul80FWMLvavDXHcN7fLp2gWGScH2bRjdFlG
tAHdjo50W0zVOG826494gXcriGqqwKDhifETgPXmOJL2rK1DYuZBFITd3KuJvuE4AXPDLUP92IXF
pcymagpY5EKovf3vIjvNpEAiQi5RZ2K3ZvqOrm1KUU9pYyuXX5Ix2F802Mhvt2hSWMOP4eyXWPG9
Qg9Ut3ADF619Ejyay9wYFo0Y6sqZJIdLfl+n5XbpvCQleAlpz5WapTh4nZsgO8jz0m6ZEm3EooRh
3qt8wGcFq7pygTgOG1ziXSSqvIFQK9VMSzYZIw1zXqsXbGV9AVpjk04JJZS89gFuOM9GPVx5aQiC
oyRFFDM82Jg0BgESkXB/oGSYhKmEi2GaXdr8vqmwqKsxixGoX4O6tiquyfTFYGwJKju0mKG3QhPR
hYLzgdl79644mrmM4U+XHCH0o391pENbe2Qg2CONtE8D3HDoFl7kPTlqe/3FLPWcpyLuyCfcQ+Qi
+ekI2flW7m2F8hZRxBRkKMSKGKW3nEiLf+DfDZVOEJluQqTAVisnolaj/KDGy2xMK1Q5KSE5qV9N
bmQ8SKwaH5C/jzXzirdsYsd+66JODBvkJm96JT9ShG0nO60qLb6HE8kDv8iJwjRsAQE6lRCmVMrz
j4R+/ZgoOo4sCIl9oGmkUcsOrYQKTmtY4qptPsXs630OIcYuCAApLQAs5UWiHz2oT9ak2ryp95x1
UC6osButRFAaeOf3wJV9ju5xadIkWL8c+cpnNgFrV2MKQsONpiNV9Pa9/YxTfZCn9mClcSKxXArp
+sWsasatwDNygMOG1SErSHkCxxJI/m/PV2pHWmybNwmXNClMWlNd1xuqyooKK5wu+WULRFoYkQm1
1caOmyTzZH9dslD80Rhy3suOa2J4oSIKHQKWP4ITJdeV8JGGviKazrYno0icvBZObq6R89BHDE7x
6Phsd7CRUpAINb9XxNGgpDZIdjlK0NO85m7WMhg5DO4rVgwI91QkTLufp9jhubbb/1vhuSUvRsFs
vH/yyfcVN8AezQbu3t88eIsN7bNJKvnHGDMEQmWof/S6gRxXQ1vDY7XAVZudkR501/hOo36mQ/uN
8WGRlmkGL+PAkkg0gBdjtRBv69gnk1ipGxGcX1iccMVeImyBVCo8wwhVhKl3e/SMExy5/DJmcafg
WdNmO89KbV5VP5O48kK9Nc+61xd6BXWGGhHw2QpAAPTCLd6/mGcyt4OSg4nAuhzVN041UAGyxb+j
e8OT26+GIj96TX9mem55lTgu/IbeCqF9bijKPeINrT7qF7S6noik8gRwG9JtNeX7h66OoonvVS/3
/3Yf7fMynW/obCOheUyDZXXtzc4DEmwpDG4UZsoxPGFJVvGMGXuH+j3LHBDpOKWunf+7eHr2r512
qYB+kHjkN0A0HwTAYEczMqOEs0Y13Rp/g3wKXvLhHtHh9TKS/sq+fYbaRYulSCo/q6x3YmtkhXg4
LuWEkqbFHolUBc5C96BJ4ap7j74xNcbghOJQuXEnlyycKVA8WDxstla63gsdVvkTT+/oV3OeAVBX
N5/zp64/yNIja5LHHD3hIbAXv59u9mCfhQDbknhUrG1Z/8eyvhXoIQLIucHJIimyHu/wz5bV0JKg
G6jblpZOxoCl5pXEqu6YZatXdiwokunezbpnO6rYi5nzlTXz5LEhRAPJ578f/bqCAu3BQb6WsOLY
RfkTqBVlopvWwNp93bHoxxuJ7guJtl3BnYKJFtBdopTGQwMnzWhdZZQFFSa8TXgzz86/lQhu5j0G
9Vrncw1RY7R3KJ3nySTkwkz4PLubL5O3c1AGee9yNGJMMlVCxz69cmTHf6R4X3KJQZDtsmjPxheJ
sXW//6BdgHpcwpCxiH9ImHH3088loq1WL/B/QEvT0IK3UMnhuzR4F8B6JqIapQf1cgEnSmbEWOYq
2f6iW8OdDqByoZeuHW667YKY++Ad2d8XmVOpTmgOETshitFlmJG2TrMl3N3ZGI9Y/L743zEk3KVI
se0+lB3pRUPnLE9bquL5FPSML7hJYJrLfZGzuUWCK4Sa763i5mLms64Cwsb1cLUBlv29RRuisVzK
BptzD5jmGxqcvT1iMI5yX/0o5b/xGcMvBAchcQ7ZqHsu63NRy0uRiKL6cu0nUNH5X3LrrKyrxJe2
oeZYP0hdT2iTUBXMIdevbpW9lsJquRAET4IQ5XTwfzHG1BxmXdHlMeMnRYw62G2Ft9SdrEDt4nM8
hlb6CMY6WBOF1tZULPE8rNenZ71QqQ/NZtmqdIC9j3GOY1RNrz2NTv+n73RWevfAifE4bw2a64yN
LXFcMVXXRlwkQG/QFdDMXE80rQXzAWAzWJJn7Tz5zZUHMy4XmXYdqprK7f61kfK+yJMBYNILpE36
uAVPEu4DQirFiy1WocCLGtZGkF5zFCBK67uRzuUDfwPJwA9+KEgrMYIAzWlakNMX6izMGQhgBZMK
kIaI25Gkh35jFs3o64jBxkJg+vUXZIXI79q1NGefd4UdiwnLLPXtkEjJT3E/ex8861KvXJO64P+a
zZCLaSgBeD2dKQbKa5gT5eP72pSJeEAmCps1GsiTv/zADHNcEynggVYl13nIswsvnuJ1H05U6oCT
NMeibYBXXcgoCKV17YJbigVU/yevXV/J9uiPKvurP0et/vBBA11GReiKwY156SusDsHJ/cxhnOb9
0d/NeWTesKgOePC5rUBUO2a581eP7tj2h9DlFqW3uzhBiB9W93tVOwvWrX+EYrUdNq5BFu+TQ0B9
hK5pA/RxSsH+mDDeSTq/Olcc7eM38q/apvmboYEJt1PgHmCHbM3yHlHHh+Q7Xzwjp7IeWzRV0Lqe
9psKLf+nkzwlR9stFdA2JViVUI2I4TkBXSauOL7DMwukYk9XahWq2YSG6Kn7tk4Gv2liZHVKEdNZ
RWeRp7XP0bHAIXltD8BLRAgXaSfuG4oo5I7MFQnvAxJ/DxH5i3QVYb5OQDRf7ZfGLGx4etUTxZTM
gtIEphV3Mey2dWJ/zCVLmvNV4W6B6jJDpQqwwMnfbk1t85Jyex3GufxZXDObpp+uu2T0NOYMIoa7
9F8s0SanyniIUHTUJUKe3x1kgjPczF+dqIMR3dTa6eE+i5Vvend+ZfUXM3Tup6qgZD7BTIWIthD9
leBXG1gNk7kYqzYG+IVWyW+UlVOem8ePLTUlZ6kI9gTegNfNzV4LkWbZAOEEzQWuLwg/TRpM4b8X
oJkPhs5FEgpk8t0Ybn5zNIGJ7BuHBSWeiz4YU+I8+dhZQtufBSPY8LN0euJlirE8Zd8wiJwdcv/M
QW59BacDV0gvbsSVDt4tTof5MULCVw7FxIRXk/o8IIWqCd5y2zbqwkdggoA922Zo8Z3rKKF1kufB
3aniY2shbMcPv2pi79x/wUJkMe4HiFdWSDaUCj/2WHhOYmUdLdUBRVre5pAy9t3ZBuXDshpSJZEn
2kOFnzuLewnZjTUKmIrPDzjL4VfIXTzroGDhBP89d9uHvnXfOyncDKyM11IE28JtwuNEI0Xm8j+M
MZwKni/MUotXOcx3J/E4gbQj6Yojm7wXEa3joTxySPZoYm5bSVauBW0K+SsyBC7uFrUu8EX+vGuV
Qy6dwVoNJAubdB9ObK+h4+394XnQJuATNBJyb9eYp2xOV+rdrK1NCUljs5iQCxmNkfVMoGNEKrzu
r5hmmFz1xtaaUBjvgHuIa7wepscNlxkZPlnQW9Zz6Ipgccq95zSmvJjh1Piqph7YGLJovwiH6Svt
O9wPdppBPuhYXA4GZ+mcg1uRx6S5u9RqHKk2BS7MJBKezrGr81WW0ud2TOLayXdqkfz1S3i/V/zS
ZFSxnE8ORnTYWrCAZZLB2E7JDMY72XwNoNd/E68M3CQAhNQbxUiVaZ6PrJ9RGVKouvBAaXfP8KUZ
gNCPjoDJqytM+VkeaGfMjLLgchf2hej0eSkBvYOdPj2qTqgZq7Rz4yeyD/WKFmQmAY4MnVZk52QI
BKgfcmg1EaIsA14LzR4PYcGtVCXJTInL+OlqkLSPH56c85stsXUcUJ2yZ+u3A1p8CgR0IBpXWa0l
LRpUifn3hIE+nfd+HP2kPQxNq98sCYVIbwjEHQN5A0mmftnSdnz1nb4H7ZEMfBkp452tslR3x/CV
cVLUH374gjY26XDXUOPERGAzLE/IdRdWvALT1YAhog3GA2oHNdMcJ0UROhqrsEFd/AhiEAb9KFER
mDB09BlIEMXfXzIwgDAcDSlI8gC9T2A0+72C6hrtz9L1Rtx3kA4vNdwBuLInURtpFpq4fPKul4Sl
HitDYz0o963ZeRhL4dxwH3TDLZua7pIhnuJvHsQurQfNM4fau66rChOZk4cR5U7UNDpVm8EBmnyX
YoJ33TDyqV5DGyvQpru6a+hAiQh8DjQq3+ZK/c6Yu0dVfRQQ6zyJ4gthRY7API7ikSABD69rxLBg
5Yz1hZZMtAcpeUivZs+SRZFVfh9Z+XFEMTnFY1V8/CL5fWpcKYy5vcCzIouw4iCyy2/ym8lJ/Ndl
pJXr+iE5DApWROmMKrruESa5F806Kmqce5I1ugq18DIFwLZA8nLAf7itOynizhwzLDybMmeSgWQo
CliFk3JAEHUzLDEoam+8tqTtCKkaQUUucnp66Ai5yEZHvt/YTOy7+TmXH3uRFouTcOUL9nh7mEcp
2ETk0gTAnWCrzyi9eNMm5fSc84+jDAI88/wwPcsBbGvbY+iB9a/ohHG1IF5ZsALlxuU+B3awTVfw
I3FyyjAwgq5QIHw45iVHHFq9Swnetz4JIR0+AUNao4VtPTeZ8ic0RHd20nN66yd4RZRUHpDWyRmF
0hWnJTBVFmpCnaM7iLSa3ET1uraLH4cSOOksqwvkrmbFrTXBNcgQwXiEXQ1vDnXf+y812Kkr97f0
kmNxK9AQqeDcXDCB+I9t6MdDX2QT/r6g9fEu4XEAdO49nz9GpnGTcXhLW7bI0EHRpMil3eJ0l0pU
9CKcAKkrJkbMelWiSDyaNuLyRPvqKuf+ivwVm/ATn/2k2oaZ/b4Zyj9e3yfsbiYpaKYumTdOkxkT
7wVpxZSgdEW09fg8UYR1QmzOmDuPYWuHQC8yp3lPsS44en7bkFFDRLTftHOTsPjbWmKOmZbEOK3A
Sv/FBKd1N1F8mBcMqLVA+BUFDJ6sCq6Cmo8QsCQs+il29uyzbsLV4ZWfgjeMp1cwmKbvC7YO9Wcm
LJFV9WfCuYzm2M3ACaGqTj543Ph34QwlGyhGmZo9K68gPjEVVXY8DMiHKhEGnmzvm7Wpr0REhEVC
Kqo8NQ+TZIZhO4nmIUjCzJeQG34ygyNkxK2GE2LxtFP/t4qz84NpW4rY5wIT3EEpUD0L+bVfjGn6
lLNnaTDe1EwxpGOHlZQfRdNXm5bJEbgsPF62fAON8aXbqsvWmqWGAsKGx7teQCs39iHxvd85j/Ej
3jPS5PC6crSwyIxOpfdH3CAkMa6kV6raNq2jaOn9/ZyxmTtEdN3ct2QJsSN+g9bxiEeVbeul5KHf
M96MRj1SY8WsBKc2QloYo9pSH9c/zjfm82RZ8wK9SvdOAijtSThHKa7yy0K36KIMNYdSWJsDjRtN
akxgd97qK9BkY3l1WiyL5SvktctE1znZdrqtnOKkY/5zmFcr3QWp2+1z8iskiwZKYRy96t97Jj3u
/Z+1xEt5lzE/wFzDJXZ/TzZxehDErWwxvu34ZwSwwNdmT3A9FgzseN55hcgmuyCRk6jj8S4zR9p0
99oPhPOsU7kIBgETQG+A2F10DUFcD50toUgizYxSStnQFp1krwDNZTInMBELqbX8kcxH6qrpnVD1
3RUil3554Mai1mseZCt6/JIiFAHDg2GyXBifBns5qn4C55SecmVrCRooe0Pqq+zx9/HE56l5wE7R
NkDZ7DlrUuiJbbHx9ZdWv9lZOX4xLpXadO4ha0O9f6f3rxeDtVXZ/GQZIrMbio3KDqlN5RScujhO
EtqLumR0zDeryDFVI2C1j7Bl/kk1rWMaMLlXQZ8+Dovj3SCwhvBgbXVbxmZHykid9gfOeTfSCt+p
vxYaXuQ072COFMwaPQCFTJTqnExBoxaWIw+QrPs25lFeEsCILBXqUY8BCj5MLrC+e6qqZiKvexR/
YyTwLl391VnKZYB2EiSZSUobG0BdJV78q3Mg59O69etEBdWVgNHDwcm5sT0c+MYViJbNK7RGtY0D
IFGwBPbZsUuOWKjbk/vXVvAQ9ORJT4xzUygJ4zMre4CSW7KgbJI3nEEM19zLB5ptdDEsFaVbVvJI
W3ejd5Zk71cATc5qkSLX59hdJCkFU/FuhcKfI1q3h3bry3NMHyMl6TYzB1YvpbntgitFgso0TEB8
7eBQn3WracrnvJsTAugyCZcgOyTvw5jsIn5Vmmr3tezqH2TzRVBlGrXC0EY/Bjk5D/YYd0D+RXdH
Pss7P+vxkyw5XmOKZK+HG5cxtbGBk7AU4+GzeAXXkTEGMAVg6dnE/Pk5x8ejHfwKR4ZKvFL0VxM+
qh/s73ugflJfWHWLMK5u2fw1jFHkA+y6V7+mNU0x8Iqcbfk70myNemNLJueKHgo3+X0cxqn5Dv+h
907+IglMSD1ZHd3Z2eRPl5jKCvH9qj8MeWQJcpDRYaTMdAmtIuZC/l2qtGgzr7BrC9/QB36+itfR
iUZAHwj4Rf0yI4umc492dWoG5LFqC+MoVTrLTunRN81H0iiS3FsWscjZlvY0aBZN+9uoZbAT0ZOf
FQwU/WQ2vUSIHhIXKvB7whvakvVtyGVS1rgJQqvZsQyjYUOOqieMiSvw6bUUAWHmTdoFtEoLMrXR
EDSfzJdPYyEYU+aSCaxI7fqDyBAtOe8q95bRZBv5wxYg2QhGr8/XuEL+JscHRfjfDKfKD3xUx15b
A5a9OjfQQDSrkuzRue+EgBL+R1MWahWa52TSizZgMbOB1iF/YViYAKm4CNpoAgBlOjsDNz6UPHyq
rMnInLGIwa+blCwdls5f+NBlC0NIIZXaQzhTvFGRnOZGa7JRVu/hhtgQhRpIj+1sQU2p2AJuZ79l
AYBJVAYxN547+1y7dvXWsvVS7OcSE9VbXAbJZMwHj6BFZrSOD8pRQhfjbNUjY50sFj2ysxDpzXth
04TXf/nTTx2qbgTtnNsOkRxt51aj2F1PHmo/Wl+b61yZoGo5+dKobyE2YP8AoeU8lH3F0vwyjH37
PoH5yvp/gOhkYv7ny6sIbpXSQ8ufd6xkEJ48mhCEAAdNwyTwB55fnUg4DZXZZJ91WK0pYYtYzvW4
kAuvDMir5Hp7pve8fgmsTY0yJBwOuAmqAgOW5I7XBliH+ERhXj9tk0yjaXjVaP4zd/oBb/J2dE4R
/dej7Qk1/B9036Ibfh9RSBucVx9H0zE+zk9EOudZTZxgCMJKe7hskYRruuUvr8fMeIfqNfOjMp3a
hyRr9YtXSnILgfzE6aBUmrcQFPOH5hynZXy8GoHIX+RLzeHl0Zcv60YI1fxTm495wk0fQYOtHpll
Wsq52WAK7maUtE9C+FFTEpLyPymQH7ghFEwkqU8bxonrtbUOMyXOToIQNmfLAwwNj6p2cUAMb9AC
alCkQB9yzDWbgjX144rFTw5lSB1VJt1cxUMAnHspE385zwmLVqFaRMKoXdcHutZmptM5O9UuMlj/
b7EPITotlwZyL93MphLSPQHSD8giNXYvRJiv6nqACr3Hx+G1gahE9/CavkECZ1Mu6whojslfO/P8
GUg34uptg+UJlgROjeA/Bau0kEEm5ydD3wR1DQsAXLcCDte9rF/R44KmVkUTcOIKAoSo5Zn41pvL
X62FAVex//yKcFB2fz4E5eUNPPzKQY8OBCxAYjGtwWsliPM5iFgb2eTZUNrMdpJa/frc99/efrYL
NYMOVmNlIP1pkgnGvC5ER2xE0cOLkxRMyzum9kCTpqIz2Yb1OV4vhteZakkY1udmrdb4x7qzBQhb
MYgaDwi3Vy9U6Z6rYzaNgGj0lNHh7shDsWmr02Hqi4sJ1uko+PIwk/Co4MJxNViN6t31EvZpUM3G
y/onBoxeFqIANezQnfdr4tsoYcjpN/uMHpAjL6T8Xe/Y0XzRou+H5ZqW0DYnqDgt97PSfhrToGLe
Vd5EdthnrTclXKPZ3Rgkj2MHZNh2lDENbK2Xf6zgzQw/GsgrVbCBqxMInMHj9QVIj846sh0tpR5l
qOtHiZpI4PW/WyHb1yao0kYV7pi1DzuO91dZFjqLgqA/IYRZHoWYelweLimfM5QiJuH3EBbVSBeU
X9lc2wOBXdlqSHBzyUE4I+UhPYud0KL696egi+hgRgbXzBPSexu3eF94rX7krypKfP/o8OFUE3HP
zDcVa44Kp9b93QjXJMmYnPI57ptRqT0I/CHCkzd2aS4c4sA2SBf/dxYVvcCxefpfkanCJzfLWIK4
h6pK+ufcMcH+hNGfeJPLHPg3sHIvjdzXrRyJXNV78JP9ZJXsnvgQDB5limMipkGgha/QGaCjgMg8
+GS5DLwcqneTO81iZt4KzrtBNOOEyzuddTel34MjdayK9D51OdvazwLxtf2EqASLlXWRh9kQmXGV
A4TxE1vZGO9H1RPRUMUtq5io2iewnXStHTOH07VxLn01SMDywJGEGT4GFZGX/GQFrL/u9SSHOWHz
J22WgZLrzaAi5WTYcuiDtGFVTKGRNJF+uelh/Sm6TJwZUWEtn003xLzqWN4eP+oIusdLXZXEZYfd
bO84Oxs8TdbJn35PRUCAup830mIHlPxYUcp/JJsWL7Zbq6VQUlgsiX0u3aDvXIavTNuzZdg9uYsk
1fDAKEByeZNKtDbHynnXaClfootTA/5GDEy9AaSX0HFTqzWpYJUnaLGd2WWENeGinqxiXN4fVqrv
cTz77ToL2U3tYv8jkIpXwb9cLNGj43qzGfmDWD8iFMd84E0ErXirriE3VrKG3/CbpJflUW5V0o6c
xwQ3Ed+UJ9RAbo4NlNf4/JrZMNBqnU+Bear6XR/snpEVyi3/iNDSemXDKNzgc2toax+9yHZ11KAW
mPuKaJ3LUuN+/rrkif1ycmgObOt+OXKJyVDfSzvOupQZeK77JUVO/N+7Dl8lrByZ8JovUN7lsMiB
iSazr7Dm/XMX6xjSULFzz0+c78zvZpepo9AfAPHSuoPeXRLcaOSuwgrPvQDuhFJmKoY4ukt6BaLJ
XklCWriM2QlURCTIrKEKKbk7PZOYuUAxqJ0ReUtStYCAbeURANa5hPG9oTsAhNL1TPLRnPiV4r9s
qbQq0DzOmi36VLNXaGRAlCF5pKcsOVlGt69WFUoh0kUuW0xToRjq4/k0MpAfyxsGuJFOydnNDx11
iZH1/bNc3CCakQOrNfamm7WJg84TsMbuQcNmJQk30bbLaOezvp3rtk31w5n2WEknI2/hr+ZaPzxY
XPio9xDSwEHtK4Hbo1f1AVbs7YoBG9kzKdVYz4t+QwDcN8XbIOgNKKvmPk3CC3v/n3fKgDq+pDS5
wdJDAc3TLVAMjn3qya1/FaiHsNZL09Sh2+4qKIIE7dPyGOi7NtWCyyfRJxSm74WXeYfj22UnIUwX
081DRcyVOCvEU5i/6KON2fHhY84jWbZbzyBQPzfA+c58DOgds7ajV8rPA7tTSD7pp4PDmTX/XLhi
gQUx76CnLsK357TkTidHqX0mBycqq8ltMMPgqMIrmVOz0zlT8U7ydM0YSo7CvuyKCg04FufO+I+/
UfRXMkxht7tnzagyNH0Dt6/azhm6k7b+YL7IdPohUCHvE4fgraOH+/wq0ItiHgkC4fO5dLWkQC4d
eDfX/5Jq4xRdxnNMr4BIMQuguQoZB2iKTiYC5AfoNt1/lO8RukPfnMKj7Kl8+MIhpuv+EbwvTa8g
Xw+3cY7dX8hNr8LeIQ9M5eOOJGAFEXtQ6P5K78M5qI+6+P/C6VI0ffep2JOpCOGvid70XJFuduzH
MYcEGGWhp2rgt4vSCiTS2ktStpJnY9Kg6KjtXOwfyVnzPSJAdRl/h6bjIY2ehlHxT8i7SiUXv0Y3
4rdiNMZmwJ2LHYe1ASyYHPiQRsWCg/DZg+Xa0/O+rJi23JFt22KKkbnSQLNZI450tTUg9suKBjq8
Ut/VyeEbsPTrfgAWewgI8jd86r7+KUSEC1fm2gNZspHCKMcS+aJzjcmFyr9GVJZTIaCEfsQU/GSd
SsszO7Y9M2gLuIXzfMzEU02D/bMdsZAf0L48PN0r3tnVXFr7t9FKzmlNsAzGVjwHh+dOOMXjUADq
sTWyHNNZ37UBYfx7KMf8UwDcNiHLEmjWkEmIZN6NkzLIW4AAJoEAnbKufaibJs21JYnziY5Hyx0o
2VxhMmIOciMQ0Rg3nqz/DuvpNoa3WvmqAMa1CTdG517ya8yHN2sijzZO4qBQ6AbreskGrPvduz0e
QT3Ofe1uejuZ3oTtkj2UcLDD/+Y8cqXZbBAkYpI7FF21gmS1hDeiBOys5aXZdZaQqfW1i8dX/Yak
b9tCvyU31qAYugsOrpYwK8/dCLa2Y+vu+uLT7hQhaqAQ7OqMe7AXhntNGnKyzwA3s/pUOF9bNeaQ
Ctk/rbzKRiJ2CkXyciHRI7LeGsWunpckb6gjNq/zXT4oOz/6hkjzyHdcR3Ey4fitWKXMQudSsEQe
g4MgaRMz0BgifxE7DsRHMBT+E7aGZNoJkK28mbzIWCR3VPK+usrLfm30NwR2CUIdIcIFn82T6m2c
NNFXI+WY0GzKgSVn2v6IW5uovCOIBUy6bedtOcMvCPBljvLRWtXnJdc6zPmUJvUWlyn8D/PFNKe3
qjDkYp7NNHC33KorwIlU5w41YQVSZtzRnrHnHInyVUHHzjB4/ihinUuYrHQfpMtFLao07Ludr45e
bhaosVMLfhK+j/X5UpTB3pKYnnyrvInbSfr8d5MIFG/meBeGAGQbfCWdQAh1kriYKBu8ZU2DoZEl
ZyfPQHAHpKDnwNOTBWM8CZ0sGDF5Rndio7U4qVq+XbAIwOvGWEhq5ooIUTYm8isJKWVdPItx+QdB
ZWoKzA5KCjl4VUWNfq0vpccotkZ4ojc8F40YpyEIe4T3ALH6CeqJKTiIKzrMEaLCq5Qng8GC+OBr
4XrjYMDrok+53v4cAxBjWRoK/BXZDaxn0i/7qny9BYB8xVfThmv4LA5EhWSEV+OVLBQ8Awkva1Jh
QllMoJn5OauiKbqLY5NAGky+4jhSxQE0kAal0I+JYkKF8bsRl8Ggd8HfD9HlPIeRCARl1pnPe8Gw
GECo3nww92F31eBhEHMRaK/PbN3MywBYgxPZuowDksi4j3BfuQvE+ULC+cJQv2qqaJyLDeEbuzEb
QCKmR3gTTtOfWEtcxppYuJFg+JKQdlQIEJEhHwu8GUKxrzpUUZWCkfA0dFx7nD8L957x3Rt9+c4H
OdWY9bJ/GPLKuPQ62L2G7Qr0vZrzYwE149M1x9N8WHflwUMmn9yvkcf/miZEobT73RIhwbw01ryn
PlTropq774XVIJ3HzuDOH85jMUWQLE7VwtjJ3Boh1VSR88W8TWqgNNpyDUaj9rsregiNb/SaHmFN
HIUsmOjCYiuOajS00Y0xBji3KRUU1JDodwDRRbbY/rPDocwEREXcMQSTZ09v/nnCyoSfMFS6ahqX
wSk38U5gkP49fFrN6LL7qrWbQrxO2C0cRpC5Vj0jNNnL+YUBg6kJl0QfIV1bmOZ4KEDo3/oekYH7
Wp+LK5r8ocXG7J5O3CFiUtDq8XQX1fUyHBP0gZRFNpalIeHKdqvzphepps88Lxpg2HTl+S+fdfvv
ItbxQMacpIfyYSLEUPAN8Vy2Wyc5tZNYxrCs9jKIqZbSukVk9wvYxJSg5ctLzAOXId7F3SXtyV6d
e9CdAqDkWJjDLk95l4l9QJH3xgRjCxqEjhVJvWnOY9Ovim10V/wK4o2DGrb/pfmfDbJuhJISiU2k
oFECNiDiB3qbeHPDbQtNhpnlSe1CnUYb2iCefhOXZgBycPwb5I3s5UIk8M0aJORIA1vgAk3iF2xT
LF+A8yzY0tyiURBo+6w832e2PXhgyXlwzZLnX9DQSOQG1LIrZHCGdh1RBHc9oXhjBovukKt3RORF
cXrUrljleniRf3cACL/qKnCFKn7u9f06WIzCd7g/51JW1LdF813LKSVWvJwbHc+MiwyHz4I7X/zL
tLS1UOrrLjIRXDSj9IuHzVs5TKeb0sMhr2k2K4AlNUV+89PCuz8K2XEgvnX43L68uQwuTL+LY3XP
pd2BKG6TGaatjPrkKX+9B5+k4/nhS9xOT7o5Dx6ilyogUHc+B7n6QSMGCXn//fzB0970dPQ4C4Mk
wYX7/xc8T3t1UQNuCfSI2B/rJqvICYwgcsTWXTumqo0l11sQ52FuN7wJ81eieTuXg44pl47PbuVM
LFm1lbHTRRWaetY8TWqh6wdx2X73X0doSYm2Co8+nTBlAjZRl081Z791Cr0YLuINMxMh+eN4h/JD
51Y6xNOkv+JJE/MYvINd46YHlSCkV3oKwOlQjkZHGc2b1d77q6EzAWosNJ8S7QbvP2RMxhstr8zz
BWqfK1SFVlkZbh9gCCJm9l6PRm/nOOmjYI2KAlnYTBIOp4OCZeJlORUqcB/eeZwb2DlGIK9pKk+P
b+zS2BL2EFi+XmM+mplxwbk3pOkZ9PGO9Zvrp2GBGwFfl9+cjDK9XFhs8pytp7Id3Lq/U7ZUlYrA
vVK9FodjnNGBWhOr21kqZ1u5M+HXAmQrkoI/mz5cqMG5hOKBJR94WY0HaMGXLX0h8RWkP8hG29aV
vLRQuXk3Y9c3ywA7ekoWKFQ+lghUDJ+sMa6pT97Z0+stmmVetoGodYGl271tYzE5AKGhrtXMlVSK
SG7x+rjar/hcwehluvbOKMARGMo6jv/KDAr+w3p9bw0Q2eJgIJDsHlGRSTpxvlfh2hNybgevgCD0
GVDQwGEgXBBWAhrVl8My9n9w7Sn3oJwBkfukTIEHv297SI5huQm/6/Q76vi1xKQjugLSF92Y8Omo
RMUWjDMqJYm0SFzMt3xMD3q+XP49yqQM9Thtgf6AhYp2093Xxn5c98YO7V1faWSWyIKmE4Z1TD/x
nQpjf5pJ9NcxLDzeCjru0+E+ImK6LnCNU7p2229/rtO87BY2HB0utbb1Cnj8fbeYVJYKTVOxNn6I
DHrBK3T4M+AF1aiSPNSM2dRz52wVkyFTsPFtDUccESO6fERCh36Hbl/CQjSvCRl2ZBTR4tWr1rDx
efwTOfluSBgWW+6tESb5nLDu/woRVT/fik8p4iub194n69GFiKXIt3ceKOzxKne1yK8VSy6OHE9J
fnQNvD5QHprF54FHyuULQGITA7AfZPElD8NRV5Bjk+4LaL9t7l7SQbKbxvA3g57fM20K7M2KBOOK
dMHg4+pDtlhOgi067cWR34ISRubKehEW+ofqonGRQwSVsRUr1w/KLM5fW0lg+OD0QR1FlyISQRuf
5ompuYtg9fogpHdtslu5n6pjA0xG7DZVe9xkc+5plqzbpsqVYlqa5FqrCduY8jdjgxDGLMzA23/X
2nRWLyHQq3+gz/rtt/QmjsCrXa95XDi5vRp4HiY3Um0VgLiRG7aUUuBhWsiO+sgnTANkm7f75hpw
ohVWIFOIoLE4OzacwSJfuuLv2/I8Tz1iBh1aOuyorcH0HDfIoIXe/PWmoi+yz49h9evCqUcYgT5d
8pv8jEKHFIYQUm6PPbqkP9SSToVMMvsCoXeR4HeZaO3w1xlZ8n4d2GwQJDekE1EUAcB2CwLgddoH
LnWR3Qj7LzergkLrOPxeztE1PspJciggNRh8rM6k+U+roZpoazt9409JUiE7TRIxH4qJe39dULqL
2bRFR/21/Rh0fhbTA7xn7NGC+Ck8nvp3csIlgwiKlKhILYnkFiGier/FmdLq731fAqbVTZVExnNa
3j0Ra8SaozQwD5C3y0ikztzQWEtOmHOTzbl3NJ9y+bTLjvjuv18F76RiTnyUQfwM/qHq4Ze3a+JQ
HoROwCCdJxgiELj5KIYodlDi8suC6/2yEUV1OsCpL4AP7nwUy3uE97nCgbuDEBlk+QBl74o655Kc
Jc/scfzlHFGfamnpdaQTZGFqB4g6yLcy8OR7ME2nKrjIi68ZrXSOhUglC+z2752i9SUBtAZRbCdS
fnKt5Ytcb5xRAflO9Sb8Q+Vg2goIPDjt41REUPttyQvdy646INyyMRxg+xGToGJmdE+4zXdrIvCr
SZm4cToh9747YAeXL7UtUVqqfcfM5fWnZ9NLiWsfy7SB99pLzPIF11PQAUCl2M9SyC5OQbKBQpQc
eA0CfbxLt47gx2rAslQ/wx6AuDV3trR41CpHNi7DOUwqweJFJRwlO01TsblnGRBvABTccTSRIiLO
PQY0VI7mGzpOoSEcx9KPkEvLG2hqy4rorM9NH1sExfiDoW3iHlYPYIuHdYu/FX/nqrgLP4mnPW2c
SLDYv2odsvXqqzfRMdAQwnPtRz6kU7VlCWwn8YNbNfXN6Kz/RoInYDqQVetFZ+vvFVNdHybrza3/
dt8q0dwMwklqfouYxSxWt56kQuPk5ih2lSkifRWMq8zW4zTavo3xyQXzJBY8wdm3GHvo08zDLhft
f8PkQDimdrZR16gTzIE1zQPc2vIu27B9OVmsa5rviN39kmik4v+VPWchRRqNuB5xs9nImuK2br1E
CheGwZhjEwHuJ1U2AlyNe6GwLBbu4JAdw2QwoRv3RvFf7vDkjtQB8Uj5KVyMhcMCOZ94/EKwz/3E
p+7k7JGQyJS4GPyH2n5JqarjO+ZccVQY/BfruXdO7527zkM0QfunsSzNyvtw6R3woB37rjRsPi0N
wcCDlzc3cYNGIjb9fvvIGv+nNP5FmldhSdHNWhCWrCCzNrC1Hr8myjBenPEx6OP7EDgZWybh/FYX
HUwPdn80aE3/bV6V7YAktaAFHV2NWQWMX6dh2jMNrbUhNJZIops13ZovIE+eyu6Poc1ll8numzBR
r/q3wLEY16f8WPkCG7zQh/ycTr22Wko0Kv61win1nR6D6qRZkxWEHEBs8b4GwjY9OS4PlUc93KyE
M7CSsjC5r4IOuf+SYexWDZ80jxMiCyFgk2cvFl0On7FRnhIGLnis4QHTvWKbXTCaxb0LXOVpYmET
Ix+Xm0CZDzyCNViiDaaFRSaZP1NzCjgfZiaA1X1JhK1T1VEWkCtPRVbShaMXg59Ts527H+g67kY6
n9st0A+Sh/isFBijamxRdBF8IaylT3HOOM1gj+Cn4Su9GI1kpDx3jGSNLfFN6WCV+nTolo0AEzVx
zUH+aeYmygj2NqVFtHnKmDwmETHU4jWtN8Tq6pPpP5K8Vn7aaqv5RqgBOlcmR82CDxKSb/bDMOR5
uy/auQlokJLRBuNa0pWmgTQc5hzRS0/Fwsu20oRzDLZdzAgItJ1YenAfsnIb5ZU0c2S9uvsebrJh
Od2024JSk6THwh4bonH5k0AX/9up4R6nYLBZB5cExGms+TvO5mZRICqV4g7N6KU/LbojdkEXiziT
t76k6VQ7CaNC+hBcpZqCtlUwXSo3VV3jhCG4PJ4Nqb/VM4Jb6vQ4MvMnvzW7KO06HjwOpak0pyrU
iQ1pnhB279obMqNX7RYh4DQuaXvEm+1k0yrti91YlQ5/kzdQlTJor9/SMQRx8Xw4QFnC6PHKihXn
kq2fxXKIQvFV0f/HWztNdJzqw1N18k8vYh/1/QVxjsqRsuipRxiSs43oHelHjy4xP+lxCkpKLJbw
9ZsenEw6DKrFGJ53hfZw8ez9yP4weFvSznzXFVdKOrA0/oQGe6qM1WjFu2ugyONcO6N/t4BLQB+Y
k/ktcTE2fR81KCm0GIY+89SdgItfRHZsSmWCrovpdLGvI0DzooDTBwNxXng0AUvNaeOj5lQDjfRl
QpOA5bR2MyJxkkMepCXdCy7OTVVq44iyRgVO/p7NEV7YjKDDk44AP8lgu4imON9pKCVOWBb4zoDo
ePPJdYIRv8yhl8g/ZfRQkuponUpC0T9IT1LpWWTUXM5xxNxCzZ+PRN7NLkVe90sYV7OfZBbMW+3q
XkRBSvPoaROUmPq0VYx3cHR0uYXifa2BOAIXD+PtiURSzhQxdYmBHnYLuNatNwgEp2qFA/CD28LF
CXEroatGLStD8yBTYb9fmASkhJ5Q+z4UeoNzilJYcgFVFfj/nVMZcy6NXBucSreiRKJPPHu+MRYe
56JLjkK5cCpHT7xR5Q6c43JNAKZv+eTMhGl5B64l9jLee1Op/jMdaNtBxm+jrnU44RXGS2MdOaWG
WNP8VoHwn4QZ9yRi1CJk78ns0XxXojzKCAVSmWQ6iaWHvIR7mJWowRTWOnE6yiv2RdZSo04IwnJs
WGg/IIE+u8dNiLZAfabCthQuE02pXtZ/6sKoH0ehx7MUbnNXj/zoeVcZY+iVOU7GyWXaFEqfalXf
6DFsrOZXxLm2hoSptS45wWd4vA9izOAOrB1cfhj1jr+Yw8WCXNcl8ti+qV5R2tTb4hmiEFbNiw4O
bvKvnjwxzM3I9HlsgU5fNzLGEdaf9UvsMjFJegaw63pwSr5EV8GsAVU7COna7RFQNc3Ug2cYX16Y
Pbleb1Vkmzg3gyLsJEurtpbhmeceeapfbb30Si6YBZNYGRFS3O6fQ2cTOx33ebYr2xcC1+OXlCOO
EVZVICya0RsVOM590VcUKIk3SLCQePhs5N2mHfA0zOpGJO8IUPXgAd/2xRxFJu5ANpQCEfZyxdMC
uultIWrspjktIWBH0nmqLREM3G8jntfT65LmtcLNGFC6+UwByyR0l6LV0J9N5nIzMMzQ/+1ljVZa
GbtS460fhVU2CqZ+S9g4oGqLfZkEPvL3l3x7xNint+glJajKFJqbPTdepJBfVH9orEFcGBqHnxLX
+bxM5oBpCxgjlQTSb9G1qVEOZaap+jWE295IqP6BzbQKQSEQubmI5/Ij544EBCpBH1F6L73dCnhZ
e1DCeNX4/UvPYZePU0xH7TaL91qopwIiX6YAgRmlSQUDCmluDYIFUbz98sNnQ79k4GNUpiKlaawz
6ZuA6lxNpPr0n35VYkj5SAdcbB8NoxbWsY4K/qUt1d3uI0EfxsQ8iieXEQokd+undu/Sp5ojVTI4
Q+3+Pq1KPJWfnIhdxb3k53D7M7qg7H6XTWKS8tbGv24/qGQN8nz4xM8tflF0D+kZUYOkEHKqWVO5
T0ndDwqjCt+pfX27nvypZiIaKWNlgrlHjedH60zQrcal8J5klf710ke0wNj0LhUy8IGYt6PTWHOx
80DLoiiq8KYsFE091nN+MBJkblyI3wS+fUj9x46bCb3lTRTiuXV7+okGycdkuP7cYkXqOpQCEpZH
Q2VciBFH+tOig15ad8WI4us6luFXDFAhWenXm+ZJpLoH1Z7eNnC2o5u7aG7vbywJcHXoL3sUYPHl
2VwFlsGhayHkz7z1AV4Y9tIZL6ZyOHhQvs0QBv9l7raXRliTm+uE7cYpk4MtfhPupg9uNm6ZiMO9
LvObXnMnemqmgzls6zwnwTI1SzifBTdw+4qgVcMyat2Q2UCZzNWhRm0IH9oQCsAK9EjaMbgvYT8I
NmSyPTXR8Gd+olHDHCoX10Drer+J4pZjj0rBJdPFY5LWr79GPShyOHCNlDv4QL44sOx0khHc9cuB
gcJQ8wZOICg4y2QQMRbAXdoEXMOo4Fg+epNoeBbWmP7YRyBmITIqQ6eBcfp29dY8kfsR6I6fxNnA
sAM36/ljSPhf+oGA6Jipyig2IayQ/ZiTt7D4wXF9t9+WXrCy0OLWVvm3SNrGk4OR8ey7y4TFZnI9
/Hzn84S8i1trlr0P2AF6DS2w4FEzy5rpD6fIkpmj11wpD6ByDIwDv8slpC0d7eI7WKLSrmbpalVI
oA/Qt1Gux61yo85EI4g5Rk31vC0KKOIgee5okC9we7wkdr5v13ZbHgu/Kxv0s+vGkqP2/pXn6s/y
Ok3ev0/zrMZoGP/OhWwKAZHg/7v3hK7b/fo/2cPZi+/W3sXzId5mF9X3cdZSIOxFhUuSRTMiEOll
g1aNlpiQQ2cFRhyLhJ4rj13vhSKGcX2EpXK81Aojbr4iEBNwl1OiLWOumaDt4Jiz9LLr/TOeBani
S0Z/B4hfx91lItlDO2uPbIHEZ7Qju/imeY8Fo+NP7Yqtlp52MhJ/+lpwYHYCc3FH5vCA4ynn/bp1
7gUdpvwzjwv837lUanTK7SqqVmOrXVFsV2GwDQqBmYut2asogursUVEhTnG0TDlLqdezILOy3Jry
akajkmsASqAIN5nWEYvrOdr6iBmcyvCtOVF9qzHuPj3g3ryXr+KRi4w7wM5Yd5E6YJVPjiICG3P8
28RXEnJUf2+/7vTmRWYJNltLv/DQ7mFiz0qtPCg/dCf8jPnJIoQ4wZBpAIiXe6FguMjY2hxPcQeD
SbPMGrPHA5ZVtHS5AjObb4VzNgVt6XjgnpbZ6I2En+loI1iQtjUoM/OlPt0TgVUSI99n0SOjedj+
TE2BcwxEaFb0N1S1STlye3EQqFG7iodAZr8xXAKb/5q3tZNl/4xiQmNATHCF1Uwc4W0hrrMlYvWo
LlMzp55VQ5wao1E3eYHJAwbL/nkXAsImY5OYLiFVH9iW13sxA9erGBbgc80af5TDnNWy8xDbWuCJ
JSofZjyM/5/5uFmY4Ukd4CsEFS1kXIblcy/VafJwvk3dzN+VtoV9m/RLP1t7BOZDGG5QMQ2UWNAE
+9kBgxvk7JdZeKNFt90kh9wz8CqkWFnILgNx4PffUla35lvoe13zWgvO8LlNPSm5OrbWpEhkOY83
an6rmuiTNB2r+vqctDw4nF6mMy413+FPQJCYLXO/f4SCmiJH2H1Mxvoq8tinlBEr2MSARy93GyGB
WcQOEvgefM/9NaNfzC02+KL3itP/3792QcQ7pAqXn7Ed/AY+QUarIVYn2u4So7DF6M/5Zk0fvidg
dYLd6zRwWEzHq014ZtuFm3Jwz3Gskb8bQ2mD/ccOAzrbikftncHYNQlDtOFdue9qOs2z6HdvFuOU
+r9CjV/5ergeFSIirsAmWJiq9skVKojFK+1mTtYRcJfU4ATl54sxJ2egY+WAdPunefoiXNPv54/C
lxOz6z512fsPsahURlZKePk+2aWVOQaUJMOGnWFzOxfcxGOXJ7gVrNi/6NwHomiBGQTir1WaRHRA
f6JbVzFf00L+ux88VlooShdo9/WxYseVMxSHX3z4HLbPhBMwZmRG2N2/+vXgpWCikHTQiLUdlv7z
pEMYKNxNB8N9vW4V94B396qMd/ji36n/1/ya4cNv+10qKuUeZQAg+qKzBF2kQFMLneFo/DUiZYGl
grbmTI5MYiGT/DrqYXfpBCPdRGlL8+ykxeBfaPcFJfYYAY+6WI1piOoQXuwB/DdyM7zeChP6t97y
NXU93S458nw4hNH0w8bexjFgsGI+hn9IcvQX3gWG6iZl9RO89ugnbvEg/9yVGpRZNeFgv3S6WLfA
6NcitTSctMPlVaWAIFWL5aF+i1G0QpYEAvGMWGtjbJB7r7cnd7L9MN0OBcKvcDoII1ocrTP5onf4
5G/0qp4D5jdzd5IXf9yaD+BzTa/0H4eH94+9M1rqeJIf+MIMLkV9YOENffo3R2ADsJFl6tPN3jGH
0aZQdU86phz534Naewvs8vLzTaRFTAKFf0UJrlDh11SWdc2IRztIFD+0C4cIpIrd998LrvLAN0fJ
ApdhaG8/r0PoK96K4TsOdOORSxo1ZL6EEwZdAQOO9e2K7duowmnLf6PIwwZosjV5Bmc5t1hGiN75
OlO6cyd1QfhIySzz1f9qZjduUoOXAdrIWR/ZUT7ByUf570nYE+2qLHYWXMAfH3g/V5cWuh2V07m8
eIb+XQVJF65FxoFcbBN56OQZ7T3To8FDPCJJ/y+DHKSnQAcbHYT1nuEVn1giPY9t/YVDsUNkkwfm
LnBnhdfPjkndgblGke/kLTGefinQgp51G02x0pcOsymp+CFQgUL9Ux6sOFG7YjLLXivTesX+7Kmt
ICWg+qn23BjaivVwrkUVnD63hEO9p0YNeVvhYY9O+FrSg5APXNKdCT6ok+addIGb+GI1NtMOqAmk
2KdtjourwAybu0lw2w7gGMG3Wj7cdiRSs/qrYfyCMNBb86wqF7kbAWqqxpl5T+DjJ8rDIvakDQGD
T9PTuVOhvWnSif4j28SikuIKtTk82eS8wTAootqPIwfOkyPxPseIqqGwRXsRbppLJr/cHv7vVC6g
YLpR/KMQcDee+g2TXuQlzpHsHXwNRXPiA/rtaS7dz7yIJDNGRh/NmMk43qnTYda53jNYwmpvuGQ4
Q4/q+6MMVNkTipdQ/NYhPJJqgjE9JO7BA5vHcqX3OQ2HO6VYnEdrFWjiBzBiI++qllgOIG9ERq/f
CeSTHi20IPfIx6Yb+sX7oWgEB7EDajgYgY8cd0V1NybkAOr6kS8plc7eMljGCaGu12O1b/2QTr6I
eIBIHAO+d2jW+v8RdqV1VV0okZod8wSfHY2bAE3z4yk+LVU2mm2xggg6Gr2kcE3f3JAR18KKiub8
CSFUiF4Xr8gff+QY8PaXq3JYRtFeZDZAXoT+s4Rebi3N8jpS4XpXmse8Wq2FFBeFUnizKactlAFr
k1/v5iH3irgBLzTND52tCxC5AnqSTkOvOVl1NDIbak1q10KmU2afjQEEbv3CP9+6fAiQQyileEpi
pPcK/SoGsm19IdVTBPeXnRj9P/G19IpPyLF0D6/2IvGjxxgNSjoNSwrPbCHhafHWesKbRwTb9kP/
2zHt+6Qn2Kz6cd9fEYamPd6iA+oe9aukFJVdQ1hb10yEG0BOE2+vgGDITNa5ez4UU9U4gSgE8ZAJ
/bBsPvNCnGmo0hL9iRC7ElM17q78AyqlC923PderhN1qO/L39+/+pZjghRnHxFUqVs6SJSuRlyv+
wKdvmOW1kOnJv7Qo+I8o5WN72bNUoos/UtR8yB78T0JzcusNURE1Ye67/ZvEYYX2Z+qID9yAp8C2
hBfYXOZKD9PEcpUf87B9lTcZXh7qjqnsjBCXFJz7bx9mXIrW2ATS1QjeWcFEGmHz2c3FTQTotqRb
BtBRyjX0kAsamYGrbpI13cwqjNWP6y+J3CrSooCVDrZxZ72JTe0jjiYOdW/tMGfzlGQcJbSXXZgl
Qdqa0wSP/51TK/TlX9z24rOxxEoYpvwSZGfChZIf1KrVSknTD8GviV2OzUDM2gwQ+jwmhSS0lNUN
NeLAMZS7DRZV9U+itbYdZI1HQTBZNxEadcaslgK3N5ITPNKDCQH87HeX6irij3zB26aYbIZuXmrm
Ter2u/AIEnypr8DeT5UpcEXtJoyFjPW0yzAlPacg9cX6tGFyZc1uj/Dxg+PXZJvjjPY6pwmHq6Y6
NbbFmRRAMTNqDyzMeTD9NmuNp68bWDZ5mKTKqbVN2AieZR8R2DQqezC0a4bgJmepqiz7IrB2iOoW
z9Slfet9SCW7u3NyxQ15Nhs5Onqlgl9MizIW8fbhOBoP7qTjacysQUUtdIpCwtg8aj9/qeKtbN3H
NhaQbCuxetzFq7gYmUbRwElzQgxmx8ViWBPZpa06vSGuDrYqLe3WbGr5TGJ9SyQPFuLMBsNOyJL+
7P2QiBYhgXqPjKwks06Lml0EC0yFVsc6yZvF2hDxP7Hi4ZeNbe/PI9bWtghCAJLE+LDhWAvzrXPs
i7pT4VgS7j/EndRlRhGDkOme7BBeVPwX92r3FaTlcEd+lHIvClO5Ub2t9IaoillBsvfwXYU8/X0m
8yI2y0gwC6xMifDDKsoG4XGHrvsjp3+S49utHd3hyIxHy/53k3gPzQdQrssayACdg/zk/pT52rwU
sjRPfME7PRDO6jvnsFo0vLnpAornqu9Sp8KM5xFM56FCpsaIm0wqKQY6se898BLiMWpkImspQ/fU
8jPjdnq95qHlkRQ+7gAQR8ZXxql4U72mH3bPfD1dOnlZYLB8wCkNdb7Ms1FxnV/IYOmkUwG35MBe
fKg1dDW1KSqbxpmgOsy+QE7FaSJDv+iJb6o54dmQvStC/7naJEXuK6viIT31jnOaeUBb65OkrR6p
APmbjbM/tcs6uboMmk3Ru7vyR3q01xh2jhye//WrbVuXqIAWf4qNOsjYRfTMBDy3/WgQCktviQfB
R/YQZf/9W9cKSP7iaR3z/UwE93ik8QuIre27uFpZmwm6Y2lD+YcwqXdeJSTQmVEJon1KLQ0tqvfU
n27oACiD0od17J3V3QsbCLWebm8770eD/Th/LSJMevc5Mtb+YcpYxHKdf2tBuSdwXkJrU0Z/SIH+
GT+1FWzwMr4PycfptLvzc7QstqZcBocfVXIcAqHXLGPPJ/PUmhyTizpRRCG7uYagL3nraQzbOAMZ
ddpxtiSz6hR35n0UsXAZgODWX590B03n0720oAacaDP8JRi13A3HsHSPJ2W7KHXCzRkvJBHgqNol
tebRnf1Api1tel/jueh+0cvOAftZvJaFK69qUS2n9DVr19tJmb+wU5EVj2j1PjPNfKkvkBgv/9o3
7qlO+zJ7iDEsCPb5Gm4oN3yH11966GoLE2hI34fcxbSttswL5gCLPM6pKudJDR78wYwpqqQaWNHq
tdGJWGUgtXb0yVI7UoyrraSP+bJtI+cuyU1ao+8djCIIaDMj59crYvg1aTGez/r/OaDDhN6ppypP
2zAMbBfh59q43K3arLN2mfopZEak74oMMbKh4HRdc5FkiunrJauAKVIQxcyYGMFUg0d1bzWTL35G
H3mNipkWX+VcrGivCN/CBcnYBhl/Cl+sptHg9CEiziGnxAcLWzctu2iR+9vtfETFJcqHBJX8Rdnh
DJkmSeo9Jq1VPBuUYq9Z5/m6AbTF/aPxwZHEIsr8/X1pl7Bpn1EvxVcp7zA3UDSXMFXftbeOqA0A
0qyzybTIUadgYN0exxCC89QdSWgvVh84K6DbUd4HsC5VbSo9dLeFq/QjZdotVXB6xaYu0/MWORpA
mLXwKaLISUEqvnBuMadE2X+IppNwWXEWClVG0jVlI/8P9rRr01kVP7lqU0U1Zh+YLwQgD/kORtoZ
40nHX4Gt+WWh3LSzVif2prEdRsITgg2/LKRqdjr5h4CvRla5vYKonZL6eUugUckYoMDhOFiUuxoG
rqkESaGeZEx72d0u7qGETiV8PaQAZC60ZksFzj/gtVF3IQB5385AN3eRyRt0rBnNSD1EVvCg+Jgp
rBXDwCRxw88qMw3C6Z9SIxoInymi6EiEGajnBSXZ8BFR39b44zdjVFWYbKIJb9ouOTJb6tCDe49f
pMOmYw509UYNJvR1nqWrjbfJPWkmyT2WFiMGF3Tv/zqXVdl641P6EEEzH0aoXWC0YuFb6Y8vHpzJ
yVo+czS4qrRLtp2ABvjDZ/iZyuuise7KWKPgA0igriiCvZFjXTs/XM9XgHqOg/W53chC5KAZm/O/
F49lOxkYnAM3wCRLJRvmfw0xyhbMxS5W6vpfuFcDjmtbbi1b/Uqew2itNZwQRrRHxzp3+oeLG5lK
CqtdVLEoEbDYVyhr2YUwF9BLI8SqSIGVk4LZUwQt2GOiWrQUkMhMDCNwTvrCGDaSpVeN6UZUmfGX
wUBkblkpp/aBj0mbr0lDOqterEpqyYJJEgsvaI2/Z5ZswCIFjYYYlqKaqbwgV7asFfxXfb6eavpp
DLR4GhzJ1WyAs+Aq2vPdb5l2IU1u0Tiq1gQppTtNwg26zjoGAxlQQRIiqTHj4f/tpBJR5Rh5w/t7
2f9zcMOhu56+u2c676PGCJG1m5sRD1mMDU/XTS7Q/YxciYs8tETR+6o4up8/6LJVsiu2D8wh+kxY
PX1uqRq7ETSxVE+4ZoClqVuGWX0UMRMoNZC0FWz+nb2vlljPF5sxx6YiFFpeGqU0F12WmnqAqkqt
9+im8TLrxirZuRI5Yvo2qqNymO/SkimmYBf8R2XklLXtnsETcaQoS9hsRQw0gC5Vlposd47pBPlH
PvGtwBIQwbvoZ97phCwMA0Q9kQS5Coh4IkJAg9EKDP+fS6xmQo3XqPQccjbbXSRoU7ynEJFgM7eE
pqwl6IcbeSyzlI55eicWsbS1V0IFpAhuYUfUZIsaGnAmhgRVGpHw+QrnIC5/oka9jW+cgg3mkp3o
nP2/4bDy++QbSP902JmHix9C6/Ll8iCv/sTTZVIZeG/AKmtGocQMZmMhpda5LEFS1I63SaJT36lD
4VoUMCzsQjCHDRS3+Tfjfh7m+jpvrU19pcLsN3fl0hLrolWXqUqROf2GtKhkO5rXW2iQxpbL9YTn
fpRETh0ht7751Lc5fyvRZVxUpkz2lvCyafWbkGRCY0D02S+mISjDqQaKHCIhe7R+sIRq56epfzT1
ceQRHYyTRF7kt5hGsYE0jHvoD9Jr9/cTrT+G4gCqPbxZX3XGaHFhlUdIn5lidHKCd0GPXNZgjy9G
wJwNb0I9hXtd4EcrwiRGHJUMKEIKuDW9lym8GhGieBNztYD8djivYkVKzKl1uZXiXDMXXSreRvrv
0KpdBAbzao0oiK4c6dZ70A1jZWcDaPDlX3QgxLLXbbprzdOWlKtnN4bF4ja8TFDpcnhlpJDcCNnU
ed1zy09gnOegYcT+KwBTbIHSxXRe6WmGMD2qSyHaUxEs3KuVBGRMkd0IPUknlwwxu9KhTI9C8J7E
GdNlp0JwhvEA94zULxh1eB82lGpmHst34sLw4xw37m28c/PR2lK8Z5IiQaf9VL4ffIeoR8Aek2Gy
bh8Ay/ljbDV8/jtS2fp1a7oA2pI3B5n9ZGPPPz7//dAUn0hYHsKwj8oP9ig7bX7OK+5qhKQtjqE/
bo6hHAwNE/vwQBpO9OPa9lAufIkVSoM4CbhZw0SEj5UalH71S1hnPyRplIWDkZyYx+TFhWajXl1p
uKqJtEX4E8Q9FR0FZcUzIG9lexMVOPY0ghE389m6gfXz3DnG+0RmXiy4FZSdWNWcannIdYxbykwI
CRz3lcpxnW/FzXzyHJfscx+6vfuFpMWPtO97dYw7uAC11mF1d1LMv5VsR16byRe9eoI012sCIj9t
43SgznlF+gY0AwMCW4/OCaA2VISlvMdX34K8wGjVo8gW2bsDpAS/d+Ze3LpGiQOvIadUFJ1x4VPi
aVI7z9oEqHreSdfgsxG2AGkq55oT/xtiLYNpkl0pSI8ZQRso6tSzAGH4/E3WQpRvJvywO0ZvkAeV
29qpTXChj5xUI6HSPh09+kVMdTgqd1HY7PzfxgissG2+YeBrVNFlGaxGiMuIfFPCpWxTJspKRA1D
uMOlFeFSBtBUBOFIUYZGzUpYaAz6ieTBScnF/KpDzALANWxaKZoEdJQHphB1oWBSV6Z6FpHP4W/A
utgEGHevM0jQufeQlnkSXedccUYVHeT/bSpK66P3IPncGY4GTnsVMTGSXrY/pWUD7zyB87D8qG40
nKwPgcVPQfRjf1GmSFghq/vGaYkFggYNA4ZFPwGtPDkMuabKYx1cpUdHGQ/8+jcksCnYxtnJBYlb
unl+SKZHCRyorioxS4DWC4wb2lc8sWvF/G6g691MBMgR3nHy7cD40diKMMV92Og04X8Yl+GZhr9T
xHZG0QwOW/Y1wTg8jmz/WGQEGHUFOy53p8uIKbqFY27jdp+mCYgdKywCU7ghqSOROnzwpXKvJbE5
wNrgIImJB7eJa+nfe/ByHCl2i5HfQyYV1ykWBr0JgPOrLhfJi8mW3PRWJlXTv6tQOyvEnLTSsdja
qV76HDxNYIBc26k62yA66jkMxa4prh6eruz8EYKjs3fgj91BVKdGdJ12KUgG88cLpztMEgt45Rwt
I9r4flfhzVXW2iqDQBgDYUU9p/ZexXyy6qMuuQcPHPd6H0fx0dIj/6fwQZ0Ml9dKKYt5y38z5VvU
8QxPuzJiBYTaUJ7FTIkgaMF811+8hyIW3clIZNNfQm91whBMunciZ0DlL9d6hTI8VMI4vH1pI6rC
x9sE6hTneJYjVOELf2F7AYeKMXyqqWkNnxrhKnQ+/GiAWs+dvw8ISVbpr5N1Z4il+E+sk8mKCphb
UXj/vBy5TXl2hHQumlt4o/yZFg427oY2WWSwvvRTcxYWMY2B13PdO8tUip6aFq2/wAeyj7Sl7NfC
ZQt9CVjZnH23E8/9ai6JpRwTNWdzAzxY/06/VPni2aX2XV7YA3P3O63CwFzHerENKTv2Ujd0oYHG
Obc14UFDYRrNutsCFDhw4yPDOMCDxMR/C0vJirQBC9EZBybkRoOKP/T5m4iUxWK936lTSr1R2Len
Q0tEHn+W1KPdNEVRjnvepK2jWW17S1QunSxOvOAD0EqZWZMHNMOnjJgwiqjW1/qrCjUww/8OVDCY
wcABZMXoYAkxNMwxvWoOV+rbbZzDU9Ej9bfR4094j0H+ZHIWTWBkh+ioKoQEQy8w6Z+hO53GxZBq
AOdvLhdscMsWnzNTear6FipzGGrm5CSWbykcmR4WMxprWcolOWoJeyBZFnNDSnIPblmqXXgSF0Op
tk9NX6Fx37KQQNEa7gdjXb2NzjRYDor3bndXon1SYApTZNLJTvfUtjzVjxdb4kOKUOumzbebsGzw
5Vjw1FmJ+NSHfPBqz+uRHzr5aLRqcYedUDgkZ42X8IGjAsRlGjmu8cwfITbiPzWBnFv8Emo9pyZl
i6XnPE/5RK4Ct9PB/IYoBGkGTB97S3Eyr4ei81Q2t1ZM7phQQqrUxantixjygWIsOVhrPrfzrt5K
uG91p+07Ezs9T+R0fVH64r4M5ldFZrmO6ExfzlDsWfy5FUiMsrlYyTjCJSCa4FKiCYWKG70xwC99
E1TN96ZXDKJfoyntp6AR2tPuorTEu0cnxjOPDPzY3oJoFEJql2p9lwNgeqzAqa8POmD4EvfEzxPZ
ZT6XetT74S2/K79infF0ELsuENEml6wqNoSlHLY+08f3jcMYuv1fs1mUxusKxtXGRQnR55eL2sYo
vFaeyanX+7Ob0GMlZK7ooI61NiuXneHKn0BDwIGOz4irrEfA98bqpliLm2yLB/xioSQ6m8HxwpOd
M88PXzzmQfhfGtkySzf8UgZaYuGI64g2YFvtPYjDgJnsOr4BzUuu8O7Vtf2iFYiClb7m1HICwjeP
ji7lEF5Zj7DOrhESyfsZJZ+ZVusrUSfzvqw4gbc6b3SqbXdU23xCdyjWcXpeOVuuVKCHV7T+URfo
ZKZA/21M3LmaVa4DiYB7VSdlsoSTX66d4Dbg2OeKywqi2McvSNMjg1bxgBpjqTWqMUz1uY6/Gwn+
cAUohdwReTfQWcUua4uvkvKtSdXfDAGpj/GthSRsuUadL39kTthqy7/AiDvZbz/cKUIMkuVKf6y9
jo3kBes31D/Xd0JOj1VHxq4FLMxYWxO/XABvXH3hLTJfTagRDvkrsWfW0syu0hMPURqlWEXsn70J
2N/3nftHgw4cHE7Rk0994KlaW2OFf9gMinqBiVW++6VsXc51JN61K5toLmsZPPK2bO/g+O4IFYsN
9CNaKG0nyeUPDPEZXr8H05QrGPg7/9x+3nQqUXz7HwUtrfK3Zv888oxIvV+3C4Fj2nYqziavXW+4
QCQMHNbyBAHWqGbx0/rHns9DQHOl/Jd3M6dE8slyPJbp5yhxsJ4GuN6kh/tHzw3i/F7kXuObotsc
z++CxyC34WWCaGkeCoJN4Im968TiSvT/0bDSGcUsQ8/MEE+cJPzJydGPvVH7M0G9hetGLYJydoeD
zzp2CG0cAXyTvVeB4dmqvWQwJZnDAb3SwvAiiQoxp/lfRalTHSGkNGSMtvFWzpb0q+DcotNurW5F
VnN/G2+ssW2IaOXUTeOayAsaV39YBRLTU9M+uLDU+irTQ+RlfeoO6L8eUC4t8QDFIuy7d+dHoJ2s
hj536fcH8fn7pv7foFanvTDD0u6qrnge4rauAaOJ23vOgqYt2YPZZHeYY/QmBtqbxk5chpYgflXK
EOVbx/Z/HT8bxrNTB+xN+GIkbGbTgHDw2OmXykRQVkCRONji84YNocEby4+f2ggUhyDOKUbXRwdR
cRg8UyhAUZjxjADMnXvWhjzHcb9DL3tHq/bxrI+di+hTNRu8l6oPUYIXAQNLmkkLj4WaQDHpVU4j
Z7Db/KlrVXf/2tpy0iRa9LYILV4y+8tV8ZsuA0FOsnOZGh+IAlNHb2Q+2XYOEAFMsrcCtFXdGvuf
CKMKDwbgehM1cbi6u3wD8Dn/xvQWBqQa0rVbGJge0NAW3xhsQLz782+QKIsnyG6vVwiSlmcAndxb
XemNh/UHkzwveKcWl3She++aOdDntCPly/Qtmm3qNuU7D+G0Blg5yccFKjOj4VV8T2B4xMuikTpT
+3HJ0el5XIQG/BZXqY+KjBPZ8GZZZ4e+b0xuKTgs0ls/Om2862B0SggGl3UA4K8Vxw6VoaK86Hg0
5pA7fGwqRbWkCI8dcRvRnRr8fDfVNB8K+faYrwRzCyzvarlwet+/tO7fUJNSZ6n8KvObbMSXV8MX
E2C/Yft2lluxaHP3lBCsTNV9W4SWJOUpmu/EasRmHkfrHghYw5zKVqdHJR24g4MgJ/Map2KYt1Rs
KubmeXLMCCaiBYX5GbJw9LQhuDqqCO3AlQsiE08kLfDjO0NqPbFmS7fpU/Dss58ha92tfmHI9/S4
Y/vM5GimG4xD2PlfaPIdOENTiQiJpQ+HLmmpa1udMJqiqGzh/9JMqCNcf1LJfL2k36X/rAhvVXlz
WqEFzwt3z6cwyO14RiL9OwjSeiTL6mJiJHprii+Hmrb7hZrbdFwfDoNsNbL8aD05XnqWGs/GZ9Zi
KWowR3xc29SsxxYloIJipwYAWqCXT+KmXzZu8ovqqdGXF3HKuJ9/fIYJrLVhXQq78CLDvbeIT+bm
Icf/HFK1mlVSL4JFdl8LxHdYoBIPs7YDyAyRmyKW2pWPr9JOklhR6afjcSkaCW5dmanUDOL4R5xY
2muLYr2F4B6DebB1NEXArz9nJmI7ILYQwFp4ww23OaVk5b2o8RiSAN/m32QpPHXS3oZ3TaxObc6c
PaE+DgNn3gis4QmvWMZ00EikScE8kzRLW31lzxzQAwCuyTgFO0Milco6ZJpZhiEd1mZvqHVV23i+
4nonGv448VYO7O7eufQP3i0CJo///d4AZopQXLDWV7mwgiqxptggoJsuV6yAmQrM53pXW7X/fMY1
ge4zzIPKPKb93QS2z43i/9ocX37N0Ld766Md8V1fT3wn0w0kr7Q3QCvT6+FKx1tgEGReT7ctvkvO
BU7EGXu37Em9xnMJaJBkBnkKB2yjCpWoAZ2HLBnSIsPKW5Es1PCUXDKgLWyX4bpbxZ98g7xdTL6T
azfBuviBh88VaEiL95jLXapTZiYCdIHy+xy5yxfH10hDZzrpQXX83tJu02RwuRN4nWDMElSg/DJu
N5GKv4O8dAlul9oeG1leB/h+lNR+kMUCIY1bE1ie9vWUyTp01pxAVsY/dp/fcADjQOXn2e9222RM
oo6lE6RWxp6+SxWOdTsjErO1PhMBE/K0luSeBev2c4xdfbDMC6tkgLQC+tE37bvyIO538b534DWq
eyOVH9Fhxv4PZ3l4NG57DM3Y0/Xe9olOuRz+211oJoTZlvF31OLlmBlh0f+OGce+1FArFfMEXJ/b
S+XlJ+F5+g+NR5Mt8FYCciUFJybjCnrOtTuSwnCeh3OfYi5bT2sDmaBUOmndqRrU+uJ9y1iMbf63
K8IBGSHFqFmqqRzzQSukk1CwJC7g0u7wTFVYc2vp/Fsna5pMxqtFt4Z+wqf/fO//xd4jt5WuJENV
WMqyP2c1MYNmbRKxvdi1e38wk43bV3yafa4UM8r00GWX9cfFssgdREV7gKp+nuTekXJTQ5s0eglS
IRzL6NPcsROwoElBIPQq3vifxQN3eAchD4eoPjzsg7wmf0xzm5vciAFPNz7TSO6UWLHRP6Jya3Ny
fe6cn16LPLP/xG1n5mGW3EslHP4ZHwig49XMFHZYt+0XxSK3/4MUdfZqrtPfF0s/QxRLdFq7zgRv
Itn8CWqMggLXqwG84o9Ivi0gxCMNeN6RAN4mgc75XQLBFd/Ief5E//7POF4zjZ0ugmDtEjI0W2Qb
xl8mKzRXJAqOZAv5zQslP8pW0frxf7CX5IKCCPjetnD/bT/6K+4iWt4nGFg1Ui3M/DXX5wLkA17N
fHEc6KI/aJ7Hj6mtqO9ZBvgXEGRUHsBVtBNwbcYE5fEokquy3S97wSuhOrDw05+GgBaOho4JgOP3
2tdqZqxgw2iC+fwCJXnTEeKjCNOXx/uQBjODH/5/XJWWNlZjCvJwP+Hs5bd8nOZR6cF9gBsu4w94
dms7V/7fgCgeBPkg5uSMRXBYzuqce7Qvvnby6HNboVfpCjFdZjxGK6ypurFSyxwUGhipD8fqLGk1
xbQ79Kh6hxjhAcDu2g5fmcArbMX16a9CbYwcLrfWFNvLz4hdks31ZuVW4GL/JrGyo0uTVhd9umlX
PSBDBl5+lEanzkqyN9otxvSi3mvBaSjOCsyLp1JpXIQQJFoIiI4sGp4xaM/YaMeKkA1rgotVubWo
RCB2LTx3+NrBFQCs54Eh0IXweizxNx1ptzzqxOHf2Nf6uZQS+h3sEMb5p6iEihQl0aJ4XJ5GNvOC
FkIPNmPJ9sVl8p35zShX3+XK9lNqHluZhxsFCAh/Uzwe8L2mFLmEJqe6Mo//A3LfiIMQyikUHRIi
JSUz2EIgIlNSt5lVfeEF4TbTh1NkzcPKVuIFMgZFfys6mv9NlDfhjTF+aC43NZgFdl2kEk+BSkyO
9iHns3WNAYN2N/TNS7hLZbrQg4GYu6/Uw0M5VXc/PsJsOIWALCWGTIdARL1qkiJY86vFrDROytfZ
X/AH4R3jQqcEErzGT/swMbZ9dbu3jMCpgoOQsmKl3G2kt+B9sQWVn6LO6RcEkmETlWPh4MzYCt8n
6deIT7UzvGnb2bucbs0Dc3S4lc/Lncj0c/hwqVs4GJu+2yYOkgXZrE6+S7RW/CD8HMLaUN4+6Xmp
HFAi2c7wshFS7wqAdAOSpM96aOexwcHy2OpyTD//2RFW+ekXXNP4ACvOPG9ul679BEEXY0jw03+J
jCyvYLHC/e9rc5TSLWe63cseSmo7I0Yvo4ugCTwv9dT1jf4fe73Lshat3LdRLExEtp838uDudB95
XzK7Hr/BOs0WTiw2O51elA0ipZMUZd8COvE4BPLh+n8QGypQPf+BkZvgU4H9pDTxDCAi68+H0Isd
H/tBcZ3f+EXbkABajK1y1H79WdAJHl6auA+5LxJ8PMqGVFfyePLn0tezaRJxomA/rCZXwTEOoIg+
/Pm0G1L9VzBS4aqVPAVgkO3bWPyZ5a8wKyqn9c3P3VjIQk2bagyG4VdHmivDEDh2KDTqRc0BXuE9
D5pI3pSzwKXWcH4BZ0TnzxflqoJFY8hButymXP3pwbjolb7GXzqK2sC4aQaEAH7cAKZRZsIbyoYp
w6T0KivSLzfFU/26wnsUTalv9mo+KeF5Y1tc9CxO5o2uCKT2Y286MBAinAxnCg6lJhkAbs+iGBc/
E/ryoteSlaniwazaZ/FefXgVYBv1xfz/yp6xMFelYzHqyEaFFRNHO+itB5GHUrnk7//PfYzfqlvs
eVf3g3z7YFT+c/6sjz4mfwnlPaWxG3kBtSq2XGYC88n/ckABoeWGmXTaNwA+kHDm8RL/8TrKlDFi
TAewgcY1R9US8WauhSkCU6QYuJAJzgioVN6QupTyD0BOnpeF5AUZcgWRKFOHdkQUhwlmWCYFatHo
MF/CjXdJkCXvHR3axEJCWrfOC08EkseF3KlRq0IcOVDn9E3zXXRePb3x3PGHH9BkB2fqPsut6B9P
tBSi6VwkCHtCqaKNl08rLizc4FzA3L69Jy3zhf65N7uDLyPU6HkM/2M9U40geWwI3C2nZwWbTI/l
aGPWNOJat1E3ic+LeSvvPZ54PxpyvVh+C/WjdgKvWx+UIx3cimmQXf7D162Qb1+OekQrKOb0cg/O
K1C6FqzAIy4S9vEh5jtIBN3yGMskLnK+g9JTTNBpq9rQ2veAxiLLPIXAT0eVw9O2K2JJA3Fg/7Ed
bEMvXXVcnaSyWk7C4afHXmWl0AwQUZlH8NgYCDTu3oZcAKwYXSTfI/7/IUd5je/wkS67juEQd5Zl
4hE7NBUFdXuhGDHqJucg21Rz9Arj4JjXcBLa37bMMf+9T2H9eN1bjgu3PX4xm+5WSQ/LWWnP7KJu
+Amc6CakiB6RfGur+ebk8owIs9rvSE/Bo8cqEVJ7rBnQg7WX0EA2GH6Lcorc5KhO4ORsA5j0pn3d
1NpFcbOKPU5vRUw+y337tk6e9wOnX5phIXBEvyDGsXuKhqgkac6dATsvo4ZQ1oQdj9JNLYLkMGW+
z9vGSGQFlr0Mvj1aLQJQbJ15gcPxh4yYi3jbARdhoxK1jRljol2vNwe6uZn4gZaP278Y+s9SITrw
LVtCjkZO+MLY6AzeQ8BCJ9hRmrNYOHBPkVnhTcHY8w+nycrkuG1pBjDH0Yt/KtXzPOLXp+CsXVLk
TyxbVmkZPEV9Gugxs4KOJKjQJnfUrO7JtOmtYjR/kpPepOH6KI45n5k4zgluG5FWeZ1YuUxDfLON
ZDn54pYQosQgunS9+czXm7BS9GNvEEKfRWmfeXqsy3fTDJnFgHeP24e7I5DSsf4V+kVMDhD6m6ye
dcl9EzerkbmE+xI2JUJXbyX7KMMHhySR01ZtdvSqEqAml3bV1tyJpwq73lVra2svY+0YLDVexvcq
eRpb3E4pC+s+r9pCpFAO/u0Ad9oHly33kiVysSJFUZm/oa/NlwQ3yAoFQ3M6RBL1xIBaKOsdNK5P
IoNvuZS9yo2ZQj4uHsS0JjRZgsEn2GZ5DjhftL5le+jAFZE4ZU8qqtEiHOB/d+OrO/xLWM4IZ6eK
uUQKuhv115YF61HMeisT0nmyVKn2xQB8XunP26I9NyYjZjE8Nn2QocZQ79C6bwbDsyIKGCxy5DG1
n0hWitgaf7LETZ2sEXjX1aA3Z1YDEudnh5ygqE6SkdoeuwDynbAMBrqLb3LJdQowLwOprC3kv/ZR
kdGqhSnA6cUg0gc2G4pq3O/4/0WaWTZt6zOa+w01SsJEibtzOEOY3HTvNVCFsJ47DJ//D856o0aU
RdKTVrhZwJTCL7AavqhCFz1xmBRVQlc/y8cvSXVM9cyg9Abt/4zEuJ3W6eESVVwv0sL/4UTLJgjP
pnBfrPQAuJx2LyboS3Mggsuuhcw/47jP7Irq3AxerOMafBwzZCBuOD/QWBVvtJtExVspnd/UV3zp
IRAg9V/EtVAnpHsptFEFkxrDurbFOn6K5+FIU6CIbgNUZXWbG+EiWKgr7EOSlz/DF6CV7RZsNhE1
rjt0xlVAYHW5PDXA4S8lwEjl7sb6AoLHl2UzX1Yv2j4vYoQeigoOmwP96YLdr6uk+pi0x0yHjWOK
YAPNgxvL+I0S+L9svYzyUL6G1Scf8X79T0RDp2ubi8aN/8UpY5ducYGvIyFZUJSb+YMjYRNGjjMX
gZrJYmp2swwJOl5vPR2Ujjvg3L9vwEAl3yxsxLZdGl8ak5lZuSHswsNNwHm5PXjChcgEe+B6dto6
1ITuQ0v+j5svvIFs/0tqKjRUId5rv8OU3ph7jas15kosNljOrqefBoqdF/q0o+gqls1C1mwVJolo
C3KTzMAy+WJ8CvbR1nHZzT7peupZ/utMyHmJXvlnTFzCQ3p99OWmVq0we9coQFpafjzgs+zoVopS
gZ9hskKmYqMwotY3emH2Bnq/yvtPdwnXOIMREgzN6TjElZZ0l5vXTwcMrkM+UF0fmTEqTSqwtl6F
L7i1UP0K5xq1s1usxshYq7FFvFg2LcKVEWJtIRIqflvaiBy7kyB/IZXu4RRBCDZ/RwzeoX5+m/XA
XNxtjhR84NPSVXOoOJsgOJE0U4OxWRO3PokJez8BnQIGZhva8IdcSODWECX6zjQYN222GPGfsF9T
eZ1q4wzIFAXDkjcw/8PpM2ENWMpYloI44wU6cWefdDfaivsgeNvf6+exwp29/z9+l6/hO+i8rpD+
/1CIlg4D4V9F1gFCMZkMIrF1qXqCuA/FadqxaUtj8d1dvBlCyncPP70nQMa+mO7ZUsjx4RwA5epf
p5Ea+pj/vu3R9SmhRsDQHp5I/wWXRobHaql/T/V767AvNq4qrsf9YyzIVIzsanPAg1OaVK97uaUe
rlcR4uLDSRJBXDI0gJSRHpgtM2l6VRWCkC65nQHVShpd1m/RrwN6xcopxHwnuYL1RxW2r7qusrGV
a2AUjd6nnj+9RlGBmmz7WGGFDiBhEM5QU3zdDcWXjCh/IGZ/zBXfUSR0aMh7rSv2obCj7ZDBMPGZ
ZBF+jMf8hD4QixggoCl+pZlm3DPDhP/WQYnF3N9ZdPPboilE6YkJ2LDXzva5L+JlscmWEg5oCGpZ
zE+lJpTEdNLrHzz965iqo9s7bhoznP+YcSorM8vNxkWw5nYtuU9PilDUo4EhKUrmr8ic699NDLVE
u/3i7ulrlaRq6XSSkkQG1BCUogVYRChWTtY579OUbk10xQjFOyL/UJV3GxWgwUaKcG6ufS1Q9u3M
QLvc6ORAB7p8Yrtwd8DDKRYkBrULJED7SYDd7NmkPBIY2OEwH2WFZJYDzIienxCOice6VW6KA/xM
GzPhClPqv/DhyCTn6s1v3vfsgukudiqcKWQbzOPS4rUapGjM/DLH4n7QYtf08ptsc29pt+exHufO
InQ5wyTQqE4E3jXoX4SU6AS2gi3O+l3xnRFAtmkRc5hb28741XcMjiqyEsxAk3BDY7CIuL2FeREY
LDLX1662WJVCT3cPgMjlQtsZZ0Of1yZI5DKQ939ruSEkULIbT2IjUtu4aKPZKJ0Vv9ArFxfj3PFK
WniuKn42+Dh/+cYqsFaPaGr0pPTKbnfE3jnkcCi0ltCyAeIcNueKeCStqSJ8Jw3OQNFcvv05x39G
etR/aGMjhVVJsza81VpGKPN8SkdQ+bE5ajey9msdGILKQCRLtL2yNo4a4rl/RX3dfaAn9HPxyw/p
jnWQvih4iOHGMYcVf60XYaINhz79BiOGGJ2CitvvO9DDJGu4yCauIHrUv2ZJ7E6ye4bGl3Y6a1MG
G5fBxKRLVRuNhW7VgngMR+gWjGQPkrTOCYxkwntflEKqI2V2MYNYy+8ztg1qpkJzSxSFmbZU371q
1AUr46tZSp7mS34zqCUWx0MDTYAN+PKGGHE1PWf2NeyhNAt0Cx4gT6htvEeOPQZz8osLYLlbutRP
cevrtttz5uJU1DsiOCM7kEQKJw4KV89btrvjMBlTmaGBCj5bK9MCVKoIieEfKRA+jnUrZHMtMHuf
AYgDVacEVlKnqVM1VM+fXUs6lO5mT4LOIYEI7bHYum/CCldv2VJ/pb0TX9qq7ITncLQVDBQr5uVV
L8BCSAnrHmtKwCpOf6XGQxm1NptOHPrXHCqUSojO43CVveO7TPXoVfWurAo/AODkg/gzFUZh6MaA
T+Ngdwy+6SpKZzbvYTNZqkdpkYxvFDvKAPKRcVJC3tfqSBANYQyMxQqljxRBYn534PwIcGF7ojWH
09Ci6kytGiSITiHEPFXWWxgxmpb+rHSsMykBB01lriobIR/TS0N9M+9tYsBPIDiWn20SgT2QtgDY
pAPEbxl01zsZmA0dzSzFN4o7oGu77YXXF7xkg5sSlwzxIbUmrxYvlcO2LmS41uDy9r8yLzIpQ2O7
0wKH7qhoftaBg1yv2Z/UEptA30DN95IgzMOvBGs8JvJ5LiyuRqnkAZPpJFVaaFoXOdODb05HH5Ee
zVbJE4TeitrULfcFdNknU81JtiX6DmXkWZVrzufZUgFEPFxEVHV8n5dIWP27KH+yeJkOHQZ63h3L
TRpJrxdRXlq91GjQtQnnDMtkprFdEW81XLYSt5jjeuFLDa2OV5ohQLTA6hNaMM5RReq0fASB9YWY
orf/Gm0il09fniUev1DuHn8DGaDB4YenJpTR1rWlV2Z1z1MsUM1nbTJiqDpjAxoYpsZgigeIdhY8
SFZFrTCxtslU8TD7ue7DGmKKYez43gbiwi+gyhpxmDD5tJCs1uiCjcEyluxA/z2bsm0IsvmYO+xm
hGGB6R6yUM1fLf+DUpBBFT/kTqGTtmFiDBb4uak/psSOVEhuQjfI8+J2usGl3zOJin17lRVgkU+d
0D9OVAlNE2GlgozLQX4B4ABmEoHcHGjW0Ba+gfl98ZxbVSRPCB6UE+4/JlMfu5iViEGEYpinc9Cu
ck0Oi+8QMRc7dhQpUvzG7IkAzK9fG62kwfYktkiZbKRxA6LaAAJ6W6mibwnrZVl+Pd+hYYMNVkHd
iXkEGsUT15+5P6r/IPBzEBCZuofdXsg7eknajy1B54sEXu2hdDUv9oFquVBE/e5D71VYLs5Qta01
4Z4Mg/nh2jMfYVu39srElPPdkj/CHYDjLoTgC6fwaGUhqlHI7ePmOr2o85ZBG+hoDkr8XSfI6NSO
LWY+X56Ed0ni8BUXJ5CkBTVxmQMlCW697xcX5ew/KdIShcU/ezX28DpOtLpdhvRhPJ0ayveaMAxO
5XzRgmWhIPFRsxaLsUkrOF/0LrmxSKkdcnu6xHwWQ0dcrElQsrHbpCdkSxmUgpY2ZDaAPKXYUbv3
PIFNwZQzhAjMgDSZOgar8Hd+PzRy3xogMzNXHKNnxQSCEvF7P2J99eueAB7MgItQ9M5aNU7bFVt4
GjAjIKGlXZY7MmjrAwfEmLx7claLacukZN6MGu7x2gcBGa560nmRSo0+ACATAtWnTo4r3+1GzmQl
tzZUnnLvlSiMFlu/OAkpXttt+nSBVqDURxKKMio3W4M3Qz0cEPPCPjEVqvwWFdk7hxYX1v+hCvam
tY0up3cC/cOuqFGAdJ1Y44IMRghN1PXiOGzGhtxCDTkN/7wVZN+hZ4QxDYk4UrjX7WJVQhVpUR08
WUNc4DuVEFwYLGFJWZkx8fZNNx/r3ex2kb1y7iZMEyB1fiPjURTrtJntLGW/eG2pvpYpE+mxGpNe
ikfELHcwUq7rtpQkNapapjqdXBT58B8RDK4ldeZm02pWtP2s2wM6ORM5iwlqofziCB0klFzWeY5S
4c/hfbewrW+EbBDR8eedWUNcvToLBVULGHiIF8e41A8IsUFMpCdEn54OI2cqSjiiJOFRJjuMiZxb
j1FboJN+Qou+jpEBATgGZgCnfxLAl7uuHjCutSss/xC1t++r6bOeHjr+Wm7nTbq8P9C/nfMWMTi7
f24+wbiZpPL5VRCoN+KFTU4x0mwmIaJV7dr4O7Fq/Lb1+QO7tJ/cc5wxFT1iI2x2WxvJnPf/liry
6QcunWMvcIlJp8gNd6oTuCRtPeguj5ilpASCZ0Ux7vyrm+UX9l9hq7d2HFMtzngqdbkyKEy+NZzI
fnXwqzKRI54RgBJrGzXpBgWlXUG3Ubdu8KQM/oypMetyD0e34JOe8BcFGJwDxUEwiQXWc5NMPymK
3bQ/c38zCecd2oizr6PjnPoqBbg9Ed9zVgZoWrLbz+uP2pLc4SbnkNxM4AFbEgBzZ+PXMlhF2zjS
CO1kqi/YnYgkq9yn+zlFSLgvCrYdOUnzfaqJMFfRSEKSNezALFqEqJaTJVxaR0/ioghg/MWVY2QZ
1311u0VDNt4/CUQmUfQ75+I/fFUEIJqBYpCLtppI5TN3UqMxYiKtXVj3Vt3ORkT7TyHXgTxUURQ/
GX3x6aSdIbVZv6IMUNCctMzruABqm7bpf0daa5fI1c0aGqr+p44KBE8znqWBX3enaKKZLrRTk4Nu
6SnQbqsP1ZKl8p7wDW7qSoNmAAy+2oJ+w7DBrM0sUR4V/Ku8Su+Qm3G3BGYyGGEno1Poapl+D2TC
oZJgB9pJ9wReC4ItxO4SEWZWJ84NEB7wKOG8Y+DPRbqxVDx6ao6TtC4qQKQCJfxgRfgwYLjnWDJS
cCEu2p3V4xGODz64N92zUI+2XALB9OmnetV0SPAcs3/w5hw7+7vpw8jwEPZbhXqP/ByJ47a2aPTT
x7j95miy4OkcG8+PSbAU+qmmnhgg6wekBUOf6H/dcnwd57jS3+6Ig+UZypy8BdoDJHFkX4yxm0Ku
Nmy4WeYbXVeFLjnwOSoX/yivu1k1/qEwdRIbf0IUFbtoJT+b8cZzF5SUc6sDuo9thTvC3CnGc7mY
etWBf4mJXLTl99MdV2w1AC3lrv8EJIXh5y4IggB9RwJug2SUPS3FgfZMXvp8OnzzkjJSESGLrFrm
0ZGhB9rgoa9sXJp736aB4tuwRSa/5XWuIb/WHTSXoGVQo0reF3ivagFMiMwK7jBr5GALv3gxF37z
oPuuv/Tl3ZG0NfcT78ujbxBjrdUwe8LU4DeZvLSl/Y+UHKvTcfSTveI6GfUB4V1a2cl6ZBNNv4UA
JrsXTQt964l8mOADgAC8sps/z4OWTpXPhSr2mbT68UY6zPbiMsEQqhozACzpE4GxYdckFe5tNOya
da/kSY2UMi9xDX3L0VX4EHJcEnfjW5OVup8WKcUdA83Wyp3RUhi72aDf5Hr9asdVNF+Wdh1fMU+R
Q4SV1P0eMtARPkQHVugA4YQGGSPQ4hKTyx/oBFSv6+iooT5EkDd0n+f3TwVM30ZcPs8V0PA20f0U
Z+eyQDFVGO6t03sP11yMY3IeXS/h2XWlH7gzlv8wFCxyt6L9ZTxtRBnZ6gvFZe0KUXUHqmP5MkTK
24k8bYXwRgoLqmrYNwMSbO3Ep2l0DVeyuSAGxp8EuQVQd3zeif+ECyY6Mk75G20s6xFzggTuMdry
IW19FKOmLPg0/E1AlHpCw9b5D4/rkjPUfTPKyxo2/9RWaM8LU/cwdqO+CM+iRERtk7fV3IZP09W2
XNSs/yoPhTZ4j9PDekJz9s6CA2K8KiBe7IpjNPb99PO8lIyB863o7yUdO9+rkezA1TVEKsZ11s29
7U2Vf6c9uZYa8MT02Co9RZ7W3YdyEMLY2X/7+V1JK8MjjfmONSttjmR9YQl7tWT1PmraG7vzN+/d
iLv4g4KIWKhEZzCPNaSCqztsKo+Juf7JX4Qgc0TeXHsNcqoh4GGLh4p1hMukv57cN+QayfTpoP1L
Q9mkhmOBT7wqK3eRsfasnaWpv3Wuhsd2aXKznrAw1dyA0PEXDHOwaim0nGrZm58WQ1Zo/bpEc1AO
MMewq5sPLParGJy4BSL6NItTPYzmifoDawLcejXaSHGZKhWbjEGnAZqQe7mN0M5FVBKJ3uccnmgC
7YjWMrdwCRKY86xIQVDuAoPjJ+iRqQhsyNCot68pKNCwLn62DW1qV4rjpJB60vsYY3PMOB92coUN
NbkamS6BDTiFxUB1IL7xIlBiRMib8Cd57IFTfD/7RVXzglYJzCswndiZ683/voK2yP+FnYL+/+yh
W3BI7JLQ1Mu0GS+9NFJFA5/dkJZY8XuLBbpv+x5ac9Mu/UsDdYlvhSk5bg19Fb3gV19jsP8L6oFC
YiZ3wGfa3YhNIC1/HbYSa1SqGLYLHqX7F/UEb0NW5MyTaGojWwROi9EuZwTFW08wgVR/NWxXusKx
mwN0uXiSun8k1i8tMyi87k9g4yV8IyLO7BZJb+wulJPz3ygHv0VeFDafiWFyV6ocZDtLiKeHHySH
LrBn1oxY2WdtkFlynfsG+waNTZFU1NEpncQNeQTsfE00kdzPELxUyYf5S10XTCFYUlzLsdH38QwK
npyG3XvUUx4Aop0vIxcPVPdAIqZLwAlG+8rl8QzhxkQzT3ZGnwpmNgeeQ/DChXJ5MV4Nc1WAyaIQ
GkfitMqef6syCnNtGdXNW3gwBm6k9gYaaH6lSQweWkDgb11t7eCPyCQCnRTRahXAWH32QAsXbA63
ku5nQ2ZNfAguvKS2BtLRRi51LNoMl/+yHhHcryypFe0TT9s85y2W3c7mZnogr59X4oeePo2fk+td
xqVmStP6gU4nqLW4n13ToGpSlFJQDsZKBF6ZemW+0Q7o5nAc07HKgsyKLI9d4rpG/ZOORtyWOMtz
Wl6IMcAhM+ntEHVzhxRE7GcgRIlkseAu4gPSJ5V7YWvGDVAiQNLZi3Ieqan5MjsMKFUL0qJZqvwy
FOYXgT521rUcN66oSMu5f03gvhM17RsfGl6jdJxMtKutEcwb4yuMmZVSJVIEPN1NbXgtCYjpF92L
jgt2SL8sNvXv8zqozflKHjrpoHtalAMHu6nkapjMrFB/XGwY7zY27ARWdcCFikPsEiBkDVS2HtzC
GplOSR3D64fsReUAbLwjJkgd1Vq1jNPsBDijltZLzCVkOuKc4o1tkdJgbHcXS8vL/uaxZZEOF5KJ
q2z7DRLuOOXkMAfaj6fr5e0gOBXLd5SwSAfPP+5GYrnUxvPMNx9hjb2cSlx9r606o2/TEzPhdvk2
CSqFg3ozNYN/DATzKBCeK7TSQIoSKGfedtjZJL9XgDa/0b8krKwopU7qmwV2kU/6XQeTzZqRj+Gt
G64pMRWJhhyvIkJNSx8ZH+yVvtIyIIbGRIQUxUCPaa44NTCr6JsMtjAMKcve1ULcAz17P61fMoZI
qpiOAyEu7bB3hqcFWvWVwQydO6/pRrRbpkI90Vbp9Yy3EoX5k/h06SCYgisKKDb6Wbqv1iiZol9z
lDfSuy2PBoKhHK6UeEUBZFVhNWsJjLE8SSn7gWR5TixbJFnT5OFyd8EbzuW6Yhr0G0FqTKtWG57+
diMt6z1fFM7GpINTaA/uYsALXO4WhVzKzu8fKwmBGUPkKrabTyyohus2FPOX2mRJ55k9MViRitf6
56e4ImMoEqbUFscqF1nKHYawIolOcpMyEXa0TkA/43HKQsBaaJLl0cq0zCqPgyuuOPGMYsATI9HN
REZfVAhAlSi/qAy4i6LOVEeQa4YYmQ3KXaVTTkKMZy7P1shVMLa1qE9PwuCcogWh0h+qUDSOZTOd
oRru2NAdtCHo8CQS+z7NOvh3N0NLCHEEPqRkpEbo/r6jg3TTX6FJPObAbnBH4dN9qo7s+dF6S2jm
dk5YwN99acgTFpbm+jPa8e2+YXwbKYmLpLA4g8c2tU7Eyrmh6b0/toMvMSXtocr98GSdbIx+kZcQ
T1YJXuM83dFBQKI040Hi+TE9S9J63mlSZsPT1DmN4Kl2VX/EpDlsXdDPWiXW8Hoi7Wob6utvYqbd
Bb807Agp3l1nOzvdR6fzGEvgkvCMW86yybNnKbLMNu0k41czfWIABCPGIZiS59N72FUq/wLYAc94
A5ANMYJDYQleWiEQUU9jmvydM7Z92jQuPWAPGGKthROLlWA582vDlNTr93YeaiuUJ80zSspkUd70
iZrec6nMBPUKzZwTWlN7lCljilrWaS8Lx9lDtOzhzDINoUN5bJDV3GiwpU0FYtybEcFyr5EyIBoH
GJOSaURRpI/P7r7vwtDFRwsJRUvtQCH1xWpLjxIeP1MQrSxKexiURM8EZnHwtgHftynGLGId0nGR
JKGV/uPiiYvkwRvfDbTGBk95aEvYtGGr4taynYmDN9SKMbune6Xo3L6sxL+BJK9GxD9mYDJttqR+
657kIr9AcKMtA4HOAEDa+d2CGGzjBaQQ7kXmwyWh9ybkAJbznaAeLtUmTe8eq2VHwYm1PB6IVeZ8
Dr4C6loFjGjG+h3ENFndst41UOmLFx4GSVP+Im0SgOkYVQ/qNDJ3v+9k2bmCoXAjb1l0CO40IWTY
RW9w9JYBcn/mAp6gfwsvO2eQfkYEY8Ph1nFtFo/qsmHW/JmFjL6ALDVtKQKJI2bayWoSr3huF1I2
tuciun7LFbYj3NUde9CPTKZhtb7AfQVJIcNLBQthwKlclg4R0HI0xjGRvD6WzxncmqYpnbV/olsS
SkZ4iFDR88b7+pvLfaJvOgWCegCyY4P2FYOGt/DenlXYx+LzIUqwYQ4PN+OKIihhbzFUDRiMGmD2
J3VvNwymBE/4a+fxriVqynJovUIoO56xdTCJE2Kxir1NSa7gdO4lWwGRuigea+p5tk6osnqmKh2o
DmtaJhbaM0FSYiWyM5gR/rgLVNF9448S0Te5fCLP2Ml7uTLZ6ZCK/ZNvoYfiSvW4IYzuyJxTez/q
rN7hLDZdRuB4X7NO6TkIvmLw8E+Tz9wjY9lbv/+ZhQfXMlp2SPZQAdulI5JrVwwmugjOyxRjuXf7
So11iZwP51/T16xSdZrYvbPVlyDL1lCNS3iozNpPr5ouMjAHDrV6i+ngBEvq19v5NjKFldcu35M1
qTfPX9TbJ/Ad/zr4riWSA+bA5xxk1dW4InmocZDUPkgj2+8al51SNv76EaDsXkm+/iuJU8VXHZeC
tp0jI5/yIq022sPN/cX/xtuDfhA1GAW5zRhZImqA0vKO8wo6yNENgsHw9e8qnF4/h2w88cQOrXWN
JG25FDIfmDCybZKjxoiM9cOtpw05ksjUo8m6gk/u8HSME2ZPu7NAm/CSGwAv51HCoqO7iDgfW12I
LesU8Ar4K3QT35lHovnDekRaDn8497plbNY4NHSmcvmh++7qNwhNwbJlUrVW0k338T0vhM0fEe4G
OPgI+keA/iAiSWRQFzA14EhaWw1YVxkk6kze7K7U4ZGNBGr23BA59jrVbMktj5tkwO5popo4peo3
47yBY9suzkd7YPw8rN2rb194BnMxWqpxbyc7QGnpF3DhZ02nHU5iKI0xjQDfpNgNWlvk8aqsHxT9
MtbOiPBGRNvKZ+RfBA0hu1wE3uStzz5LziAWrUSsyOiakmNCxrr6tFraF95oI58I/QVujUVayvjd
qFM0D78wSbM/OwhcMih5DHHWaYWfmflsAq5b/2YyIrpQdPvzMFX077qss6K+NaKKHqkTd+wCKqp/
pFaT3Nc6fNHcZiInpKwugbt/ID3+KPCWzlwN7oLNe3QFa4SvdRP5GUDU7D0BLfdA78OeC0S4Z8A3
WRwXb1ZDznqrwMbQr3ij3mYLf/UB8LUN76cLh9N7RdV8VFSVfOl3diswwVvoRx5TRMlEQvR7ozxa
ZXsxoRUPMhTQmLAtc9pncwbWq/J/rF4/4Y/4B+iqwhOI0mfZvur1fGMsprpJc93t7v1ryGUN8p9s
UtPwtr+AjOwMOjOo5EXkZSeo3bMqaFCaoYqfYWTa2dWpQCRw6Hiz10uYfPGyWsZ4+vjyxW3QrfoS
TKTkSyieEzxcZsTRQn4kGkghrbr1uTMNOyryPCDZp9O6VCy7zuQ1vMf4Izim17ySjSfFO35pB1A8
W0Ufxu76SPmo9RTh95KTOwvN44mBeDx0vF+Wz8GdU4XlfGWeE1uVaKxIGwMohZL+XJQwiPW4CP+C
Ezw4aNFpezs9AjavWNbjAuIunajYcS8qX6gG7g/kDbUIA4z4I0ZyCm0sBHAZjDMKBkCCnW/8sbMx
i/tMnnpRL02R5DCUNuRxbYo5RnULaotbbs4tengfrei5JEXQzJ23YLlyPowNbZlbO7+kKB0NxQ0R
eD+lDd3oyH7XSpI/+D6m6VDwoNVSDAn/5+lHxcaozQiNtM/l/jtfkjnHaNoOEmdPYHhK1u30VYXO
yQdCyS27qKEkka4qivJOUZLGHfegtm42Mw7SrWuHeOXU2FMACrCT6ZWH6sc/GsdGBMcMDoykcs1i
7fIyXMt28DeA22J8vts7MZW9o4MjZBulfaGiB58I/BqfI0wcg5Jc0SEuZl9CuNuUTbncYzRP3utx
j4/q3Q7OT3K0dOoLPQsB4tJQC8uF2aNZz+K44tjGbFPfdSmURtpbyCTkuYPG6TbzGa/kwd194Wfw
6WwmRW/FNY9d4ayaAcbzDYNPJhuhscXekPQpRy50kvCAhP1qh+9AAp0z+MEuCIX8iiGcnYF+0Oy5
ltLS+noSZpCpjaq1lqTiqXuClvIbf2i2yf3de+Kc2foE9CsC4TOmbdwoP9VW0YucuXOnhJ9exbKs
+BIfmkVh6n+zl+YgZ+OX08sNT787prgJeG2OZjlJkNf+RkaOhetrZe73ZdgxnPNOuZOz7lPGCqZv
WGrFtg0oM5JaRvCy54hcm9bctEa8w3XYt3DBphhH6h/6NNxs++PWEAWrl+CFWj+1k0OX+/SgRBFq
+X3BTBFmRM1s+HNhJTqTdaVTm99vGLEId4MUtxtmwYvNvc3dhtnloffLqwl5K7MZfzProXKup9LI
5PwPuCb94p78jPn2zkSnaouBoKQ/kN8i2jp4PjGQqBZZwM+SV7mCdOQ3n/pkWtfCIP6EaE7qjyZZ
+r68ZPPUoFfdj+abzOQQRY2gNhPdXZvgw03unyd7+Tpdrng5XwO0sNfihE12X6dOWsZyOn4WiEPj
qPLFe7b1V9cBbN08ds4dHtJ3mlV2AFzc1dZAvlbjFf4VXXQoEfXpnRYj5+NZjxqO3tK4fDLZUf3z
3cy6fQIOCqo0cW39Kg8jpBiZUzGIJbKboK2+ZJbze5ib0QL6n7jG0YKu6RuZIDJnwr0XniaVOgx8
hp1d0MTewUnU1nkbbPXlMTxZYimSh4RRye4Yj/KLbq7PUb0sYiwWBlygfCc/ANeUXz5o9OZYcyN6
jos1SAXd1UzYcd+3g8LNJS44jruGoHMv4J5nS6voTusbFYg3KYARQKUFoE528CPB7vNtNI1u0noD
yUaSxDtbjbiy35+DeqH1T8K3pJHVG9jWb8nBR2sPKwg4aF2QG083YT6oiwVK7j/LT16JdJrcZ3n9
aSCjtCm9ynGJTFtbz8BvjRMzz0KWcSmbSZ9pEQnMeb0lqTKw7DVYZkwzrVWznV1/gL3z1mQvIhhQ
txvdW2MmTchJE65T6PJ+jR6+LrECbQGYy88yrYDOW5LKqXUxtREjyGJtyCp8WG/JMJwz2OHF3GDn
/Bbzm7ey6MqIap4YrrXSh7qLZ+XppATBl5HgDlSjxWop5C7mzENSqJKCu+HztFfV1veqG3Q9WICn
w+GGGPhyp877dvoSDc3D4M2K7LNvem43WWYv9rAAGLqHRuY1lk31O0fu1VGUIrW7U/q1dSM+JvNW
34bfVXPzjerm8agxhWZZ5QQ2GXhbkmbjfi9waB7ZwoTg1vnJ++bKWdA1+dEYv4G8GD/FdEEBQp1o
nMaaNEG89lZ9ukp0uG4ImSJPzqV1F24tZBij6tQdQ+asdCZU5BV/99bWT3gvglx1lC+g83ROd60Q
L4gtIx/El2lQHsHZ44yvJmOci3DrPlC5+pQ8t+ntQ+6/YOzwAk0arYYbkfK8/kyBJL1o+L85bBxQ
9Tf1Sf13x2lQfeVbbLxbLuQ6SltVNDTyRhlvGNNp5HHuCPxyBjwX26m8kA1+nXk2pH1x/uZmWAuM
vP/PYwrnD4kVgNDaTsS7dyJ+T0VS6rnGSvRKZw/5IVo9ceAu53J3ITo/kiY+pL9FdTTmNYF7MDPh
dl7VGSj+ebzvunXPY2SQC2KmA1Rf8yJ4QD4LLEuy/cOS/B0l819W2pTsgujBAG7a32ZitR2MwOrS
E3Vg0MeyTz+KidtJTP//XNwDnSavj60UJ6CLrEvvFg15k8kNYNJybvzAhWW17oIRqYppE04gmBlF
Dnvcc8wjgxSXuk4AUbc5ZXKBOtTmIGyJfjaIBp91ASrJldJjwIByLohnwovwn8eJrLxjdoPqcYRU
5CF9i7c6sg7LqMutgP4/hBVXuut+CjDH7ml3wrlw1N/5lipYxMAgrDLd06mgxbdX+LhZU1968n1C
vbayOwNxFiRH/9X4GBIaBRTPlcDFQgAJQ8SNN6QVLhHNIyU5tiqsW65TPJLy8avG87KhbZWHKzn2
e+d4mKPV4tZH74DmN/aVMAOgSPXc5TU87ESGlTIgYTm/dJ9pADvEgkWs9tJz5lKS3ivgY+65sb50
kyzXIVnqRjBrGnwYFgcYV8NQalAAVAoXDV2lQYwOJDOs2+gQQS6ium0z2U0a3GTD94NAZpxjEp5e
0oQZnN6WfgQ4avlus61hKA2L/zspEE09vhSfeTccmClAXm+giLDHHvIvivRqWdL/+ZJ045Tc6vYJ
uCASs7r5J4HSE52EBOzvUaBHSlvoMIEwDbpBd8NDGWSC55OxXgiwum3S7pYm3NQsHMQ6xW6T0luA
gH0Z2psMYZE9tU9eXS/AjvrRYwduq5QXdSsdtYhM0JE9T7L6K067toLbO353989qe9KxSOQ2xYvF
1G1yR19RwBrtK9TdEzg+Sw5IJ6Zc9ISrqpgML8Cy2K0dRsdanEJEOSBrcyGVgR6qQgw7yM4S0blg
3gP9cN2nd4QSxuMx4xMTr/ubo2LJdmgjUj6HLAM6DRlJg0ZqbeDiwXPKZtNWhzhh2rmfYdKnZbN3
aNp2s5h4M+jydfkKMbLX9n2Tk0lyCQPdTJfNmSZNfN8vLrUk1w4LnUvSoyvn5aLAU3uDAMPZ6ISt
vbWMjhAE9jM0B/LB1d7kVjkj9M6dLSLKXGRBC4K/XWFaTxY9av6Kx+/eHGOMd9tBOc0qGW0sCetq
cmHO3gPIgnIUIgRNilU9YhuLCzsPU89yv/e6q+KB4Yd610nEj5DeyEdjHESovZRnSIPb98uLoPlF
PpBDPrDoi3M3nx2WN3hhz4MOOM4SGTZ1J3L827jVS1rwJREHPStZQjq66wDhP2RQqod+/SNCkpFc
b3c9FyME7K+GqsusxDcGFGuBSkRlAv7OKKZpF1dGjet8WCKfyhn5vWsdLGqDVTOlbIzc7Ut0+Gu7
etv9G47iqCFQhqNbvrhibuoqOhHw6JshHcMLEpBCTNEs8W6jhRd4z1zpEdvrXmgRwS/JxTGgkNLs
ZtIKzK65assnA7eSX18LtJamGBMLBcxjpeEfRqbzoFN+7LDt4V6c75iSQPkWC4z8y3tBnnBwFta3
lewOmvZqJ6Ubp5B6bWgiDyxQI5czVAyo8uGephragcQcmjeSClUejvlqJyODUH3tdZuDWWnFP++1
EhxxmwyzeW6SrTPIwbRsT//eN2t9sM7/skCxfAc07joEKH1jhWidPL0ekhhsQgAVdwy84y1uHCYt
mpfvdaiM/eWX/KBi813muienbG378VdgsDH60U/CBPCpDPLhD46DLoaVq2sbRzj0R1zgH8yAFbG0
F3fcHMZseqftHRXU05luUOF1RRiLY+Lm95qsPlHLDpXNORXAYuMp5d24ylYO26aoxyeVu+TCdGfX
hMdADI15BQKngEpI6c8Z+Rciu5YCRaWOJhKZx+g9XC5kWyvrygFqg84iiAm+wFgMDJ77p8VtESrX
g8R3HQ/DAzh6x67MXtjtvBsL0bfKu/a58Q5VccgSGGSNuDv/sPXdTaj1xW7AYrp+x/liCOO56JTz
VvdXOXq/E0kegxnASJBCrK4WgSj6cN4qN9VYvOuKA4c7o5bzDml8XEXRq3YMPAk4Q065N4mpzbYL
34AoRbhYmH6gEnjs70AMu3o3eb/lTQRmfO2TUTNTJD9jEuX8U/UB3yHWtqbt5fZ5pYNnyRGqvcLa
ixb4Qm+JkX5qZdqfaBLJxAw5wNSKHmtjFeZAIP8FM7na7emHJ1PQDyhDtC4LMm1n2tMvYOFwpJnG
BEJUN2HNaLBBpgGmer2AQM8wXC4HEzd2IJiM3lGuqhurmE0PPcgmNDhGyjmfY2cBHGAbghBTnkaf
nwxQcEk0TeAoj0d4274fHT8HXUiitn15nF7CoZqs/AKBkdBOMI22pl6fQqHmAz5axjI9cu5vu24g
NyZZVZ1MjGTj++ynk0fiexgJPnZ1VMMGTAmXalJv59eO1hLk1dLztKI3yhZziT0SeYFaK4aqVR24
YNJfnKX9sdcIOHXNj0NY8/lowW6WQ/tG2jT1hdoqFBj71AqLVuv5HsPiqTY6LsuCXKV8VS1P5T6X
NJgSSyjVFs8icYN4osMsgpdcTkB0PMnXZbO0k737j+kd2CeoPtrq6Vnm7n/IxYM2yEGj/ebilQDu
2Oza37MJNPUYvYkSUihRiAQPvswutTD0ywD158IR5n3dUaT3y5FPXaD+HsvAjzKJOB1V4jXD9ex9
2xmVj3MOoBEvFbnaDph8eks1qGlEjJJcXRoMekKj92oRKNLdp/rnJPbK7Nq+N/IjTdvgjWV48ryr
/FbAjga8IPMja5xS1RsdgPIcGijsP5Pm9ppE5HNISDhsRfPRv8IruOUbK5A8a3Imsb9EozmYWnYc
oXPAytx0u/4T+nbwSZp82e/wXhC5iRSK8D/HISBununZP9nTicx3vTGg+8rmYSElBAAdzWoqG+2g
sFAC4sTRuhZPRVzuQjgInxpcctAE8t+4339610pI7ZiirRTh2hHu8ESt/3GkHvEaip6zaRiifY/d
D2WWHxXGfa30wTbqfvzc6cvM80jG4vkfLpmo/DzUGx78OJKZSqy/ERyNzrw6/Qk9LjqQWEO53Np6
9fp9UXIMGC/UOfs7C7jY5QsvacXrdiJvHfU/UzDfGMWYnwk/0y42fCl4/f7uavVpTCmdeyBVk2HR
HHFshYrmw2Ekf2sosyDowlHh2mKbM9q2huBzgHgz1ftvUu34M7fsLJN7ihADmVwtGIsIJX+ygAhg
98YSvHO3vVjTrlBraK+Zpn+DLOmHM99yOIlLkk1J62bMqG3FmTKhciSUujBwLgT4XmQRVAqF6v17
atq8gSJKUU1ORMw4urZaTrTL2M5GLwy3aPneK+9to8mB9g4ZPDpCZ/3XJpSYbDTvIOplrjjFtzCZ
vzNbc39QPbhTeNiqACyHV4jByGkQLt7R5PzgxwD5b1IbB3NRfiDygmnYRuDyslS6D82NrULHuYkI
SMDr4cBlFsby21ps+yGcPNtkZGVYbMV1tW3Xtjpo66MYlWzPQT/z4wdJWpIUdsVLIa9PQn6ukoUM
B6IqGbgK+FfCjZFZsBU2nIgz275gZL/i7KTMmXknCpaihQbom8uG33QdN18AMoa9i5VvlGEkxgMw
aK4WoF9hMA4kzz+Co70dmj7GG2JrnV0EzsuGCzNsOLVwbC2v670cXtIt69Qp2wCRwoBOySeh4hsH
ha0AcJsWPYCw5xZdHoE4i3BTsT29qI91tyCM7avFhoVXvnHmykWs4JkAYWy2bOom7y2/QfEBorvS
dgMTZC7UgqDQ0LI2pWwYqgAElsJLKi/U6LBBIAkePAFJK8C/TrbSDBsmIR9RWWcenX/modfc1XJq
FErjVzVTdWav3+ThrWoM4SGkN0WsYH2QqrUFm7sS+6xYy7jSbZ927+4TH5bnvcmT3l8eSfzUV0zd
Ov7Aexs7NLPnSjkZRgqOtjGzUu2Ct1AEauESEZ4WbHCP7RSn9UPOqWAfB8S1IYcv9inVhsaD4Sa/
NV4vGuDV2h1tvHqPez0PrbRE76auDlclO0bQojWwYW/G2fl74O+svZaFDeAF6pzkZEDS6wJqwDs1
1R4JrmHYpTtjSvHS+4YsMhi21DmIez6BSL/qE4QJGA4dIz0kVUQ5w1G2WngBpAc7lcVZh42XINYZ
8DBn/xgFi9314AplaP8N45OZLIKypHwoyLEHTKCLi/cs70U2PD9QN1S98h3ki5WklxjHaOZCo+w0
5aErJW/D+x/joiYdqkUipplRENFGRUcUsIdtyPBGwTAQPaqUcjNUID6MVMKp2+/BIj5QHYIO4FnD
KcWIiNn0nnqKmb6Qc5PPYhF2zt/a5VVa1ZeYHEK5iYxRT5XJTdPtIx1yxsEhIcby/HBn+wW22fDU
zQDPsIIpRqkY3NjcdSfHJ/glbLD01Yw59Nr7r/t+d9+MxqzBLxklrqFR3Cf+yqhSJXmdTcy0AdLA
C4UZpj3tPR60hgkKj8z1kCq3WcULfMLZjswHXiJ9sNWVz54kxd3h4LeKJOOYAbBE4Uth/vI+1ycN
oRMrD3bfy6wLwJMZHOPGYzlpsInj5oQ/85E7JYK7mYJQWlC1CFOlrVN4ZLmXVVJU6Srp0xzaKbu7
MoQGqL1bArxOoHgmkzmNoSQX3eoupf7V1aGfywKysl7AUebGZ/LJbAZ4hfFOBvaCb9eZcEYFKm5a
BAogog0bMTWy2/v0ko520tXaynKmhV+3JpaGI7wzRXCu3sk/64qBknTBaCLKtyQhZGRaig+BPrTo
mamn7AdOO0YHtcTCgyIS8Q6Mm4rrBXnhK3FZzLJzJP6+hK32PZTSgoHJ3EXtGgQrv5GqKOTx9fLN
NN9gpYo3nowsUJW9Lp37lRtYpkf0B03eixDHodY9/r7TdaYcLNGWGXjokfHAQh2mNc9tUo4iYJ89
b7/YSzAdkzHqlrB4sycBC/GAKfDNg4XCU8IZYrZP/GNq6cZaqydVb3hssZcPQ3VkhVc7eNb/5bTa
KW05GrbqTFlTfyqubH4TTKZGTNWJ0xlsrLm8fvPKU7qfXwkVVbCO6xIRrjd5Q5qxJdKL8BhcAcWv
3i5Qs7YJFIil77t6ANnQ90Ux/pDOjgNYy5tDFL+UYFUupb9x7rgvcWBFwXee9eMRwW2bBOrAXidY
5BQ2jDTy1zCwXGJ7ejt1j719RFbKD6+rxiRLGKAuMJhcnfuGbX8e5S40AkqiK75qcK71tY/ISzAi
97Ny2JRZDT491uz8Zuul1M4L+1NTQNGeBJZEO1GMXWdIQ1BmnoHOiGmxzXY4mLK+6wCBkrjKw8pt
3tH1+wgcaUPe33mW65O4IIhNuUIMkWjCJ7O8UzMdpW413obqs1tru/LnfdZvAJu7Zggedg0WIqAP
iwlcVUkDgcbSEK/EhHVYKtvqI24PlueuEnscn12tBLKIv7PBV0jppIQ3n1z+i73Klp/RvLqheoB8
cdIKwCUxANzUprDWyQoHn8ox2NEgiqU1eeuMtfYiOXI2sjSJJ34qoLim/yI/JyS+OkkEML1q5+9f
uc+bKLLYXa6Xztv7MuKYyXroYRQWZnKO1xsQDAHf50opxW8SbTFw6ltWJKD0aPlORmu5bQewAI3R
JiHd8gTRm+kTZN4pXV//aov8IiEg84bKUlZfM/w27Op68jh2gOxUanvo5LpWgEYv3P+nfxqSMoR2
fAsyyKZQ4uuCfKMuUz/HLnLkHym+wmGO22gt7rbrM4ggAXfrSFxhpNo+tg2/fZB6/tttodbE6WoB
VkYxYYBFnYMZm4GUtCWpfjxJ0cPTiv9kNNKGljV/ivQkT/CvPMwiJ4/wQUIgGHwbZKGSddWMgOu+
cNBDLAIsNeKBMbYHR2ZNrbBq1OHvMCA7JTE9lKPjfv5ouuj+zxyICXsToBSE5v2z/GuuH6qUtVBQ
icDbpHYXqtEDI77g6AKFIbAjAmmI5tbGC/B/7NGa5Qobgq8FgQBOd/WNR0Iye0jOvfXD7Rwlqvt1
TURnd4FLjjGo3eqZNmOSzua+5db/mGbKR0xDcJz4GTGUXlk0/MRuD4RybALX3e62uMg4PIhmChlO
tBHwFpok8M/FnpELz6RXhLR8sUUbzBKncjq1w3tqJMQXdoRhjP+LfCAeiP+XTrLG1sxTW/PYXgdO
MhXO57Wia2luOIImFsWmKWAFso24kekbaMhD0kHdaXVrezLhkJ8aVaX7MrR4SJsJ15YDRn/WGuBK
uSyEs4By1qBBzh+HwMXalx7LIIKAIL9B+dRAK2e/PN0emQBOgzXHh4M5CmZm1AhDI0HmN5i1hqSK
XEAMOnVPXR+d3i8VBBJT/RrWBfS5N8OFIunTv8tj1Dd/BCrcRGNN/+lwo+gwSWfSZ7HRkRVsFrj6
oFz0/5tX5sEkpZ+yu/wBcX9tzIPY1ptllB+D/OQa3HqPJntqI8Vp4m3x+pMQripqHxWAbT5RgEiD
SuLUWCzVWBDmLlK85zYyEr5Of95E8H2LC5/8vCzB4WkzdZfNRMUDY6yWf8WIJZ8DWMaF3PBsZIkj
gGpFZNzglMRxB73OsCcxkT8w4TQxGf355hOlo9xa03moNVVoawUWPTUhbSv8Y4l8NLe37U/4Bhb4
AB+IOQAphdsEIiK7ODCLSpfumdsP10+uBoahUR7aagVPLXvwjHeqjuuXu/z5dGn8C30gxOuifOmm
EMMxr/FHjRHWzmonaOwO45rwU76F4DO6wgint18nRtdHK4iJrtwZTgcXcOqBVeZu3EDIuWKpjOhk
0H0qB8YqMardioqVZKimJe+z1qUI9rThtz1SBcCuBvtWNu4+o9D2zF0J1xMkKmqf/F7CruagBlDQ
Ds1iAZVQG7EJiGn2VDBA6tHY9HgsMlodI+2eA3njPr8l+i06m6LPOYi8ceo/TND661PqHz+smeXc
ZjRj8VGVCCQqZPEjvyD/KZgL8nEUqjyegP7hHPCiXoY+at5d43gpoPi5jCSX2pGTw+8xTeRGOPn9
Xt9rjywpZ4o8Stli58j7fwGhM1gZPffzsSktNON7XLLi1Q9SuJjaeoVCe3LJxtrxl9avNjaGTGKd
YSsqiFClftp8o/03wRuYC75/bAJmJDGu+Cz5RYl0xgO/KuXlKKsqwj1sOpo8U5ktPaaB7Cpv9D5N
M7HAgrIWD4UPmlsvuyN1IuFqL2aOtPiPpziUUt63LEAG1r3yE8cXKReEErCK3wJ6MQt7vzMoH3di
PTNyAXH2OTUYAknR1uim4haDc+530zTm2azIS6/4lPxVHdLlZ5rR1WUA8pgs4acqJZz05DJtaQJW
BGMYnq1LOoTtG7cj249wmyA30JfAXno0vfRM/HiEktyY82omt0uEmb4WiUnh9xF76+HR1qH2twqZ
7TQrVN2pgffsR62UOGf7jN4ZCfKBxpwR7jnVL7i/2as32MlA6JgrhXyzso6InQuTpzKgqszMnkKS
IGToS4zWi6XfwtPDC3m9cHyFUZzpB7XraILPiUdAgrPFRe5PaTr5HMONFklUSJQjN5X5E4tVlpyH
QvBDPe8Aebcch6LmgzaO9RgIKx2NRGlnuSau9GUkLCsVTHMF890TiEOEn4qrLTewe9PshwTeTYDy
B/43CoVY2dBwJYspdG2wWN4Izwsut/IZh1itf/h/RPnh4G9TqCIi7DqemkVMTxwlzXUcmKrfPcyl
NZwsMqbH9rgmXiI6egqETh3A89Ox/WiUWp7y3slCe3b95PejrNzm55D53a953MEkQQ2QVhRNpGN1
MclRx2YrSnWJtuPkHglfnRmWkTh8fbHgkcpW9QS1etHDEeHOvTi9Cilf+6/C1md/OMByp9nup0lf
viRXlNzxBOK8o3aCAgxMEcop5SWkYabi2k2rwAh20CrzE+C7rnuzeQTsCwLlL6g0On6KDNqgg8qN
+85b41hxQVVPn06uo3JY4TgnvhnL2foSDIgoyfv4EsgR29VdzcqeZqP6IheMSP8kJmbTpJIIwKjo
QHNEuyEl8hzV9Z8JX38C/y4Mhwd2FImOvdgcGeRm0N0cTm3iNDPn8Y1f/of+1n9jqvFUIHLXALTd
JT0J0BlfLejMg71FxR1BWAx+XTJ6WctZjH6rYAFtbWk2TPazfP/tH9QBrtzGnXfizNtvgiaLu1cQ
jaenU7uIKELonM3xJHIezB7LQwP5XNVUYkykm8RBmOhgREzHL2ZerurU0tPc/rH75eFaruCE5oac
pXST8OU6QTyi06SEQR+p7nFgxThTF3JPOr55KwB7bu53xzNxSl/4MgWTCfa/PR2gwA46rYIun7wp
uRMMyoi6fimHp50UheiAQ2Il4XU0AG87uMg9rMA8F9aLI1QcUAUScRodMDyG+xgb6GsAYUo6qIXy
KlcoZ2mTBoWU2VE3klBixg5BbaXNFCr165BYIM6j37+K/XeFhVjpNwy+n6aL25AB90sCx2RoKJUE
RSweXZgX6f7oGS5cHvjEJFwjmzIuROaXOdcfElEPq2oQmrYbVb+ywlEkkIRdbOn0JOpRhtEa8JGk
FlJOfg7UgBhyd6d51VRWbNFnKrHKiYDh3e2LRWjZBglz2NWur2xOKM8/DaBCHWMzGse8DfBRlHZg
boi7NoWwxxYALAj8LkWnJfCBJ1tPFOx7HPdcOhdB+TSozVDEt/LGkKEfinVxBIsAnrJZxfJvGlfe
PSdgTWWG9CXD34CsPzTazsWFqeq1onX+FC3IeXgcD9rWndIvid5N17xPKPe0ql4YOVZf9/NM27N1
R9RmvmfudYTo4PLaTB4qOiZQ3rGZIjnaW3JXaPMSO+IThDzJDMlKqc1PGgbdGPQvlxyCbhBgaA6Q
IgVZq14aw8XRP82x8Ywt+WUBI1KDlCVwgTpYOYWr321gPD95xBXyHWyftaTguprqLC4ur4TRpK4Q
UYrVIAkXCfibxC8kK3749/l9CSPkBFRR/JFACx3r5XBbal5yXFGPQtVrz40YdTFrZbPO7wDerBVh
ogm4nvS7AP8AYHch+k3OYYoAhflbcJFiGB6+WuXtJJkfcPj6z4z8WyIMUEJtmJf97JsX6DijShPn
crEmlK2Cymxome99mpWWgYXMgPaDE+xbWQvCjyrgF8zJaYyLeWDTT7PuADcc8iNtd+aCoBwrOZpD
URLkuTN6fBxYzDw0EQ7O8+71hFL15FSGyIYAhFcx9EBjAInmwF9GdoAmXYxlXSl53X1IRK00WrDz
L1Im4tKl1rWsx+l6TaZ2N4lUYSz3mHH6JP6pLUvfLfA7GgUtG+JhPpdE1xKihkw6Cak4a+aLOLS1
HgDVVXEfh80wtqqaBw+5p1CN0/4I88LoKkI583rt8EekzNb7doXW01qO0CiuhnHCkT9vFLtEEMGY
y63AGnJyCO6FP+lp2/IYgWpabRf39sTSeDki+AlT7BjfO1XdFsX0JQFpP1WcWv3qKEQSo6cpM+ju
6D4XUV9zUyH4NQMpBpW243WG3pxlVIIKqktfedLjRY/MgHZ9dXN7OHF4jk/FR6RdPD6CmZLdCyzJ
IL10cpmtHQyAyViPqFh0mru/2bIXsxM9DWwVxEXQMxnFLlyvNH+7Dhxk1oEgK0ap8tQxvnOsdq5X
Iq5ZSUyldn1Pw0Gc9RYLaT4umg8uloVf+IiQdUOKiLdTStL+6DOIWFethp3t0gKSLcQkhlvbIcJF
onzJXYOpSEvqX+hKWk4Vts4YDdfT7It2CuQFkYadQOa4fCg9TcxGuQWjjQy9gZFAe2iLiGbaEwao
/nSiLgOfvGNOujpdoAUnjPK8ZP7N1NTwouwkeq59J0bUrVpgzvCdhffTpuwxV7+p9WHBQTFPWhM2
xouz1ohrVGeQqjXKbh/rWicRheABu539FLsHt+O8cFWyaeiUztMMBzYJnHSa0vJJmSiDl1siX6aG
QJXkZtn2yRNr/wukrJN2MncOgfiljY3/BDDt8Kp2m4j991gijbmDlqF13tCdjKQWOd4MnWUV43mP
Gj6Sq66aabwlC3OAUa6UP7803/XerFj5zihr0J53lTyeJClgCpTScd1IGDm+RZn47ApnbOLCxCBq
G5EwrlxLxYeaqVZuBAk6/6E2PgYFR+TBe+VR/R0rHUEs6fFpdzH8tTYXQK+ELR/2sgL9Znlscs6G
GnpcAUKahs6xLEFT5DsAfFClOkXCC81L3d7ggYtmg/iXRDsurJ+mF/44x45bgd/nO2Lv/ox01jRW
xJwnoR6hlsVczyLtqzXz+jdFUov/GITEOyZJMjvYCsDiT2kworC/ln9+bGmKt2gQ10zG7aHdjceN
uI/UVoZ7j1prprk5mShwXKN33i0hIwrBBcAqmmKigrMy8d1lod3gcLL1pX2QZP4IjSKyxu8uGPrx
XlJwYTF8JJs0N/YKHS136XMTiTVhJrwVw1VbA9YJnhatzNEXLsTnPjFinXo8BwTGiasmmsMQas7o
MT9ZEpxyWBWHghhKBFCIoAJ87cCTtwXeS8XD5rKgRjljLQ4mQBPgaGKWCSxwGUi803JfHvGhbAj3
ekkPTDs1FULQd/rvuQbXVJbCghL4WJ42qEA/whFyINyOO6L7KAH7w0v5YA9iXeqkO+hdmCxrriOU
4/0GwhyBF1DYPdxUNI1uKEmrSVVo/q/BMa2KgQm8bfxqDOKtfLLHpBIoZfiWLlJ/RpTEFVl64s4g
Vy0gX+yvwofUFOzDuZt0GFl4+fkmTCwn01ry/NUo51gD0QE1h5PZ7kG4CO2QFRkOZSaTaq+yhVp4
GHQI/GApU7T7eXjy/JjjdzLNzeAh5w7M32LQthQ+KrQVu0RQdVwnrMA6Pe8Ik+OV7t4SQ7RiPTWZ
eL+aix/f+nugneisKQ7kJkWgoyVy7TfJ04xFvksRa9oNSeDMjHLNVlsapsL9JgmgNSch+IeRf3uD
/JgbxWSD8MY7VkAubPHs61eYyECT/Zvo9zSCjfldkJi3KYjM4IY6oORmndab4tTCjwHDD1rr7wMF
MYJjt+gI5NWqrtdpY4qihHVQdxQ3PeHILmZ3IyXS8l/Ify0nziXLZXbnnjwGi4R9c4O9dYJ96GbP
yC/ELPqRIhzREG5eXyquxDSnOT0tEDKlhOW+GM16/llqHzzr5Rx17G9MoaZaxV4YYsvXMyxD+/U+
WnSTJN6Pp8euwJ7CJEToR2GaouV/Vz3wEn1eP9TZDt/Q7Rk1qT8Xg9HbCeQsB+7j4RVUAQ1AGX1c
wJzpmbq8M94gxcXpttC/d7uqgV74IGcDszca0Lou8J2lionVu07YVPdCwz6tiSrUMkFDta1oOPrX
XJR2DgymwDS/LTR+h/1K1s5r/Hjjm1qQni+Yj9C3BF7GesNzv98Q3JKubkMVfqVM0uA1S2ERamgX
6L4b9Km3wUdTXzb9GB40PQH2GgGImeEPjeqXlq8KVNapcXTltTAFE/SSjfKNr87sHFKV9JzNKNVG
Mx8OXZbJ8t+Ey7m1T9CVTkY7J+3UY7m4NpKnSZHwMUlEltIMXscK/1A2DTo5fGScD1f+hV7FRviU
Vs03pKd74nbQx/Prl6OVEnavvsstJ/DD6sLmPLgCzxzSB8UHoWrPYE8Z8Sw0kcmAisxbVHpNzP7M
MQst1928M5+YCM/4+GgJTb4bniA5z14W/7S6o0EpiTKjcK3xvTK5SXGGtYFtwx9BjH2msbiegY4x
HfI8EyJDt7ImLVSh1AHre19LeymZuL9D0oMRqHUmLM2kAKPCqGMjjAzAGqKiVK0oPjQxjExhCUME
35pnOh/080luH8SVk1eFzYcccZZOxb9fTFOHxNv39aGomWJ0NrLkoOLt5avGjB3VkyigEkWkYc22
Cw8LmhaJj3wLI70h1PIRooVfMgzVbqOiP2ldsVYBmiHtxNBF5j0fmADSAPmlEH5TinnpCn9hQDGM
nKWFWOic3IuDFXHTNtb7zwgIPT0Z50gCg73VpUcZif6rh3t4+lKESBeEJSjT8YPBB7qNHO0JKtS8
IBnkrFVp+f1/+p19/BppqxjOCqSy4KzgCHlYwn+IlkQ465IW0W4WIaFH9U5UG1osD1lLDmLERx7F
MjPMMuBL/YHSNMg6nEVeHHW7VcXtrJSVIubQDqYaI6whpIpKERAC1BBwCLV8xINL+twJlqevSaHt
0Mi3qgmmOsgkpu1o+9jA3BQOMt2d5nXb0TjasCvcYVJ4zw+vi6+UAnYbF1a2pkZXJQSrXpivNI7i
IjKRKXDVmYlmOD4zlEorb2emOYWxBgian4Bm/KEzSq1mazdV4z5vJZX//Z+jub7B8IzUe3t5tR7G
DlczOOR2rd8AWrakwGn01VBZMC4lYpNxjfxbgUEUsO9GuOknAFGV+4qKq1mucguOYwNJ34vn05zG
sdMV/lVpMy9n5IuGASUbi4jXFv04aOiGIh7JvxDudN9iwUnP4rLdm6kWvnS96j7qEjN/gooPSaB4
mtA+y1kBgZqaqRDDKaUTEXnVZ1geFrzL0R4wmjmuN1Z/4OWI7BN/ZRbUIEKx28kyHLmAsLcTbbWr
8cirZUIqui1whNMg4AMz+oLuYiiVredzaTEGBACJ6jwa35JlrKHLtcSe+IhVFeyR8Un6tnKESDqI
ithDupPA5lw4pkbWiq+dVwhiREwCIN7z7TnJbhf/AdmJet1yJhPhIVjdb5qjajwqH3u/1kH3fCmY
iZ061kn3dBZhYugkp1kbEbPvC8RaV0s/XOoMrDLP4Roc/T4ES8DYYpqvQ7h9Gf29T2Ukye+bUzwe
KDlAoO3WqKHfrpOX0ExJOGShGyvJ9klNrUgR32S7wayvJAf9Sv+hcQ0wJUPufnho91k0c4dfYd4x
CUbAcX0ycPPulJ316kCvUFqEZjAmTBB05cWz39nqRb1Ipu9HDWocGZ4muLikkubE9+z9mH6eNcnz
ABpflj+HhVbLmyMHfOmMY0EHwyur9qyEmvzoFwU7Ylw3y3iv3qcfRo3m7PvvGv4x8Gugfukvp1eH
uilOVtmBrxV07rILhf7IiPnwY8j5HFlYFHAagfO0nYaCz0Zfzy/L7JPbOIQ8HwQMRJd8qHW8rLRi
5ZHGhKHPxE+oM9l4QGPyc+FgfRUQ3rs5HK4MNTMbkTMUbd2attyh93T8nAupfNF6mdD0VwUmNXeh
usGLGg7JSHTw35z9qXITDWA0eUcsSPBQ5U/VjWBTh8yWQ9Tpkf5Hns0TfZ7i0jX5GumVc/v/OXjK
Rgeb48aW4sCT0VFOSgJrONl8ANbbZ54FG5HiJ7Q/XuSWEZWIzGQW/kEw0cmiebR4FEeiyfIXoiqx
apxUSWmBqCC1oN+HspvgriU1XuX0aA4FkgAb+Jfjqp2A0/eDv/1WPrG0nYOzAh+wFoA4DfyeHQZk
ebSgQjmRBfcRWt29X04yCWiqsBiVWPNvjCMHDr+UPH4LYkI8IwtOx+3TmSF0ywgHH9bmuA0iCXXv
seVLUGNuRCBo+xlno2QQO39CBIOqmMW5bB8+a+DphzyxMhX7y1p79oJWiJhDRdFNJq0dP9CYpwbL
17IVeGDBJxat/bdtFYD5K40BR1Ht0lKuADc0pb3w80crg6J5cz0rJV1HN4fL1MNz3Kiie06xJ+JH
zkmq2tecV1JOpIgAQ4rAEho3IDYfIyC5c3cZ/xPgQtwUCx3B19BtsqCr+VPzzb70On39q1QJO9Ut
D14w3d5FdTFoyEE0Z4UQ5Y4Px5ls62BAYzwYSKRInnQ74TbdD/2HbsgdQ88XWutRhbV5VRrJ9FEC
OMRH7WN3ao4ZTU24LXZbZ5NzAHATfU24+6pFUlDfWTLi7M7jIx3WOVelQ1gndsRruMXRqF2cm/Z+
ISBA4GIwH78VaMe/zody30kCPusSF9yUSKrbtJVkkqJNl86cnYbnN19o3F62HNKI1Rufk4H6qcbL
YafLwmvNubFbSZs5baOX9DQCXLXyG2HXMcOUS4n37Sgqq+lskr5qzXGZ3KacNll3Xz4Jiro2i3hw
MzmMGGkplFY2BU1486NkNnkVDVTQt8Z6LPelhFhf0XhbGLznb6aVfqcqi1fdK6x3P6umMHliKjdN
N8R/X9aMsbeQ5ee3Us6eE1+3suRqcnczOdecMpN+tnkL6tlCx43hLw1Gtrkxp2iOED7lkdfZGWXJ
DGGLkPYgOwwJGeUjTfFtiWRyl0lJoq8T+QsL+oCmzfLMOrWksxk66TzsjZ0YrJ25v0xRMowU9K3y
WAok3H8YScaF7E6GyrcJvGgV3CzauXQHAK17OqgN0nXNc2my8LkeCtEUfckI89crQk4tjZXqIXWi
s+VNMr0XH5vxASwd8QMK3rWAGmC5IzXvEdcqm0vl8N+dUvBFiR01IT9qdBvLQIIXjfQHJh/cdKwp
K7l3Eg3tmASdKgejp04yX9TinSxVZsSfDI3tCApV0DWts0C1n74naxfb4kPvScYKR5a/xrSsjay/
Bhzt/raUNRPM9VuY5l0yWTJ6bfISi7AFrQAQpJ9++ApEcZY/zzT1n54t/fhZiEMOeAolsWy1ewJN
euLgU1n/ipquVQGj5EdBw0XV81yFGe1wSyfScJu8+Y+1WFUBiyMVcGrJ5TKccEgDoas5Fg5gartP
2E6Y+qYzoHsHHXsb/OoXgtOnxAYL3EoTF6K/e3vIticEw6kvW7wAkeHqZkCwrKJsYkxpdWKAjOaz
igW3P7N/wenJHS2nX4N931Xge0yuUixcsXQfkNPLH8mb9vHkYnQK3gycrWnRRTtFz2nWVVN7wrKk
AJxOTbCljUGLy5JiSi8Ik2H3P/GTX2997AaV7DMfQUXWaWQTGmEgOyqp0jzKejwPuHL2V3Bi6nhn
Dd9ioWbGsOGp2q/dMGl4W0a/jyj6rkgxI/M62IoRCCXTMpXQgzh9cDMFHmIkEQ3MEvY1ww4GbR3K
gCr/VC8EhrPJhgOUx5+60MrIhEuqe4M0NSvqFyDkN0MdHwVqW50Z4X3d2HzU74Uf8+bqvsfPLCq/
HJK3dWd0u8DoToHs1D+u0fh/BrDg1uNhhNeJKLgSkQEU67g2oNl/Ab8jgThTSWkXYNDUFE+CatO/
gAwDcNORb25G+0hdvyiZRkfzmzmM+5+v4Q3dVRz87T2E3h16dEQGchvZmTA42u+fASkoVJ0brLo8
RfTLH8SimcJ5C7v28Bhh1W0KkgAv+PAeWTpSOzuAuJtag/ycw+M5G9sgtlIUiOx4z1viL8rV+w7J
kQuvDP4ULBYkSNCsCGAuuP6LqOzjiaSCP4dg43ER2pf7wmdntD9DlHhUUn5J31pjzirB06/sPazZ
+OgWToG2CaG2/GWI2l9QjpbFsQ5GYMjTWINw7F3Qlh38NxZoYooYHBEb09wCA/whZI1+T75wyF2J
6gbSZHRABDYbimnxpgvK3+nEG64NsjqKVnflLwltWNWbXYx8Cw+hDZeVRODnKtGgRV1GVg3X/9XN
6x7oHidXYmEDp5SjXEJYJsLsEk4sahCe169RTeWyhCL9t4/pWEg9EkQXBCYaP/dRoxt4Dqc6M2fF
0E2RnpYBcoN6MYx5Z5TaQ8YThm55Etg7ZuvG6thQlokMLQceuwQO40SarpHRHvQaJRv029xwYQf2
0+859jPKtngDfpe4mVVzbWJmRnTW3tsafaBWSYMlYKlaeK99JwYk0BNQZgWE8Ed/2mdeT5gxlhAU
vWX8boLx/wjA4miZTsRSkuvS6wUnjKmGlSpoGr0qe+GgpdB1pCoITo+nf02/lqtE6EmaF7zURokr
VfWElrJ8BmDNsKjc9b5EXXsaDzx82tjOrhNkckLz+oY3jsC37imzKssfzrcnO5GMNKyrzHIIaXfy
00ErVQtYD0KqecFo1vT/SsKBAoucqGXFKWG0FQi9cr8EOX6C0HTarWhWZVKS8ml/uO1yd/NobOpL
Cj8JOW+EWFE4+uTdz50kkNvWWq+iwACj601NN63v2AlzzBCegqihWnfXgjAN//hYL3k90dEbKVTg
+Max/EnKo7cZKwet+L9dNcVWr1i82oQR5Wr2V2i4UHBS88/opiLloB6N9kyhN5rVoEYBnVE72RXD
kZUl7hW3Dnq6qPgvZyTcpSylrBYcJTK9M7JEmoNdkeY20f6dE7UZo7RFAn+dJUH81sXE1xHaEuDD
auNBqpvswNWeh7jWCrs0ZQkgL3wLlE3lkgRmcSW1CK89Qzk700ORRblFikNlxf5NMFYK0YEJY+T3
DKTdT+/aNCpvE788dO4Ec+Pe2v/W5b1Ra0joBXNBeKGKWtP+EdCENFLiqIC1Sc4/CUS0TuoSzr+e
g+Bc7IttFjK3+pl/HUhKkKAEOKRvrZi6D7md90aQrwkycS9omVc8Vw8vQb1HLu0lFUarXSAnP+X/
xSX0cPZ7oTc30pmlnWVCBjgwl17bBuva5IXSuKthEEnrxlsUrJgw16cKgmeF8fehCjjicpBCeUGE
Br1bQrqXFNiM5cUrGO0MDV3+qe/j8cM4uxygGMRx08WTipiKHNtvYCbo1U6WXL+0Rqrj1vceaQPB
Ev7bY/dOx/b3K2EFDKqR7pp7J3QWuqeZK4MwxsQfGiLaXY/k5fptkI0hE14uBvT2mwmGGRv90iB+
E3zkeBoI7uJa4a1Ni42YU1fJAlVXqkgFmfpufoD+0Xc9h+/ym1DsX1Id8/DBQ25pvD8pbDFseuvX
lNMLnSWtEiYXGkJ77rUbTYhQxC8r/KtXnbsmwyW/DRO6rauagPAxwDpMr9vofKCsd65zoprUXxTd
11dXDnkR2x5sHSDLgCpdcrzJHvyAR6/2+YItqeaWmdyIT5CKgA7PXSzyBQMUzbyp34Gv8lQEs0Z2
74OtEAZxul6tBW2kMmhAvnf0H+mlHtngiuORcN5USjhjLaGMTFo5dM+83TIjVOuBn1fyHuNo+qe6
/m55UFccJ7MTBqzVm+si1Q5i2dfiCJ4tru7Qvv1WRd0lxhdnbmCQDp2Ar28HQhExsikqQg4xL5qW
+zKVJLSXrQZs4LEtghzQw/YO+gxdpwGw3l6UxGu/peUiL35hZtbonxnwhizn4oN6u5ZHmn0xWEbo
iPS3r0+oCuGB2ndyP+gczMQDzSlp7wPcVp05bImEwKGKb/y4zaF9y9R2XPqL5k7ngfIM1/baauli
UHGl3vqUSFbYsGpJsh4bt08t8/cVrzLGdR7gw/yGaiHv+vEUl/fns87w8GKcyRElnFmMBcuSQa3P
HRR5ipUzcKo4BqLk2cRtSGsaFiZYoh4NLKTzvpB3Fis/8YwtNgoGhIp4C1orgDEecOykOHompLLq
kAlVrEP+GSoajOqkKwWrtED/+qTC+jOZWaulpOTyQFrBVoJJ8ZYw+39BCXU/3oPoz/e9hBxa+OS6
ADQokEqSIklEMphosvGAZDOTX1EzLYe09UPHZFR83aXp1XevdCfmTPiqQurktFb/Jhr+P6spMcNP
3yb57NCWikgltLAwm6RMgbLQQTwlqbxqBqle6+8r5D0kgFpzmeHAWapgFQVtwVJyBWqa9pb5lWf/
VB1obOo0ZgFYxhKHJ/52HxUwX82Sp5sH9Y3bUCHHdOvivf0LM5ppidWGnk7EhOp2Q0DIlPrGAkih
4Vx9jfJiZgZFRhkGgDfxxhe9tWwHXKh/GD/RFiz5tghxbCZrPX1tEO6SOd8dSgQkhZ5Zb9SK5QAc
fdbUaKLoy/JNDGeoDpozLlD4GKajBtA1xRU/Cn9LRboTiwVm5uRUYoUpvG+TmLqL3/reWGQJFUd/
l5jnnuBfVmC4AWE0KzxYFKJap8UTH73anJ0p9PWHQmjJR4HQJQ3QoQdnyN5HIRVy9cTK8iLdUyiI
4eqyHriWeAM+Xiohlp/rj2gbKtnVQ9LO+ANuk9ipjkRHc8y/Z22whKkj20MP/nSBYh8U+3qaRfzj
SO4ttNvwP9c7qgNB9lMkG8J/jbLPc9ooss655EABK+4kK2stJlcUBJnWyBIB6LmPKkAZnMjhFokh
b471An+N6QkaPYN7DAr7lZWv2kL1RJNo6kKK0JDfQBF/g4WqJNzzfeQBmq+e6jvApnSlForhMG4Z
KbKuMt12uoT7s6O2BNn2Z1neNPecikXLPCbESg0vx4AMMjaoajft8Qw9PjvoNxExl9KhsUCGbCpq
KL0IqaDNRchnJK+32uml+0YI7G89B+Ni0BOLlYSz43H+KBOYMaTUbmJ/bV3Y5SK8YiVLIYUifvP6
CPGuGAYD4EGTVhz0GKvyMlctYAXx0+HiyEwyrHPP8IvuXmAB2lxgflZGFoKElocMHXqvhroQ9xtJ
IPFuAHjzTfxhM4CWAeMYonOo4cibxyY/PVM3kbGmyEWCtGpMCJUt0KQ7p+OwxnpXfLHzE8m6XWBX
iBs2y9KthKP3PE72ARVe/d3sIymJVdAa5UvZ5kYFKoynm1wtQnH6Wk+ktvEYtte3/XgvyR1JLC/x
iUTGC69P+uj+RhSTZu4ynbe8huf7/GY0/Yu9y1lv2K9naTx/ZwKfbvn4uOdL0V6nX/KPnsq3DO3r
lW6GofQnF4gFbZRqseLwX+yRxdjhzL6OU+vnSFRjKm9ePj/HCVySzcGl7xak3c4nb8jIW9BmLoPb
UDNkf6gZZ14JuoiWzSSlex9LPZzbleFe6Uuw6SNj/tuicU1sZuMmEyMNE6R9VLLe117a2PbD7aeO
0y2hgHMmoY0V5ETBXBGny0whZbC2LLXrxjFFSG6kXufbMQiXOZBfa65cQMigC/8TYN5wvpOkMh+g
a7PDQCflUTg92io10vhBQ989PUc2VKjyox0IofQUBrmYNOLeEcenM9ImK+H5LlfLY6tRWxWcaBJG
4UeUhf6pvBb8pqCmB1Nhn30LKV7GGinFTXSqi5ZZp8TbG3SZ+Giiyjs4ltKCPxCYjv/SXP6ilYOf
8SSVBF9GOJtCPzGZENMgriju/VJkzul3J5tYorG3fts9WAtWV35Gx6/X7o8foM/NpPFIY3ys3huw
i4fyt1BCj2fdSU7j26KRxfY+kj6B//0cc+EesVbzq6HGqTtLbSnuZAidUox2BbHvUbtoMIX/DVOj
aRk2vEFG1wFQafka6Cxj45o1MHF+341JGH5MvOkzKR47YQMuS34x/zoCdUIcnYBcaIx0Q+boX4Ft
xgtpKgZtBkHpL7CDvpCLJU+75LUamCAkqKR1cxfB7tb6FPP7jxQk+iyB395+VGlulLYtNvWruxGj
g7k8qp3E4NvQ1x4vonZ4B5tZJR/Ds5bQgac3XuecW15DcQJln6FrbO+oSTy1dij2F4sffbDiXM1p
iwbY1YiQhhhhJFS1DdqhJVdIpk+0Vjgq+s+By2h4StIgzEhwKiFKGp/Rq10B/COMIhmk/yI/+nPk
SwObjLVupUcB9gNtmaDMkOdekDfiEvYBTISyEDngwYqgu2vqPDJW08kK+up3sjLFIXQwXZxE3s8r
yUE9IQdOlFKcImaFfuCfKYIXx6Ex2gIwIDt83Q+dE4NjYnFgb1u5p4yjYJ5Ie/K1ug+rgx26w5NJ
Gc3oLLr7H7rYRtsBpHBU1EoTayiMvmN/SIvVpno7A3EhDHm/M58+gzPzNoYg2Ohl8dDjHrkdcFSy
IKxt2m3IF1Ww0vMx8PLOZUR2pb5f0F0hD1aj327EZpb9KYbGWO/C1BwlQFe4sZDGxpGSpK5g3yeZ
bdTWbNQu3OBjoGp4Ka8YPgQVZWRgPJeB0XM3TMtnH2nfU98PD7wq1JyMLjUSsr0yTfpwuVh46/9l
aJLzaDWfWuXDMwIPl50cq68hOE7giLmvSaQA1aVZbmLwa0otxx6Cm2VnkxmhFng7uNTBox/Lnnfq
4hBTSI8yhbQvHomDeAi0V8sKmAN4OLKZY3nJ36y6Ul63OdxMzSytQKuaIKYu8THqf91KbLfvQe/T
MM3zqxBAbJ/zHeQEzgjgm7smqbgXJctic5A8NK3kehcs0OZT91jWJTYK2XBzYEkMpTRMRrBqd/2h
VFTpOAhxXzWSHlR6FD1SEMUfZ06t01g1kxrozf+r6IM+RK8f+PDODly4ilSxvxzQuJQCQNGpoVq1
yUx3Eo6hP93LGbzDSuvD12wfpF7jQJFBwYRR7y31yZe5I3OhrfpLcUKFql26xA6/bNiWGlZnENhc
XQ3TqW0Nqdr4PWQPUaDJ0JB3Ozp1lkE4/I2Er+sqDTSAyYGquaeLAnDu5tABVV0vw7J6hwd40CGN
KAIsKqq+GxpgzZ0dP+qdN7gX75/uN6xX1AMsZ0bXdEqgkxONltZGGaX186XQ2ucUmr+eXogzr5lI
8SSq+TD+CcNzrz9YS90pkz16pZpm3dY8Di3YBLuBlR3xcgP0+TIIHhSkg4JE+TkARZh1LSNI4s6L
Vqmh0vkfxekTJRSHbJ2pXRYF4+p4Akh3eGliwqnJscB8afX+qvR3xqNqfhqxyCg7Af/jURyPEajD
ucDE0eEQXmZpbPK4iwaTHBfMiiNkw81eJv+rUMujFvGVE3kEZD/KIm64kMMb+jGCTzKsdLvKwc75
XV/eBKvSRHMAXRPx8+cOLkwp5D8gwcu+4IgLK4xq/AQdK9BXvsIHGX3UViKCg0i2ASFzPMbUKTFg
t3gVlazD7CqvnzWM217whCmA7fa089tzG3QUiM2d2vnWSQARBRu5MV18CkoiIFypWSlIZ0MR1aS1
QjYJ8qjlVrRj9ka/+MjZp32VL5D0Y1TMPE6fFgG+/pwkn0tB6QymXy7hKQSofMNbuRZfLPOrm8y9
szYutQ0ON5Xg6OyYs0ionBehdYVZq1lZBdsNVlCa4w5EfUe1BRJoVYaXwYLRbTY8tCJoCewItByt
7xSqtkr+npUhsHTOwEhd7pxEqgh9eHLTln4hqg6rSdt1x6qQIZrmugJhzH6Y16x2rHEmp1nlkESv
/dMSpIXC5pDUfXazakZ8sHRUSf2gA2qsf7F8sqy6RXxPVMV+rCwSdSoR6JUI8FSkPMcO0gQMeAYZ
Gs1nS4/SQv4iRNj/yZuGGU77lCEPzSQsCjLdHWrwliI3K5OQBZy5GJhhlB/J00AT5JMJHxOpK7Ir
F3pIAcDlc7tWXI/blvpRr85JcV7IgxqL4qwStGuNZA6vpXVVrPACKovqVMCVxmxoTa906J9Bc+j2
EnLh/WA7ZfFIRfvodnYVzF0UAAo988zxHmLZmb4y2FSL5i0EivltgT60OVt/ST61QR8CiDQlD4+k
zbMss5GeabC67DoHJJ5arSabiBLRj4Ted9Lhqd7rgmwpy1RBHpsCW3tZdtixoKdWBEuYkNZeC0eP
H/1t5kPL+sgeXmXj5K4wm5cwexNZQvD2+U+FCimtxMsrfkZgaVg1tEEH0v7mrWKcRZ3Rilu33yzI
N1D8SG67UNs2E9b24JO6cAs+x/XwoZRaNFdOwYVIuo3fZl5YZif88pLUhyTdFuM7rUGFntvYd7O8
+K3G0XcAVFLaaQUMt2osOXqdp1k4MwakVPzzwOGdIvNe2mmJ7aoXa81iinzGdKiKhXLmPHS+uXr1
Vf9o8o7l4aqihWtcs2po/lMRIZG0pNz0RCJHeBV3VVmz0ZHXt95cDiHyrESp2+jX/chR9Nby9cBf
nxWuHD3kDCWrk0JyuAnWh9NiYFjNXNf1wKQaF+hzyMZoik7ehzdMrDdtgxH+GPK1cpPaXzuBQe5i
AXZBU8OBHV5lYyG1x/fOxyQuQgI6so3CcRmGwNVbRJBW1dvLwZzt/aGutX5syMlA5+5OKyB5x3Qc
o1l617tEZn5yH8fFOx8KMK/DgPxz3bFsa5e52Cpf8P1A9hCfL7oTMaLYa9wk63FcLqCsC0krluqK
UBj/w6QSLzRDeX9iudfQtCvc29TtYKhdpETo50494GDiBs+1iOkBLFlMaV0HA71qXAwHUpdyEd95
5gSqXdKq+aIMi7MhDHFZuJnzRdoSE/WDkWhN4SXcluHF1ik/fZ9PQLWpQUhJLT3bbyf0VT1mXGiF
IlAe5aZd+NWxoaqzYNpj1+3312vdF55g6Xkk9jfN+oAVx5Pje3DWWeq0zSk8CG6oXSkUcjgCLphA
YZB6HnTYwywr7sN78m4AzCYjAjhoKNqV01w5h+eirCDGOvfnrN85XvrZphLM5phaFFFuR2pMEzsy
tRH8cUAIKGJTwp/gdcOTkmaO6kyOND0g3SDSqq8/79EORxeeA4LOmsD3NUXynMnXfQaWFVrZw+KO
xdiZx1XgzKdROCRh5RhTkl0bdWzuPRsSTotxWjLmqNoBYlS9fXbcXNaQx/kDzpAQmX84327ycLNh
fUmV8f/BkwatVkrOoGfp85Lo7Ni9xFv0aVmB9BdGQtU9DQJEQ6Z1N0S+wPFnggAu6ja1WP65MCle
QKuktARAvCCeBN6Y2sbtCuojLyO6tMILo7QQ7Fki3QHxXeEBUXGEyXJieKbcUr7I6877lNVc5964
f7y0mzHmFbK2KF7BYkXrrrSrrCY+61GcpIwTjqfUedxlq6pCK0HM80YftNC00NmchjeGXnr3imo6
fsU8dex7Y3oiZFb8ifI5O6szVm5jq7UI8FKBSu7l9E0Arv8qriPBTqnHlA26W9OLGhHRCLc453ZH
IaYQZsfpvHkPa+JJKWvcQZ3aW4jsoGchuGG3C1OqwNbaiJ5nTSj5GxIe8YN9uNfhi82yt7hw4A8K
4CuGHn4qgh4pVjY/EwVQGz+LJ8xt6J5BJh3RB2tDMiUY9COvIpvcCAi0iGCnT9VJpaJQxKFU1ivm
L1HD7kHbpvGFqP/3Wzk450AciIVKyd4e0nNRaVEsCmXhxln4PPIb8H7ItV0GgdRMOnjYxXUuxaXn
VzzadoiDScAOMuYlxoB3bS1mCC98tMR1AnbnzMMdAkMhwlqZ8TLm1aM9Efh9+YorDc230zwR/qSC
UBXb7wszW55C9veft+5nJxXyv9R9vbyZLBVkdkNdNMpUNIxS61u9ctaE01WtzSO8Lblyh5VJsItx
z+18Xqroan9uDkd+G9Ohs6JU0raW5dWnmjd5lBpenG0s6HRUYq82QqzQPhw5OKP5p2UjczXVhCba
/pw8/j2j3mTTOfLpFZm9l8Yiy5Nkmrjz2x1qU+YUmK9lEcaxLQojTC3zVn6j6WthMXGcgnrTxvKb
u3aZv0IqgG4g1kyyWH5aBxikyZI+zOIQlzha+OxJXIjvm7dsakcs8CzAiqdMSTthVZ72kB++tTRJ
cyVV/7TS0+YiU+BFqO9N0V8aecA5tQ3Hc94iJmLt5PI+JtgzWVYBW8Fl3MqhtVuXY59Gc9dHiRao
OPX2p8n5H+niYrPnjww8MYPWMw/5dIQe0LgW5NwujEszEy2HdwXdX7Kenpcy0t/i6VLN3J16hdlg
mAd3DfxJgmjCrzYSybU5rGBH198llaw8uQ78FP/JhNK2oVCMLKpcrnLIipi0MnOpSvLIc89WxHay
ej/HqP7kwWfH17Uo0XNZenCeHqzzHw42tX6KPKHSoproalR+pGE1iCtdvAQe7G04CT64AR9BW4oB
pISN/9QLKBKi/f10/t6c67roUtET5kSEpHmlVaTzbizTmLs09WVz7C9lWsWoUI1/60ZTEKV2Cd/4
6vOsO9HcYm8uNTXHl3JnGlkLWCZ7LvyyFG6PCbkFphMt1vmEOjpDYBwB+h8eX/ykZCP/GbbdPJts
Tnk3jYdVVQMMBMfOkQ0kbGAk8dsq2omlZx18GEDOpD13iDVM6fZ/0DF36QtWdPI4vX2g7VybJpIH
DR0YKarWKl7UmEX/IzKnwzl1RgRAybkB02jEGmzkpR2rYB7VrY9ghqK50DcXdLJzhMqsWgiB0Vvc
pWz/E9QJUjyMlpneBBvD33xHCL9FID+dm9q+GXaGAZD92TVSn74DQp01rhbFgzsONsWfrHCPxNXc
rbpjGUuzGvs9RgBZOiTYOCDN7bvqlK8nfuc8jQ6wkF0Aurzmcm15XGEf9fU41m/BnwdJQ1j+Tjz5
uxLcOv0TpNH8ZWXsc/gwI39Z5b12x2cKBW4bSvHy0mcgTqCZhf9WW7+X+Mi8W1D6cdKPedNVFrlb
BsSPerPMGDm9xXgWlQoy37vh3wmwSA8HIDYJ5MG8ofHm7ssu2atn4KWW9ejTihtnq17OxtLgnHcf
HuMzkOfj7Rs7grjSp7pzJyyChuyTKanQBGYqHZ4LO/KHkQq71QISEPAMFXn6fB9ogX2FzNUaimRA
mDAtsOOI7TbNjCJAFUJlpYWiIzbUpY1xHB3EnsmktIshDhJLF+xtrWXMbFa8oQKytgkNcoydfg0Z
fGDA0jxmqtzegTCPrOC0T6PfIw3lmFMHaw7g9yAM9Nl9TM8sHNlMRi7jV7dfc4kZkxpa/ECjcfFF
jtkfzPUNKa/E/v5LpwuN6lt/saV4oqVqZc2xrxhMTTM2wmCl5PSn2hgWZe2/D3zBoDnbuUFLsGn/
2Vzoo/QlnarT62P/dXkJIKPv2nXFkuMSyBm+StmdIiJYhqdSHY8OLg9u3mLY3EsIwpu1awNBTqYj
Xdpj+MWP89cUp6tnIlaktq+1txOpKB/4nkofZea9Gm3CMJT8NZVrvQv7n/7Z+3nn2sf5DVv8K+F+
GiYRDac7MS9yLvSkQFYQgcq9NOdjUABG5+BEOiQfLvwG9juYQt54ocdP7rVb/LJRMwOI3Sdz6jxw
KIa2rBiP1E+93cJiAmkdsZ9HVu9sT778caRuy+GPX3amyIBj3b+TMxXPLBNrUTrthhqTWgBiJ2Wc
F2RhJY8CE41ZM4oCtf5QU/PAEwyc2vRUkIsKlo5Z9JlnaoShnqf/lk9OZVTR03+W8Gs87uXy2wXu
OJmZrWm8T49vaWhK/TLSQ9CyFyT/AvYQgj6J5UcqzYgkMMfOejFJvyD26+6HvuDYucxSBT2Xn1Cn
r8VY2H5pnl/hwlJ/iQ2jeYne8fORD8qdj0TVW6bNNfK9z2FpA15qpTV0PZTX9IlDsUzFZZ2oC/YB
A4ws9+X/bi8zutC6BvQdz0zZ9j+iiDLpOCxwQeHNZLlI8mibXRFo6u4DTLAtXIDsxVNbP3mnquwq
E5YwbNKkAmscRADPCoam+KBLSnYSAjSSjyA8WGQqxtDGp05tk2BzsEEY7tUPwiR9pK/Mji7H+YBH
rgxM377hICX+ISvCSh73UglF2Sc2PG/0aMK5wa2ui9qp8oSIkqAcu6NAKDnVY6OF5RIru7MICcW9
GQ18KpsLX6sFE52yz58IhIC03XED100on9GYwXjKYmtaxBsnPyVqI5Lqn/OGCxAbznjGoLpPlZX+
HObDMh6CzDXVahCyk8Qv+se4osZPSGqcKM1GoMNnCwll2j09HeVYHh8DgiUs8JNCoEu1XTOy0SqE
MS4UpfD4qBETTnOtxJTRHuqfDjdXtuUyEeKYAkxYti0P8zi8e959NNeHQ3w2IErVDKlYnobVO2ha
F93R4A2yKidyPMjELKMEnNpvJaRRKsejWHIv4h9+T4eRYy+sb/dgNqek7r/VCVTSmU+/T/FouMjd
8FyFlAJw+NmukVHTnfXIdWd8F+p8UgmfbeLFomnO1/to0DPeLPNinAql62SPYzKcdeT87MzWywIj
aZ87uIWYoJ2tvXBo1V7qMUcajgXDgL5k4uO9ofqnIWmd0PMfNupemvFjEnucHq9SvMDlG7ofx+AZ
MUmQOPJcycuWzbdEtU+P0osqvM3ubJzgE9NBZaKyMhiaCJvtEHj+lbgYN7tDq7FoovG1Ku920gC7
4tsN4cXFyugTBNBrz2GhwyuHM7mq2cJM9Bsmf7OVjiOG//pV+gSjcX5+sE8VBHhor+iDOnb9xPO4
0YeeF9GjcxG6f1Ri6qDNxeMvDSFSrmOyaGdaGX0rVt75xNMHOkCPmX/RFZBGLmrkZ37rGKwLiZA0
MvgWY97TK0mbHklQQYgru3aNl9kS9TcnxPE/d47N2Rort46GMuCpT3BAah71Lmd4anJ3EHqQ8IB7
LkBhDvOHo3v+mXSb0wenZBnw0SyXJyLpBhp5kdbetZ8DGrpjA6mbMccpdkw+TBKfE8aMKOc5rPcC
hnhVtpweqzcZZpamChaFs2Rha9r9sHcH2dx25k0L95+HovTC+5uZNg/vbUG6zrf2C/6PDtGyh6Z/
HuHcrNvPZJD7JkkCo8uYo7MyyP1GniLQDodvyYOKLG66A6dQ+60nPnERF/6TT3jyYb4vkBmJg6A9
t8HWSuS+lXzVAgx5gA7gnb25XUBkgwZUEQrWKgm0P6j1r1jCe8IcQSrGssV1jlVhNtHpjPpqbwD3
zPPz3/ft/H/pcq3dC7X6KyOZRSMUUTZ9tAq3nlrPJX+VMiLjsVjc7mIsEiH0NsmVQBlEg/blZlJd
JUGv50SZyBohyRNpfSMtkO7Gr1a/EBmrkKE7zQx+Xeg48mukHF0eToTtnVLrknJMy8tmQKSyns+V
oH1oOSfYGuv+mCkINrL2WOcpS5RoR9xgLdugQLB7OvPWnVAU/5G4H5QUvWjJ6dpDey8fikG3CNjF
iQlc2pSM08lp7Zgps/gdjWoEJ0yaVEJ/+UPTQ2MWimHxgX39+U6oNJok26RBKBQRVCU+0M/SNCOd
/X5nJ9ovKhbqpA7fmOiXO5nNVm6J3ulRTryHFysT7OSi33VNu9myYULFO8vXcvCp56chf7ZQOh28
tyOtAMoNagfka0odYdI/UmiyrEmpxh6TBHGb2bnf1SOJCvvJ2C+l+DKa0oRhP8O6btp9egpeEAd8
C/opE79Wyctvpj3+YQYqzgykFPDXCk3yDIqi5b8hbO2Z/T5oShgvuylL0kwGt2S6De9OzAzYG06+
Ly5pAYp4qor635il3QjU8/vDG/Qu3pjOA3KFPmz268ilUGmhxZi9CjXaDSSq1D9t0WmWrS8gHnqm
zLYFX3pKv2rjf/IYG5Fh/oa6Q8qg+/8uLNvrJtAoYa+iEYTcQFboermVpbs14NPQxW14iF3zI/b7
GihRDYqCHs0XKqbVwnSKpDISDGuYLw+wUx69pDNM4Dgls4YVGyr9MMWp7RgkNr7yqyql518r8VL3
aj/ln5FyEGV78j4ZF65gKF6iJBB267CUEagYclRo2G+M/46zKufOzPpN232L26Uayf6VNtQiYyXw
p5JMxxggWQjWMQhUNKsg9XPd+7SZSvnJqhADYJJ8kCEBHtplMQFLToSJqK6O5pyKKguQyF0owhcm
dmfqdNBm+FXTltls1Npk8Fm145wDdNqg0E4YVcCIbd2CRs2sURfV9J0WN8Vb6m0M8kKsukMcsPgF
dCP/s0tmginkbn8JViaQzUpBmb0lirstuF0Sj05RhxkZNsatytqmsmN79Lpf+S4iWuqp0LSNQzLu
TBrofwevsn0dEJG2g1OyG5zOH+xnAlMVSQOXoCRPTI7KdT5G11mLjNAu3LxICBjcj+VU1jhkYFS0
p4AS65wweoLEZGqHlXM88ewvjWlRmhyWdPQXCJyqjuTEyeEeBa5KIfgBRUyBFjzh0FNN/rcq5vpX
pYtSr/bg+KOC4fB6Ur/pq6CwbXuJw+AdayICOC9TEMmaoROw1V0dYEa/DS/cX2PMzk5DJ8sQpzS1
s4DjYm4o9F1ALEu/xefq3KqglyozLxui8O3rghlqFek5mBi9xLxxtmskUUZUMXTG+N+hBUeagnp/
IsATpJUe4zz/PjA74gHnHXpN89vG2I6JWBuhXi6PchpwJ/s9QhP/7B9/Ww8QZMghAelAL4Ky4zqL
xo2+vubm9ggSAjj0050DgRd3IG/983Onm5j75qpG8IJH0S2jn77Pmcjl2v4qkNIOhzZZ04t3rr2G
AM8ltAFWBWea8Z0fsuSWbF+iYJsihXZA3ICY5PbfpyseAmmTgJ8zD+t+hG9QoME/B6jhqHgI0Ge9
i8qO5XDqsrextm1aLCTJgjRq7ketxbCAinQsuEEEBZS7X6uR5sGeN+FKlgYiHR0Sq00H9yZWV8sj
9Wdn5JpSys6kxHS0Oekz32P3f/AyyoXGU+Zx+fynaKXl6LIN2RXIZPAAPNRXlIjN1SuBi8AW5am+
lbmc4usjncbGxM+z3ISX8EVol6FJNZlY6twlvTT4ICvdvh72nbQVI29Ze3bRt+0JWLCEGR6fglBi
ga9dM4Yw5WuyM79H4RDEUQdOaDe+H9UkfEMcbAOVCegXMGvNhiW+RpCji8kEVR5norQKHURNTVLv
f2J9LUL7pKUB3DufJvGmMi/ejh8MMBjENTFmTR0gbe5XzEBLB+UWmJzrxznC95Gwm3W26rFzENCe
WxV3eDxNjm3DEAyw2doQE7+wyokX/SxORbwZjr+i4fRl2n0f5A2obs5gCAMMpd+wD57Z1MDhujtu
iI8qB2AmeYZf8DSpDlFgB0nI2xnGXhGZPjzFlbFMf3r5BuLvUELDH3MUFR0O0wqcwf3/X0lEu/ve
dTxa3E7tdfxGD6sSXSp10ut9yt238KLoDFmcG9vUaxhwV5wX2C3XBKqp8t+tEskqeJO9umFW4USN
tdx5zhTJGCn7f/TDV0XaPAdqGSKkNG6uZjbN4idqpmYlZ0f1E86EfFcjFo1tS450zbInsn2EPsQT
DbOOTTEqQM3CtSY/IwgUSuGZfE1z8+H549QtKVo3bumSuiGis8ztpoZwT0lKiCfJ9oYrmmnZ+Mpy
7vs9puklHQq2M/+xdAXpFHhhfSxPo4aIVRfPh/PF+2rqwE54b0FXXFWHMc5geZ8wodltZKoUwV2O
5VKQWxytnQNWfPy6z3oS+ASL2d+MtiCWHTCJOQtzvWj/62aYE33a7Y61NRpRr8RIhR4dD8wLkiFP
hIlgHUOaszYzzGwIbAwaMoyVxYp8WqRV4syn0uX3/MAkjWLG+chSrh3Tt8cawxtROIv6OCwLmrom
JUM9+KOZCjIY8JefpulYv5GZZXdbee9jF50iH9QApCSgICSPzIubjK2W3N3inrvF8uT3GIk+B7nf
S2elaaBVey2t89DnixNebUZbGVxW6dK7DbzznvQdvtXUcVC5cAnDIJDzBdxuyk6Hkd65l5v/E5fR
CqqnGwBCpZYkVc6nwteJP0WSkHFVGDn8u6/ugMjhPNOaj+X6mWwZhlUWcawTPi7Y2Sm7UAp7Odxn
X+WPbhfoaaqX28aCT4hgje43g/D/eQfVPByAVxgwx6LxhuZ+BpZDWvSM/MTo0CjWUDwd9TIgw3Zj
PnuPlnymj4ArNAMI0D4TfFfAOCVkzxJmPDJHAUxTfHszti3mlbsBwmKMRMbGcl+ckAj2yYsK/ZLA
lzuvykDxKYg4HAK8jdH3mAKuuVCo7xZVSAs5JJKXchCIbinx1ECn34iRwmjyHjImDrkOmS+hrKZg
ImP3qWiCYqt7wOBo+WQgxbzpcOzrpd/BuODXXixl/ApGY8k5g00TL0COAoNLyABYiX+x1q/MGwAr
kdc41Pr8+L1LUeZOfAD11peQcA3HKzUah2x+tEjUOdMeULfVImlQYPZMY2jIGxfmhsYfo4FC8oUy
JgnkfT2GYd2k3foWeehZfVlznqpfn577/0FWTm8EraCy1ee1P7/rNHHLneZACH7e/BUbeQZ3rpFn
oaTDmRelZHRYeobPQVnvPRsj3/o3s90hIwNS0IgPysImtqPnkL4PwUQ97cmF/dqSc3hUK6/cUQh2
L36XwSivoKfGeNnRxUDuerQzEeCXq1kqPl8kC3g7q1aJgAeEMXbELXKPR2kjjF8g2LKU3fqOp42a
8/6LclIUu2S7vAtZOO7X+kLBHuahWlOHUHj4mDmBimVhPx/Fq7L2aSod4RvF+P3CPN92/0l/pRnZ
FFnsTq97vPciJthT/m4oJ1QzAv7M0UZKS/QoUU+u1ULCdrwJeMohBwvX0kAq3eiC6avJoMCmDy6X
We3eaD+NkQYGTyIQHgIyRga2f8MixNkqRiFd9CwEFCenDIgf8uHzZNobI/CUlmeZ04NZDpR4ySes
pfgEDP/YpldWg8hqLyVbV96JJMTwd0Jb2tvjRaBx6Q5wrg0ZB+q/1ev7QtyegMUvisfDIXkLYft4
HoPJg54wFvZ5B9yHE0DykpOWe1o3SxVOl3vOwGQVCEtild+/aIFS/YkwiJIYkNIb7lbr58/4ZhLz
cN/t9gC7GGfnxcR609EMcEbYEaDaMNMrv5rZ1MJcyWv80FAvGBjlqmoFEhmn+uYpByAx558Dnepb
sGIBTSz4YZP9gtEVDfkzXgpzOcx9cQG3AOqf4Sq8ECowTqXdOpKdCZbW5syzBcc6uRXJl7hpkrH7
5xWZ9jAgKrT+5yJnVTiJIlbbRhdKlSCv1VTKowACcZrWo2yaGY2A27jx4IDAX6JAOqV2lJ4aaCR+
6z150iWCnMy1z4HHq2d2Rp8QZKAgpxzDnXTAaznxYUByrRfRPq7e/UwrzL2teOsjgbGoLh3Aw1M6
x6PVcDs0CkfeYhryj5krQj2DptgLki9oDJ4GBPgcWSDJ9htluTGHwVW07mdGNSTqrn9e9tIxkmRg
2n4IAEHOGqnybeq67XpWgQhkZe1OQA2BPm2r477L5iV7Sz8Ye69L8AyfFOPmdBhydFjENwPRiPD4
8I4gTQVTFTKyKnPP2rMXw1y5cAvoK04Ts20XEvqx/lcGnUmYQ6YbHuGpK4KnfqjA6fGqaCbRNbHu
FoqJsMDdYuYIwuHlJmfsQt/riJTd5jhnxNEf24qfkNZSTcfVpzBE2mGrwooMjVno1OECy0UiYads
VeECUVk6FzGF4YWDLZC4SdWHGYVsgE7S9FyijaefRYWlr+Z/kTe/N5PgXPkwNbnL6tSDpWPgZBlI
DWaXJ+0T6bxX3QVYCq2sB0vD9PhaeC/bmifu8W9PI5cbUudVWAH9ZG9pdb+EyqexIWNfoj9LVruw
MrpZKbALPusoaVGuJy+y6ozuEKMjKSQrVpkh1YRSn+/5FYEjpgAqtfTFAJsS77BlPVrY7SBq+Y3k
Yy6SrbXiC9+dWaQ2J5iyBrCs0KFgUxQsoYcWu8oshVTy60PANiK9ckf2M6Hs/fzEZfnblXm2SoAd
v+v+SVEPbAFI/Ww0obeLWkPiYtCoTpKE4c8ZxTG6iZGqNb7mzKEKIaRfgSCtTDHtT4adfDe/lECm
R9HBGWvlzCSn17cwnrtZmj4ZO7rt0WiMVSVnRJ4LkkPmzZlERAdzmpGCjZmsVylEeqs4gr1U79gC
hVmDGiNeYaqq7wnZ3fkhkU92RgFXfcUioE84ueKtPK4sfhXSWM7x/O8d0dWMLCfK9IToyyB/x9FA
+b0a9rXdve8uF0w6o/hwboZdsCjLxptfh0I/AfsEraW8XZpkd25Ec25JFI6zSfwR6g0lMe8eVnSC
BAzqrqCVrxI8zYKlOcx5RGpC6kJ55QM3ouXi8aG/NCMN00H0q6mNmfpkCKkoV0v3P1+utEmBVeo/
Q+7IWa3lGWlhFog84J558Cx9qO3yr2YazRCmj5j1fwGvBFC7dP6JksDbbhV66YIlUiHETZokYd54
YhUhJu6rlJa4juRu6e9MPgpLrdA0sVGPGaKAdSiXcaKWUvbtGd/sB3+akfln4UJKDW7WBl5VxOtP
HnDf20XRV/hgSl1rCF1wl4FB5VA/FU2anR+zq4wIzbyIqJnzKSCzFAEGgHM7rmsWcoSCTJaHr6Cw
sy6dI1UI5ciWj+dfvc2d0EEeM5Rjc8PUGl6R05O1VKP93NOCLeGssqopp1UrekBoT2S6AlM1uOhx
wS5tSYUTbhjXisxDRdqLuvK+Yketw+F9s/aC5c7Vbu/PZQaP4er3viwLqdu6a6rjh/wdz02sGax+
p89LOquJAY5NnZlQZRIYN46w0rTjmLdljC3j9MM2m8SRP6DI8thnIOu1mDoha9D6iVHUe2W1p/yC
bAcDukE/EsTkA//GZCFR7qNF73kdUOAXXZN4j8c63tYAS0Q8e0FG3ZSURhyQ4/4n6b9XMm+GJCDr
ZXuqYGoIH5vCJTJpvAkc5xwnzrOrG+0zz43iGj12O36H6iIh9XtuTlaU2OUMm4ZqcbB9D+uY8G3t
HUMM9Y8TbYn1G/5wMMTWSDNDOC6+YRLUsFJ/tLXfAlt5vJ0cwPoanSs+4f54Y6ZZwJC93udhA+/S
RpaOYCgFXesTbJ7kZeMlwvFLRaJvmDfVa4ob4VPoelgRiShCiOBuk21UcHvh8yhphFr1XfO/WS3/
Reqpf2QBY6v3wB8g3UnjEHGfy6APZf/9ERscrr2srO06vWLcIKlZgHN4HtiH0N3VNH/llIpDlVrs
ENfGMyOSOP2sp5GwY8FVj4mNij+JscsORYEhBYGG/8Fta6LvnGNgBw6UDXTuUTyiUzvtIM8lKvAZ
PIqTfYtouuHuYWyggIXZIEPYGtqBZZfuOxRu5wbhCvvEIGYHQMMPVmOZDWLQXkYlbyU5hozw+SD5
3tiAtmJ64yXH4NPJYNV9Wy7bWhFdocHD8Qx/UuivIBsIL5i9hG4xpFXVkZYRkZFx41U7uLHt2LAP
zNfKqwe3JeJ8fd1v0kwwRnNDg8KwVuaFNQ6btdezAfXn8rodhs9R5JGWRa7bL3F6Im93YqXfqMQ5
LjEx1tI2YqKd1kgVtRfu4p/heE05fCCn9TiUzQin9PohTQOzaWsuVf6/bOI6hAwad5tf2XoWBkg1
8SFJyhW081Ipa+zeSVdCnf6HESIf9qnJK/wsv+D7twU3O/r+jrVtfen4oHMFbOjBY7iB+ffodJFD
aSzeuXrEk6WAYBOrjC4wYXpXEAaz3whUjijgDatSm3zSDLcO098OBWmPoE2UBqTV6igjCpIqOMKS
T6nM1PqIRJdX2a3WSCUPYp4csQ5M0N7b52UJ7p8RvTZwUtAaIH5aaaXQDGm55c5Op95Ld0gQwkVJ
A5rh+jEfUXCxwmYEaVRvusgtB3nL2HkH/64otbE90xJE0I/POv8r3EtsWNrQJhoSGDKXxk9/+0Ut
ixu897//ijmLbNV+ap6WQzru8Yy30IF087N10FEOJRwXuhndx5ZgfiJTxuEJ2+20OnzEFo8v+65B
6vhLcQiZZGLibGdVFBhPSKW2SWbQ/NwtG6Df92hP53FukzmPRU7cjBy5hntsAE4ijoX3n1QbgShy
lv5joUwbsqlqdB7mGxIes/mTb9xOgP2LjirGnGgQWXPgorolFezB7Der3iZvxc1vozP9+SDZ1qy8
8JzUmefX2xFpFuqYW5qlbLcfuWqph3D7guh2cJ3aq1zBmi79i66xC/FLKFn094Y+1X2IV7Ze6kYC
/Hru8nV3xeRO1L0WwLdkrLgSWDMdvZr7Ja/pYBR/dtJdhkvuMmRrx6ncRNTMSA7/VXJEWVsvv1yF
ImlGd9bts2XYyY5idwTepuxVN3i/PQiJ1nTUAn2Os/9VFrwu3+v2kYv6Ye3DkiY0Q4Zmh7RFB20Q
/1WfprlXIgTc3DkKUT+M8deM3kJQXMbKarzDWR5zl5ZMY/Vb9ia1vpzFyE3jEOMnWQaV54FzRGoc
iSDGQb03yr40XRrxEu1g2StQHtwg4P464M96i+luorvIQQF04Pv5Jyuh5N4suc/fdq0+M3ODOnzL
Vp9oXmqvXwCOjoec1DEsJ5RKkR1wgzBqKkAq+eNsRBA38o2auSlNsowxqbR2DZExAwPMgAi24tzD
FeDu5tHXcGYQxsUKO+hTGxleNEctZeqri3rQFBhqx4XscqOvMg+NSZYcw98NSEsGUvGu/9DdwBq8
TwRficItQqry03sRi+ShKZUzLVxBNHdhg/SFykbuIS0BhnjPOuN5hCicQgIbDvXQdff4gfX5cdWw
E5A7sWnka1Rom0bTiwkpxuCwJpUPdpmYmps3P+rCUBimaC662owk08rSzjwMkpCBJKPzOjBVQgJb
UljRHu49sBLOxdwkME7N16MCja7ED3UmByQJxO4+9VqdnQcLvF+TH4QPWU/M1SsZKhC+jMb7TRcA
ALUbY+jegDMkkEw7tPEtyeNeHPmhZHRXM32Liay4ajd7I3KbLJsoOqF6miTHTZ8f1m4q2Ebgda09
mNTUO+k7I5gSvnL5j0YZ4HEcb47BpOFT43h6n4XeTw/UK77aIpKy8Tf9nFXrGNJ6mFQ3trU8dJfR
mBBf9zMfY5N/Wt3xUiemGTjRSU/35sqx5Vzf4FR4WvXRpyu2WvdFruYLEN4V9Re6eYQBRkvgmqr+
eONVpQ/+7b6yt1ADutA69SOk8PR1xmX60Jgf64dmvBYE2Zu1W42EYzI2qxjIx0XtPe8FHRjbEtfF
DY0WSc69PzyCQ2xOyjBe+0Jn0y5vUL0fXjyL/3hNy1qsApSojf+C2pEJzdj2x17De4GYPJSluV8l
2Pb/cSJ9LsyV1odh62ztD9iB1bIgNSzC/cc2cyzUvNnt009Uiir8ZwpbeD8FtEirCp2hne1jhuME
hI3aFTwrCrhstqlnfXTAgyRnQN6mEu2vPWYYr+3WOzAyHzjIe1LG5TloEFN4bb2+Bq3kh05HtjjX
E6jZ2IndDw1a/K56hk61sFHuevAbOV0lGK+/UifMaNPHElCa1B2MGfKgEliL0/RRN5b5l2TEqVwt
+gtDhYW3rOSP9gEkQ3lAec0h2pJ3LOfJXavKYPDFOwFt7gc0UGWrkblgNNB2ak+TjOIzLgcwHl4U
l51kANX3fkTiVbrZbHfqx57ZwMGH7R4WJYqs7jleuAfZCG/i2mC9csqe8XRTqbchmWx4EFpZuuLt
UDSqu87pyCx0TmS2OJdADFiHN8xLda1LAfxhgBRfH8IG+2aYZCVMA11eH+FBjF/xIMGXTYx7G8vw
X9++lYUPtSGL/f/pZ1okRsnhiNHOnyNxIIwwjoriUmfNBspGvxNjTbN260myySQdLaOWp4sspTnK
cELpxOc0dGe1rMsGHL09uybPriz3pCHmgxZ9w3xNgeg4KN4IpxHv172F5x++b0zqbhl7rupyKGRS
jKU3AbLK5az2gcgRdm1m2EDkW7NbDXRTsVgGP5Khy9u0hvJf6c55FpnPxa3NpVtTILEGxy+58w04
WdrPSizmxsPkupWwyvUfy+cj3ZPfUY+HMfOUjKuu/OPG+roJ+DhGebkiZyEXTmi4yv7oEq9uyJTJ
3u8qFoEHxI3qHZ/teQvr+8jBSQ9p801N4lwMN96jA3icXWhhcM9kTNRjTbKGQqoYH9+07A4NNsqw
GmURhyxFSxJywlm8OUrZe+uTSOjnbogfLlM1l8POeEBn2ou5KsR+5Oi7koBJFISMkIIB2pvyUVi2
+iR3S5M8BOXC+m2+aG5mIGa93kNHq+4hvGxVdIBLysDYgu4bAXIxle4m8EM6zlyIAxqZbwuLu/5h
FDnOtCruf3bqNA/ztQZedTuqlD2kxvtvcxYFnkArL/0TV7tCy2ZKp3fNlgnQ7clBKVDl3lFROcOZ
NxfTmUaNHD4XOkoxMAKYO3x/ePBM1JInMu7P47sy6F3HTYKyEoVUq/JGWJoMSWzNaz4e1YYpfoac
FupPJh1v3IaL1MXZiwIpCnzZbQbiFcOavEsh5MmKLhOOoGkwtSo5k21S9b5r1Arqjfsbmih3UusL
Xjk8jRBaVFd1uVDfh6ebMgeSnQRTraQWWrn733uAEjnkURewCDxJFgK4g7r66RfH8Vz3F153nBuH
BP8ZUqBGP8zGO2KIo3hzqVikwPeazaZm16eo+KfEXHQkniRw+SqrXYaaLtJTjdADnSw0KwBCC99X
ssZA1VQGDdWgzqGGzOFFzMLrUTunu4rR0XI2irWhQU9hG+PuxHWFxZdZSNUP22GkDEY9sgXXJ+ru
e7t6PolPR43uq3UldCN/xcqz4jImKdqenuqFro9+5s/8c2+OSHriwWMpZ/vp4hWxH5UcnwNAXgBo
44l7UjPLn9Fv6U/nol8BJsYOWT0TIvs0AR1tY/51c8lDtqJzvA6YtFr8fDJEwrlhFnQuewC+Ci+J
UVkdOXtah7N7DPNiqg8qRSd35Hmn8WT+qEdfPoz+ni0AUVg67yGJCz/q6+RDnmLUX4pSQ+mldFs7
snTDi+k896AOxoL8/F5jfYp3eyjWsXZyt+1n5voUGLsCeo3wpsT9zQm3JqAZlmH8VHCG/GfMvdnY
s1B+WljQcIsMYFvczSoiENqOw/ao4D5t7dub+1lDW+9Z5GtvKgcb1zGx0hC1VrRzLrZTBP6fmt+T
01kK/JpOFmozOnOAhh3179Re+PRUsl2+5OWn4gQca6a39SPTeYDBOkYbS90XOEfRsvirImUjUy8H
6xViMezHrlKFFsiOEEBLSMpknhqhulplgJUo375/dhAbkQpmmchr/mjbhJQUJL8zhuSD243KAIQm
Tyf9iGa+4FiWIQTk1Wjl4i2k0llUnb9FApH8+OmftmKTDZgpIy9yh9go+FuQBOEJ9IliHGFdBcvD
boCj+obLW4FpBWEXirjur/LcnGcIfDP3fPnhLBg/ZmTmujwQpORBq2s6OPeKRTuEf+/bp8Wv6U5I
uaIWKoVNTfY4RfZVcKlMOCEHYdcHhqMKa8yMKiY8Onvk/RPWrHp5m929MRpDI1tQlkay8lJLItmP
BOJKlBeHtj6EdhBD70WHeZAL9z0iEfnWTeo/VlDyZfVTt4GRRUczZgd7UuyTNYSj5I/VTiGKxzam
RSOY4uG2tBVlgeaW0YHq9MoC5uIQ+4Oxt/rsc+34+X/m86Q0XLLO7HcoSYi16ckegjIio8cpfEuJ
q5BqcC3Xj3iQVUNbIH/xOiasW/iJSqOTYaUFoOLhrAaFAeg31OyhlfCdci8NpTXdAfZJskDqUDuU
Bs0thgdEd4+r4mkV1Ij+d6bnNv+3kF8wNXYr2NJW8xUs/vO3YdOO6llztK9QSV9nsOsao6z/+97x
4QH+Ra0Nq1Q4PVk+DLRvhwEUBkiYnEA7RaguSFXntEJHtDlGhebMLgNHLkUjx92xN+tjdmm2dBB3
a4RWXDT7yyzHzVWPuMR+3JdO5+xp0wE2m9TqBBLHly8ySpypXWzpZaT7o/WNl5YOGvuXtHNq8kYf
PCfRgIHd2R7l/2ll35D6tN88NqQqaYsUzNTYHFahnnJ33N5immRLR+tJe5q0La79/F1SdX/Vo3cI
0wRoYaGWVH/TzYp42j9xXt3KiXxgXesGRdi7ebmG9csffSJg2sMM3pYmd/TDkPw5o0pGpti4xWiJ
XmuGNFiUm6ZxbVgRKivKgvEa/lrQxcVW0F7TsQAAjrPjGE2D9vvU1kJjohMm7JuuoDA1FfCb05vl
Iw/JuB6rCIzhg9gahvGJAH6/0qoeqD5r6/BbomYlbrrcO5I1Gt0u5M5jOWdGFsjoG7m77KbB6+ky
pn1lL7l+fk2WmaVIM3R8Ub1lvLhTjtbwAPPam54J5l1wxGmlzSkSY4KOhwIvP9Pl8YEe1KwUjnrZ
Z+4iY8J98rADhDoPxnS6jDBp7v9eTbA8CUoIFGDrjt+6E1DfLLTBcAJXOJ8l7m8yGgmG97MXJ0Qa
yGM9+DJJxlYlPpbvvhbHgkwOlPB5NAgmKAa0Q+GcljTowfnvy3R5O7UTy1WiRsoy2n77409lsjNR
sEhEsUjr89bxMC3V8Lh+9H70HoFae9TtQVk25ZQXA8JRX9Oiba1kXT5PvXPheO3+abNl+AZKu8fW
HYa30l3WWBcbIQxyskQlzzr8ToqO/z5k3HNWNjisdobjtn/TdTeUxJj2IVavTYiZdhbwouNystAO
qtFPyyjwif3ib/bUTKGH+7tjBLmtTbW/m2Uqwt5jFXjRUdoAeyVNR20v+rpj2pvqdFGVIVL3vxIp
Q7OTkFn0lpoQIWq8I5ASET7H1GRnfAkOjQdcRKKFWihHUfSeRX3z1ENzqek9TYI6GUXE2MHaZ5GI
lUBB6CLpEYT9+yMhgRbbF52KKhL66pc4Pfm8J93RiEGVOiBwcdDLGB9f3lqDU1tqSeBu3IPR0KWk
yZ+A+tkTwUWOkYtzTGWAAEMFuXFM2iqSI4GXac4/40FM9dOVeXIHgHKv8y0L3mJ7G3xeO5m8V0+B
a8NNllTBM5EHvbuS7/AHU84Ho4+wT5fQuo9yf5ivkGPLrWfYk4GdHx2pOYwbo3OKe7USvOWGsb3o
ZtbpPnJ0y7qVcl4XVgL02ZAjLrkbGe+EfCI2IMtz5iEP42LK1XWbT/xlz1alXYUBP84rwMXYuC8G
eUSCStvXTRM+h9umV97ISx0oBiG1EKsnuYNQkK9P6HoXL2+ZAFiUc5rmmNz3PanQMw6S8MRcdxpB
/reL/AtvYe5m9eUa8a4lF0ARgKPXUZgMg6B1IVrLvW3CXVuZLHqUMeR216LzIr3lWHxTlscIRDx8
SYNYqzr3XOhD3zvveHkvWEeyJS11NrkG3dnvHn3xV1H77wm+JZg3NNvlCqCKFMcyaFuTrKC0usKd
tCbDBZLNDkeD4WJXrgsWTBIoU4hU9CeqOd2/mY2T4IUsm8Mr0rMWTViAN/JfwsQuY2Dsy1d+V37S
sz6Y7D4KCLOaxX104I/EEvkqNhOAkqarHgQhB1EjMaeFORM2LcDIhCaYxRHK/R0NcyS9+CgBzDW6
1GnuPpt9DRa+4YijGX2UckuUKT1Po33PWTDCc2fw2haGRHxJe3TvLrela0botFlOlPI2bmCuMnrV
QUZzMFkCTAWPsQYXR28pmDBzauMaNAV+suRdbRmlIOKpWJsnDjesEsTVKR6OGDrDEfLG09y7waHh
DRS/9KxAmb0NszflueqdQB8E+fZ8NYpceRaK2dwJXgDhrX6wBO2Pai/Djvnd1k9k1yE9nm5iqGvV
f8tjTR4wmfPwvusNhptsTc8I3AR3rrAUAGDcag76llcb1Ta5Yg10ccQLQuwGP0pibe8/Jn6evH2i
KBDOBJrM+xdNy2s8hsvruKBOVP7RexJS96VCe17p+yP8OKiecElHlHe2IOyuuEI2aBJjQG+aKH5S
KmPI0owJg7oSn7Spufe51M5yXdW3OL4CZ5lKVRjkZJmK8j7lX73zms2vcSlw78ocXmIfSr9f7yIp
wrizBLXhkah7q6SMCjyaP/O9C0lVgMr5d/DPikpfD/nAER9JtzjlmQC65hA8IjfY5J+Y40CiGUEk
ttAlbva++/B8FggDX++1WzN8K1PKZpRKbOl/kFQgsOS+XEJtD8KnlNfnPhh0STz4PTXYpIPDFCno
amCqrRU56AQhp/bCyEQQs3kwp/ksCyQUTjVcUs7W4TrzVhHN4wdciWVuZO5Vnvd5p24KHBYOuHHl
v7WdZwUx2Wb6KBpJUsdaPzD9I5GpGLJCm/4KFstNiC+OcmpIeGKKDcpIwT5PoafqXBp3cYQ2bgE4
SptzSHHFPBrO9jTYHxiTSq/Bm/0CuhcRjfkMjaH4GRzeiKeJwFdkve1VdeuHZ/px8cU5BRCD6Enh
XW5ivG2SAjkgm1n1j9fpc7wuPdOHyfpI8xGe96VFrE+9yJ3+ihRTFSdmVbIk/OT66GrxqwZZqK96
GutZCiFEVOiqnBPT+ULQ0+WqKmz5xQf+4tApYO++tb4kS29ZYztd5hFqhTbFWT4QPSD6WteC+54j
smTirZlaR3MdtG2PH7epiP9KqpVWKonyXm7IOK0zS7r1zrga7sJWVjhVbEPDSBaiOH7j+9nJowS/
Obpbl7NlX2xXRlRrs9cM4zhpAVhutE44gwv+LHEbP5wce75mLWly8PkBBlhTTlpz/vstFY9bpGXl
pKHJECa5tiE7ALNJEEVqKnNuMMjuTvhWbKW3zOpL534Iyw4//G+vUQT12zGVdfUq7gjWR05O6cKY
FohguibZPPFzWr8oMj1St3QjV66FJ5Secx/KBVrkEMi7rzMVO/ZH1lLvVRXMIcJ6ZlNcGtPgBkxQ
SHcSd3Sk87p9LioCWTnmXPqb5j3cjIlJfFe75FfuBU+eR7aipUL6Fpa/q/qi2X/hY2KMMlivz5JT
mbqf0I8GL9jdPogqwWYKcNdwqPz5eIPqPh/oJUtbaP5j+Yx9UnTW17rPaJJR+JPikxkg7vBMCsTF
u8nwLy4AoOy8pqro5n1YO0IJoCBr5yDnpDTn0fCgN5yZxw+T9TMTmris/KpOBZjHiQ3CAqL/7iml
64rq/0v6G7Agrx63a31wTpN6SsxVMY1VlsXG1M+OVikYOBs5e8M7ic61fBl/GKmHHA7sHbFA5+zT
P2NA/RRrLtG8mPIi4htf2ScDO04YKvXam0kSfzsry3oj0RuCNOU1O7YxiR1TzdgnfmkJsziYWRFk
JZu23UpZvq35Txl5psi3B7nUbI7Qrb4agkj80JgQ45/h/0XvFAtCA/6+NoLOK3xzZXvVnufcLN4L
iFvfVKlLdxqyqANJBbjD3JGGNZ2MbZul2Ehe2UKhRAAYv8lcLS96YS6JoGcPyeqaVuaB30qGGh0+
GXt4jCK7ai5I+VjRUHMxjgBbV4htTAWmCSWxoD8M1IxBMRVNGj8zKTS9G35eKumIjrMIsGKN1cpt
l9h18Hloc0zYOmwDHoiv9Qnx4kxX/L4X1bT7rWsxj8XdfWuAVT88Nv4eHNyXHjmmCFqn2goWIin5
VI1DZC8/oLzxP/xBLKEArvUq7xHXybYDOphdGUpvcGspiNHA1c5a1ebzJqmktRTP0LH71mj3KxfK
/9UxYthxinPtu/yj4IONe5TJOlufzR/RzE+Ysjt3mD1DgirPg+0JJuym6ot2hngCmOeo2L+qzTBL
cjerdX8N4LC+mASDKBusIERjgZTMipT9RlXPyAnNHO9r7Sf/HAfYe9efsb7an1jv8BqJmX8Nyqs6
IQgC+eWevlFu5+loEYhzPd3lLzEqk3wH8CTiyFhXBfM0pnFj5YWH9rAD39eqY+0laTu9a4tb/zZQ
2DQBhAy7KBDs91AVIkUURhO57mhjEf6AwL1Uad/QQUGfm/Wc0zGIPO1lPl/2Er2hQVfnSk0xYQOs
SrM4ciFfnGpqBQVhp8tU9PkFfEsBKvVciM9hBp7IqXgCp1p7H0ELgROdhSqX40YijZM77NNjcckS
bX6jKBU0oqYnzSplVuaLwjHz4P47z17DqJPIOD4BmYuPc/DH6pO20gk9xn4C4PBUi1S+SN35sp1P
gdxpmt/zygEzmHaA33iuVmQF2tTrjnNEr7u9GVsAnaYjLFGs5CrbqHzli1ewfqpY2v1/y98jzO5U
KjKh6U866GHja5zRFP7TuMcpYFoQXnHJuXCQ3VxU4WYy//EEG+S2JjOwjhcgpmm9M823sEjmmdoe
o8S0ymY71pGVCWlwzVX8eHL62jb4921caZDGulTGRAsks2Hpvyk10B8ey4MSWDC4P2NHxWqiuBxJ
vO/GxmoJYBffzfINtbAqip/yHWd4S5dsZ3bB2lzX8t48K5v164F0xJL5ii1XYyKP1oI2s9c94+Y+
vL39W4orCY6bmN3HgGXcCW22mRB1Ec8MR59SK2OSIyhy4YoXwdY7+fqmA8T1GrXwsEJSv66cmiqc
yu78TItNftMsrNOcymssW5OjIKSf6Du/5Y+kNdgMqMzvVxd+w7FIZ5EbnOgzzrdbB8N+8Tex6kjH
s8SzNVEh+5ln5nQEZirNm2T7XvxLXKHUhgPuHXHBGKa+8VyYm5LTiTKGHO9jKo2MKTkf8lUmL0sN
tT+5aRPp9+mJPqMNQ34i328MVMPr/O4N/IlATDQTQX3WkX7OsfEgW5arB+5+LS+LY24V5LXaLE7J
Oj9hbiGEgpOz93DUklF63PmnhPJ0hgcKFcOM/MQlaWmbrsCBm0fB7ieAl1wFOc6PKCoBU+BXVkVc
bjlPySpdePn5ztxAzlAkXIeF5SZnIgUxnrzUN9tvPOXeS/TgltH7+/2/EoBd6BSVQeoPKsYRO8Tf
ooJOIXgtZRdlz2JWBaG4cqfK/sLWMF3i604aFlFE0jPx+Cnh7YSbKaaWncaYUvRwz9MI/qmVwjFY
d6EVwwwWdZ3ySI0hpr4a4cG+uJRzSX1LpuNk5c95JcJFgKTr0tuMF4MTNPiIS3wcnWiJ5TV1C3Zb
8+k8e5N6vobVLA7daqJBgbk8Q0eSCJ3Xf5rYgVnoMx/c7MXCtbXCTKwFU0g1z+fI8O0D25bKMgKM
FBZFlDNYzpK5Bkjtk0bnfTBQS6IMmmBCRhHoVKY8M3spZHZ4U7Y7xVwwd8aQlryjxRq6N1LzL/ku
vS/8+rhaH3yxs8p62f7ZApD0BXwMO0sQeOKYuEkoUQPyOQ7WgkMry5woGkBJgdiS3fX0ozDL30kP
2c25sFYoUL1Nthie2H2mN8lbCRKdPjPpOtwX7SzdJTUQHcwpmLir4/Wfer10M7Bu/K2bgvPM+sn/
bYKPQHcXtFjOzNms7CJPhTRF53RDgE4CG3SXnjv7LI0nO0PjN+9ssSGM5i/FZNL36DmxyQxHKX+H
LmFNp5+ODS2hNTEPRGEpFOFPkwrk6rnEuhMPsuz7I0vVIhcgML1BpetDrW5mAGGpXcaVCMbOAZor
4fjFNGhxjHGflguj72DdC0W9htiklmAXLm0A27YRBeTixRlWrTZgF3rregpFGbBi7cJL32KM+n+9
Pz48D486elWhZqa1jNnEGpdidBYe/e7ztNAmNSnjP4p/X03OHHnop9YhB83BOaCqVFO3QGiCC2L0
BDpF7HUgD6uV/IwndbWMPAa0YxXFhCHWS2NLJ2gnMii4FnafOq21++URWDctC4yqEpEH0hsVg0W6
nqWePb6XoZEBtoHgDUcPkx9S4bs4juKp+0epyHDs3MwboawD5+R/KMO7HLMxg0aN4euS7FEC9u93
0Yobp1uf3vVa99FmJZIOOZ/rR68QWLUuAGRD+hmCr5O+bGlVvQcei3z9Lixj3hTSbzXvFYjlGM/l
3VQCKG7yfy97a4ZRQkCgg7M6VxXO29NI8Ue/E69A4PClvTzOuLp8K1VQohyahF/HwH1VJfCByvc0
NvVzNYbrYCSisPIXWzt1O0sAKuR6Kj6ak3FONJ6ojgrl5+C4w7YtW7K565jFlZ81rmBNrKx7UNQg
HmMkYDJ67FeZUgYOfluu0M1sK8UhON7EyNb798Jx+TjBT8JUsjlYQHr2ZoTKu1EDIXJ+4fxMbdK8
O4kDcgOEZKhcd63J7BH1iMamaR4BbD14yEEppMHc/bFH1ysNWiCKQozGWj7/AJw3tPcsfmcV1TDn
keVdOM2RWhF3tV3pmiFHksipgFGdvpX6BrcJOEJGvdaty5wonaDplV5NG5XE5tLQ+VjiU+BGYF/c
dIlhFNtVG+yKa5sVTpv+Ydun+AMwjbt9LegC6KY6VVZGvBnU0zzla03c4jeLzLjezQmsaVoCyuCO
PDXp33o/z1c/xnIN8Fl90XLOa/T5ItdNUgg6At9RDOTPj+fXEY6llcD4pq6ThO2FwOxNY48uRQof
L4OabYgN3wv8sbW6au3SxyLFYr9fRW5yBv5XGraSrAUzsgX2fwSIb3TqxIjFkCL9vzDSJOYIdMgO
92q6xdSAYeUuqNytLrp0ct2Wzx+I9R2c07d9wNAQY5Amvh9/qi7E+NoAFxPxO6aCVH4yG1p/bu5T
LG9L7A9pq+Q/Qd+babWJt5TawAVe59QDXxfxaYCxWEmJNiL4jYHtb6+tUxJJ/+FNlgdX11tPzzxJ
8kDnIFYVgqG+0M76Lk3vt/xVJ9D028YLM9OyBF0k61Qfqj1CpHAdZJPDIwIAfKtynayFAJCytRMK
cDTUmpUXUDPblseTDagRvLmS4bx4wwZYDsMoefeJcwzE4EkCYqew+mORXI3qv2GNG4a0cX4oPdH0
u4ycZXlLHxrcjQiQyATWIb+GRzs026hQgKVtAEXvxFAvvz/oHkeEkHJRN6hni4p0wk3bMm3qkLrK
yUNNG5dCXZVgix6Ab6Bc0O9MMULIcybc1797EEwpkI+OTsRJ88zsbLp/LrWVRPq67OFVTlxGpDpy
6Gh/cAGCV5MTMALNc6cT/uHyQ+81tNbRgguyvv+/z1dCz7yuihvofY4pfRGNfT1z1T6vBJ6SnuFD
HaEpY79svqprVYwgBhVDV0zTmRa4TrgHTfSrs+Ntw1IAXfbGrLo6r0o3+uFL6Jg4pucNd4ZSYLHW
froh7KgQIecx4yEWzCtIAuQYzwl5url9tvNE9MlPCTSId+n0Hk6WfK4Ba/PSzfEZVXGFLMxeHSoL
mU+oHi8+JgP5KJ3INCxSyyJUqgfBVkCV6mfCElVv6M5898T014TNzliXmToQ3Hue8e3VJKR9rclt
ciwUfRLeC1lIV+0/xfOJxL1poqqY2VGMmsGeFiB7r2MQNcepy3qcAFM5+5fGIi2mefeYlxkwrYWd
jv+p+Oid2fAlSts4gQJOdF5SxysuL1gstvlOLeBIGz41hQ1LqMdj+j3SHS3+eC6YtxldovoMrSSG
VUOsv6wQPxN3qdbM5i4JpVkDbmGpptePnvNVMUH1lbAv95YDicik2QPT5jKCMVvbJwIN2j7Rrtwy
QwnqAvB9JyYrjOTL53XJ3EfxnfTbx6xM7ivw9pa8BTcAwY3qsy/VmRAIQO09z0t15H6qyivWE1ZO
SWUwywKQBf5ruYeFFS4X20nJvSYpwq7EJA2thZ5euD82qDpjkRTN3SF4uDLBklWUiwzE1eKYnB9w
WCvi7I4sO5rL5+Qq2OcX8CNVbs+aoBdxGe6qCw9wUH53pqhWsNCaouQajJUkhNAgm2kw3XtaKFPD
UKu0n9jdMkoLTpE7JmWkdowp07UnbF19o4mmkunjXt0mmXcsJVPwt6uquzyPTq4mfxkbGi9DHxKZ
oOV23PCHPI9iAwzvx2IwX7q8kdtDJsHXYBBXlc5vjEVk6MjSFDRAIxim37v7M53B2w55/RBGSK20
VNzcjDYyZE0Sq47/oLiJMepP2Sg2JWwUwVzSHMk6qxlQnO/fyHzFw2JlX/mNx78tKUyWZkK621Mb
kugYt09WpHWJNojkGK5cQYD8tMN4slsVzn8GOHEDLP90JffBo4wPF4o0pm8szMOPmQdvKZyiaX8k
EtZjhWpKIK5STg3l+hDQbXJYLBJbIceAwcF3dJ91B35FcnaxDmp2G+vhS+7PrVpthiCTctb0t2/G
IQnKiaAclYB6mQZGpXOtzI/mw46GX7narFCbkNytul3bc+nPMYknyWN4sW6/6douGfK9HLBdSyAp
2Rgic9inEmnCSKgDLa1GpyGmXwTQtM0sWTgsDVhQ06Yc5hzCZlOVTttRTT3qKRJbI+XFY3o52F8D
f5Kl7wDKyVINunJUP0g8rbDpJJkTAPMslOHMYogKKqX2XFYReEpJZQXUDi+mrFMdbuw/NmRzBwuP
F+VEgrgOAplrudU7E79nbAEiw3B8opXIkjvitTmkpOBy2YgjFmoVkd5Ez/MicPsRVqwco+aYT3jl
pEFxx9DvyQTT9jkdjXXRwLwen5b8syueKfOorhAQiOKXS8EO7U5bPI7Wj7YRrAnv5i78ZTXUnZgz
gTUQ4JNmBITkN2mvZNI6qL36x24MvnfMQ8afUUVh2u4ZwvMxW/7nc0YmqUkLy+bI1AAVbZEgp4G/
peSCfv4tVCkOBH70taUATjv9u4zCOpfuyr16DS8ESNSjAZlwJFANcmDCTCi0xtKMCOo0qa2LpBjW
uslqWEstrnHZviocRKNPz/0XUUs0iobSt5P0eLWt5QlwsZsewkgqs/AI61sGLHMnnSNnQSK3Z5oz
RvOQJmV1zr+s07kZfiH+w+xw5BHpgjd9M8IdR+GA9NQNbSmkypBj11KtdDoFQkrc0igV+5du4+DP
S+k4YLBOvoOKJSF27H7jOh/OFTGGKtU+5jifbKF3jz78IlkebwMiASTNtx3psO9fc5Zd7OcYdmCf
wHajIqFkRuB0E/4NGb9zf1axpYwyJAr0pGSfIVCUPY2/lpV2f5UP5UCsoP0j1HZ/adOvoMF3TWIc
zR/rBv4DHc4B6S99lHNF2y6mTk7QcB46M6TU1mRm2fuhipVmf+0XGwNLwK/iovuzBMw2SeITPMTh
PfywmS5RjKLD9vfEGdhiHO7mK/Ty39MBlX7B4DvUmEHWRPupBSIR6DqLszz4yxvFyAd523IUodI7
rpMCJqshcnhe3DAKOI+SzwyCsIakxrzBh7je7vcoYaqrDCu9/L6f/xhwGvSSDpufhCaCfGqq1uYj
eCTQPwCUHNFBVMVsLNa2eo0v50htnPQvpqpn17vROE0kpZD44u8WnZCuSVZZ25GqhVXi4X1whHvr
9NAfOElnLz1zdDZGaU7apS6F5ETB1BqNpeF6Nnc+m+xKMjvhYUKEUyXoUwTfLIFJRbvOz4UqM3dB
gRcCXZTjf/CJyMH7HglgyTQLLEB/Y7wgAnMCcwJDD0S5rA86E1Z8LUj1jJsuS0Wdbp2I8W+daJcA
BBBjq9T5PPNPlsZfmpJ4xZdlv83zLFBUq+zxB80mzcwNEBzmcTxCkubqNov/pEPytfXX4AJFg00i
Z41UyRDMHRQVZF7Kp3DK+4nvV0VqT7yhRhaIix5ulwllyM+b3JK43Iur1xYpkxUNb4PAuBkiEQTV
/FuH/k4cZyKkfcq1QbCTo3Hy8hNGcGNe2fAauZZ/zLFikDKkdVWrlPaSOugdGSpfsQ3G4EK6GWep
9x7o0QREQjdaQTm+4+sPZ8QdRzOUBp5T1q57MEsAm3KViWbNwq2JapTMgk/P4BJzPzA+W33D0QFh
3BMtliZjhRR/5fzYfDZo1/dxbjn1cEGlFlYavm/3hJqv8qaz/Fv1VipCqeG7EQ+X3tbOvYZ93maV
rELeMvi8thuTEy32kEXKpwC3/LE8LlAqVCgfrfp0OobcU7F7svoIYZ1zbP3ITJ5hMWQINKQw8XdD
05bRQMES3avKD6hW85xJg2vgvhNFRYINDxVZFWybbKoBcgqw2g5nq3RC/ZSctk75gqCtRvgzUins
ADcNfUfURSO02YZmCTcMFP03beWhGX6KYNyk9gzkgcv95Av6bKLSrGeaNv5XGaofYcpzJt+UNzmx
ax+gTbcuPhraqNKIiuY1oFwRNGNIGRDmh/xzfKmhQh+wxsJoZumjUTsn+KhanTVMzQ748AJ9lhkk
ekWAm3CyeR03sItXKcsMcr0oyrmBcTq0ji4CCt7JFrHWwaPWww9BqNprbR26GfeTIcHUFMolcjKB
sLibjhbXzguXH49MIpOvQ1SElsa2SqKTlN0Nb7h9DrgwBZG9c5hrXsH1mHJNy2xGHHc4wtoPTJNz
v6JOST4yhfguIGJgODd1Kbf4U7fJN6elSxUWCXIRzdJ38D/LTs86NfDWuDNDwA+bYWk+LW5FaDv4
cuaHI4wY46SCPspN7cylrg0aZOsGKHvKM+y/0rKcuuWpZqoAUJADvkYRjocHY1KVe6588ZXU0Dz4
jhb5lntXuO4wWR5hnoFuU0wkKacVx/xrH5plRlq8U7LId4yNM1IYzNzEGUXizt1nXXbvlXUpm3jf
Cs9T96cwfr22fmCdWhv90UYY4VnUZ0B9cjozr+nZxXmsYSuDi0XP9x2Kl2vuXhZIRa6SrLaAzLFh
uD2hQyx4wBuvsjByf1kg1XCcrDxJO1gsyJ6gyt7XjZjbhOq3EY6b5CqkO4rJtUQyt9XmpCXbS7mG
bjsyRJ6EVYeBYO9mpY+bEDk5ixwID4dHzh0UxExl+XSUlQ3v77ikHGTsAJADSmKpRXs7vAyZNbnh
SB3J1/VIaIXBXk0T6mXQuOxQDFqCASURuPGQV2vTEPZK3a6jeGP3sq5CPV/UKC15uIm0RxzgStSk
pAsdbmlPVVMf48S06k0wcSkqKyXtfL57HhKCh+wIi6GroUt4dt/0XFTBy8D0UvqWVFvtCZfS4oCg
TfEhViH8NCfQkzWMQuBrYTe2EYwjzzgrtcY1TrbECinBICzsvQiT6Qd0c3gJGNAy6ccNgc7YOBdu
tRMhU0XcABxEFQXCmDt6fNJC1N04rAZhk54xznWV99s9yvIbvnF9LpL+BAnz6rmhCy12YFPi7Dnh
D1FmBx2rTAdKzPuheFnLl5C15jGFTLeJDvvErMeYNo3WWvysdeQn5NaQWQ65K/VzbZo7Ls6vDxat
IDwFsIAARSxNn2hvxJIf+YXD+ZnR/cMinj5vaCE3v0zzFDmF4Gyre33LZspaEEt8NBWJZfxprXHt
ADkX/tHcB5qdpmYQ+GQSOq1tEGL6ipxYr65V2HkhnDw7PvCl9pyYGhJ6qKIj/P/btU4wmrLpCfup
/k2vo+JF6XIq+zBLzBVPVQSbSt3yuf1Bp/y7+12Yw4M3MxRFnvpfexHdnGMi7B+OXeEOKddDAzMw
Q1arhf73LYIsAgzOVsUzFOqjxoWIys79900pfkcRmu/yvlO8G5F/HfZwB/2zREBtYe6t+4d/cTmt
SOeKnr++ytXV7ZCbXNZeArZ1b0qBZXLfRheamD+1Tq9PmGiE4RBU1Wj+YDTgR5MSKcR5n/e1KAp/
OobQx/mVjRQSD8yRJ7nFk5slc+9RuEsVMQrO2P3+i6sm/c9GhAXyg1418BzN7hGRVS9c1I3DRDEL
Z4UPoWaviEMps8vVL/5xItrTHhYW+eQQu0b8SUiewde/nFfqPwaTV5OlB9UFrC/dK2eDMP0Pln51
ADpc3PFWBLIUcwg0oEXr/3GsLK9BuOTIQzCzgbP98ZgNR4euPCA9mP5vnw8nLcgLKRiN3035Uuez
8crimLQOUPINugr1e0Pbc9eEJtMOoYSg4Z3PCAEsHRMfC3TL1WUUzovK2Rc7NC9AxCBEFsZwYH1L
V8dF52eRSlBpGN2ZZNS0gRNVV9fmNivtF46f0kYoxWb4R1/1Cy3elUDLeU/N+AbinLrrhat9+b0Y
piK+KoJ9sHry/3DcOFMccWIzruJHYOjjl0TYqzkSJxZAtsELTgltNXj3EPS7duOmUqxzyP5mDMWA
G43F9Q9BgMwVuRuiQMM/pvbw1JLekeBxt3V5dmiMXwipAbpxJ1GL0yroZig4hOCpVT2y15HFFaUm
oWOhEsvxYBQWA/x0zJTcxQOOzVLRvvTUsZhWRfDheWY+XHy1NDEJUep6t9aZh2C+GirAzAHMaqJ4
Jn9iAbit53+e2i8mC+238ESgWJ8PI7Yug4b/H+kIoindA0WiLdY23kIiPViRy5wEYiZQeQzdqt+r
tMnVzQUaarTUEuHK/tHsT54pkK0C20daG8/WadqdI8utrfW84BnIdijogL7V1XPCUpDVCb9cqUzy
f7vZVR92xaRivQbVWhWHS0SJSKkI8v7jkSIn/Y3C1vx/jFip1tBj1A4iGLFAAO6C4gXWcNFhWErq
NwqdDKpL2adlwcdeQNNG3r6AIVtm0byGNHSCH5clbcN8BeEzRQ6rJqfghPh2A3p/GyYhyecVcATA
BWvgUWgR4VP3T4ExBDy9xJ7GuhtGNXE2bL4cCR7CUtyVWikI319dX0xUQM+Ft1lp0CkZtS1ogHfR
392aA9FsSAS2/E6UMvNpo90lhWZUG8KjdGi5SsFoCL2EwCcOPQDR2f5vbJS93syuXzqgmpIdQWCz
5+aMfZgCzdzom5QtxUbf3PCbyd06b2lLOxqVn1UUYFDumgUMJ1529SuLmuIMbhNB5vNDNPHflp7v
icZkCoQYL3FNx7DUPSvdvlir3vgFrhc5qm747gbHc4I5moCcwuKR9O1F5qWxlFREXYtJK+0zzNK1
13ddD5Ao+MHJWRz3FmhT7PNS+wVxglpO+f5pbJENyjqJ1Np639VQXdABsze+dwMwLHmyPHD8Qu9h
AhUYgJcjrqzPmr4IvRr3hUeLOS4ktOtmbDEGN0CK9P/Co2SZbG4psy00sNVq2LPjE/iBEwDYqe65
+8KtjBpBs5+9pXSKezQyzp6/qykt0UPSrZMnmlebw+AuIDfsvu6b2OwDljwRqO1Q/IwM1wyH9OVY
uB8ivkCv2cOz1KBLDhrE3Mw+slCjbQliqHebYIQAv7qNs+1n8tTTGIm45i16Y6ICYxJ7a7qlR4xl
71Wx53oS8Rgsb4kZE6fV3CACSoQKslTqYshQGD4VhqBj32v0yynzA5y7q5onSLCLLfF0MDNVRnzD
zUkxmOPPhZLr4Wvd5MbhNqtfFI9ISvUJArXtY+VgQnm5fEVSnAxVDIKyvvF1X87/4oDaVnHJCTeE
3eMFhciyy0P30e8arlxLSeyuDouwJY6zHQ8IM9txRiKtvKl+EElBzrLNKNTzLXCZcpclvKCk4SYZ
2NiIA6YLP4XuJxTWq+vJBYNuN7bccHpTumKjJmKBm7/ChZopqKhvy1MBng8/UnmqQDS7nzJcvbru
h4EunSj4NKxT7UutvyFgY6uRorvCho9qvyTYWDFTmjld3xBvJca7dOBzvnbZpJlam/3iB1LnqshT
ZwLLn4yUoKFDRnoODCRdG6xm26XagZGOBDrFuIMhn11+Je3lPc/OJZVbhWZBlnQqptEKlcjy8ohI
siWGFK5JELIbm1P/3VfTEtZAlTJ4XRNZPw/QpOWeuBheL8XNtGBJAQjznPkuzQoKI/aik5ZwFeyG
Sa7AkIEMG4gfGsFVWwvoHB5kFTZkd59izEFVW/SlesBrMr/U3QTg4mmqtVpIfmbwPGNFJkUMQ6nz
0/80xziOfrrxm1xB4v3jI12obcggUFbo/B/P2wlsZfXMzO938n3xUPWZEQG8fy7R+0/T61go/EPb
vAkLgKguCrhMbXUzmh8TFnMqJQe9EGvPHOlrbjSRm7k2SnyAPdxfvUutOz4U9R1vFyoMchh8ox6o
pce5aTDiMDokXbc3SyGpQyQFsUVj0YPqf6+Ab6EXakST7J3vo9oc788jTm5sNQw7t15TpfuXjpHR
fRdVMLdMLtWapvsElxxKSN3zJQlRBbj7T+6fOrAtPyDiEZd+8b2V6ZgVWlrFwEk9c5/7Id5JqLHk
t2lOVvg3Oos+3ugHPuBJeZpAoC0JU/P70LyVAbnoeLmnhcYEJQyPxQdYF1XgCQ7EptYBKtEpTpRO
AHJ/43DUrt/UJkbbwO8Hbagz7IPsIm/DFb6UKBGOKVR58tQ0rH8GtBCj/klPzc0x/Z7HcdtGmQAl
yUSOdwttJBEpCIU0R+c7jpEavWuu/KrkCfqKbBxWeh9h4a32Fa+WyTMf65RKOIw9icv02VrxgeeL
3tsxbQu8iVmrc7y/DQyq7oy9oUk9BMT6vACDfU8yazuUJwwdVE0GBNn9YoE9FtiHHyUCLkH9SVSF
6ETsHrm/aVPdDzuNFTWr5kOnxcDravPu/AjndOgQ/Zjusn7nlqgCWV7s6dQ602wJ3rQlxqOdP+oS
Le08tVOVawnEm/hX4voeIHlql8M5rRN13woe16/9aGkn0ZZ9B/q2IMC1kqeLN9x5oMecMXTL01XV
9U715e2utPy8j+TNHl60MtAzysA2MojF8JLh/aqcvu18LsAe8SNekgA2AimUGOkxiXbpWPDVTdYc
HT7Ej14dEC79bcPYbQEzVPCiFsBuZxjEqo4JPXx9etLPSfaChn0G4aPFEXtVXxvdwBYhxYbmG+TH
9ndXv7tuNuSszTehZOYmNzLLCBEEEJqVc0yRbN6R6mmWhkGY+SSQd9mz7jxUpxXe1+yRcmroUZd0
u+fn+EHxNeMz5mehsFpNOUYPYG3wGXD0DVoDkWt4ldSK/Sc2MViKwy9SIeGXkdkexo/lEEjeZf0N
RMMABU6Q0z8xEr88VZS2wO+ShfuSrEKw6KRW6UasyxrAV5Du8elp/wst8T/2/xb24U2hdgE4I67q
v5RXCltLfaIrXZfxudx5N3o2Ce7QpJXqX51yaMjBB6F9vcn4eMZ1/2dNIMG7UiYlHsIh56N4/jbh
JzkPeD2hga5xC50gatQCnqMaqhzEBJQ/nCATIT8zDL58GjTlvOdMhR9Am8gUA/hIWuE4/FQDd/nK
NpujG495cwaWOZj0EzlKMfx818/PC7LxVNRy5JulnMWW8sLerX3wpYYI6TwXebI1Gq9JagGtABkH
s/NYIjTZCBmDWJPHDghMFir4Xlivvq9TH0TfQAUOLPCrBV2uk6rukKHyHvL2F1JvhiOztryBnLCW
HL1GkR4Pe5Ugj3yp2hyZR5zZyJXAly1nBkPVYjbMYkulBlJlNb5R7V3pAn4JmmysBWx1vk8ZEugA
D9FAyfshJuTH9tnNbdXW6Xo0xir/Xx1YyjKlopcmzJ1bHAnB4EsO+A5jyjqEmSad8lJygVsz5IQx
tDhgIWBiLaMzm1m8/fTOSmz4twaSaiUUaOijocLbGu5B6V8k1uVueUENbKyf4/uqg+3+NMbzdaFu
fqbR9Pym+AwR85OcaNjWrkGqEzIJ7IZtTl6GDr76MRideByN6h7QPgPT66hb/f0DgVGz4GfgEW7L
6npn0uvHTqDGTWtW2cnPZIxvPHLImA5Hz3n5NgxvCnYjr+rU2Mkgq0m1ZpnCSM7vSfcvVasl+8vR
qQOBx7nOxcw3n4stfA+AK725wmvSdtGncFSgU3TJS9nD9fzroWGDEhsPRjD8mnv97UD9CBzUjQcK
EvoMkazFiuz0xNrno5WVQc7dwbzyDqyhz4q+/Dl5jlOtAeutnjPSldqVet8sdevufH0GAMf7rvI1
AbvqzNxgM4BAxkyDSylM/W3gXmcqHiudtqs55wnF1lesnhh08WnIr+oQYxDNOiNlA8rGzQ0p057K
64eOtNlk5ZgvA/1RX+gKslsP3yHvwCL5gHYgEn6eCx61TAdFlItuQg6icj0wsVBDid5s2+vRry0U
ecvgoJjzwO5Aw9EQOz+8w1O5Zy/LDFnq/YZ/833tRszge1a/nHsJx0vXme14+Mt/T8Qp04bKHXf3
6iLjejTnQtmlezfh3VRgfBqp6LFZBz3sxSBrLToYGg07NvmDUA3j72dG/eL5xBABCuVfqhzKADQh
QPVde4cc9EWMtItwYEvAppVlUITZ67ctUBQGsdAbSfNHSMVXvaUBg9pQBfLH3qKZfnBR02JS+B2H
npdrXro9679rrY7NXAseru178qAMsPtXjpExPiL++l06kc007u/hFJGhflBuLP7rRdbnJ3ELHx1U
Q5of7qdkFxNuxV+TrksmDws+AjA7bgFDMeze+1gzQxwxuZ67qSNgfJqSIHMWRcJmuph3Fe10A/2t
CqBHqf0Y2zBh+Z2YU0beyEyz91LNuEd0cZyi+aXrOMsZHdZszmVNG91M+xG2TxAwaPVrV7MlJoWM
/3VfsnRaRQ/rfIc1WCM7k5OAgg1KOdc6jpsPkovaLUOgWlh93rIa/BYCvO1g0PKOulM9yLfcOnHk
vVk8ClDHSnRHGRKumHiPxKSuM9IocpLjB7qvwUYC68Y6+aKgrbDMxtDfZsaESoXdrJZbtv11SsCj
SfCbof+S0/DEGmSJf8LWF17DvCw3N/ltde9KlZLSl3NLPhrtvJ1lhMrpbfH4m45KpXDtnegD8c3D
8IKvQB+BhtphZJF0Z5e51WkL1cf9kUMaLqkkSkIQatcR5aLFt86evK/MDHySeowo4CkThrvSWf4I
GCCn/LeUmYDrcK7IODNOAb/gtxIq+YBBcGheQ/ob3XjmcYPIr3U77XozbVVX9VVjpCw6EshP5Uzm
Th/aUDj6n/PlXCMQqd1SmLPpCVXORMajqSikH8ZefFQLS2t1OvRLigF67K5Kf/WGiy8UTvOVPCSc
Cj/dgXjcKwEdcHJKzZPjBM4xE+ay7U8nOmwfumHZw/5ikaU+hPs1xwfnly5d2THEuYQt65WCae+c
D3UqfD6H4UH+pF3WegJeFwoIFh+a7jlqJGA4PHYPRiVM9WtJskAwkbV1mUz7S7QW9BdyUSSVjrSm
IGRNg7ycZLitJvsA+i+1WNA+iUQMq6R0c0J5Uv//Awd1zwfC/exvDdfGOTUiOByQnt2errZ10l8A
DD0pfWWlVnD+5oK6NF/R68kf0xZ2ADb5jT/lg7xBHBFcVjbzA1qWGkOUPYvfbP9AwwOdBJ9js66E
5yPE4m5OqLEj1eS8B+vh6/Cz/GKfkN7kCzANiFBMCfvK2NHZrt+eoMyDPvjLpJUeB44rXkJ4lcAK
g1IPLjsbWZ1iY/Iq0cJplcyXHhISPLQdsdOK5lcua4SO+MmI8mJHajh9PUOnotQ2f2kHLaYynvde
dsRBYWRtQ56SBqaL/NUlZDpYI8ypYdYEF0QbgDFwhef/PUVU9H25ql/2/3q/MmZ1ExXU6mFEE0CS
Nd+fc9H0D/J8LjVQS/xdYkPahjsmTkK45ncGHWgB7Biz05U1rqb3mFncebYGJIpTvOXghzdjw3uS
MognEV1cgyQLjsfeohTirkMA0Pa5PMhDbTwap6RtuRKYCnxuk80byVXE0OkIemwTPBHWxYtVrfqZ
0SnzlsQjkQhKnpgDmmptXpMutS3Y4AW67z8667zwY1KzGVCk3KIGTA2J/erE/Vh14TzYVLF8f/Wt
EFCwL5rgJbvd7j1q6TwmglO2wYNgkiNxmkVEg77NvgH/0+sLgkhGxeYaJwKeZgWpuNPc1zRgDFGp
HtrTM76qIDKSjSCxoaFE8NtCC+SRc+W189rg82eKNrDnUrDRHj2ap5wQx9b2ctj8MI7ayYJpn9Ur
ijS8YXUMiuVk30XcKAZX5JR4yh0ffx5/GWpdKgvr7X1Yr69JGZTakHarLdAzj5riP5V1VGHfrJEr
jTGpE7eltj/TKVi5MoBg7a31UGAzzcowFh7jKXwQ8XwF95VmIhlOhplY7icz7Dr6HN7jaYqN27cb
CsZ6VZ5hdHvmiC9zJ5FUELNpbSWawuJ26f7cvvKFurvpg77A4LB/GQJwkacE4h9sIPmQMQozWFl+
nW+iJObRUtpjmBq5373GAllNqERvQk8y+Nr3UJ2rwMfS/U5VhqwC/3C8vq9Lr2p5tRUImpcZrYrn
pEd1srdnyl8TxXnk422ygp5fo3atN+Rx0Umx7RFQH3S83JZuLyZK6Stfk0DBC1DyCx6wJaM0PdM5
Z3gYXFFt4soCbXoTmegzDi4khmz2lvG29M4t6sV1EgBRBjobGm6ltok37+6FGw9rewkOrlwS/tDj
EROJ1eO9YBZEPDXqXtWzv8twlPTuanMWDij3fj6KtbqGCVOuTPrZyDAF7fg5oxTiYKJ6jIvwLG7k
Z2UIObdEY4LioOjplhCAGQ/IfAMuwftqGdsr8/4C+dbMN0Xov3eQW5VDDX5X/ejoH8PfOEZ/gLFM
7glschUWPSO8duXBjiZqSU/vXZxvkDZyUY1OTph6FdMmVS0IZHzaN3jMIarz7OaH1gKgIPritlmJ
T1EN3GS2zA+z1L5rqjTuKBRBiM6Bzwil8kMkt0zXcdgOXM2wQpf6h/iIYgJItfBFTca+0+X9t5LR
+1tWAprn4vuHnTsk30EyUM4odeaOk5LW4T6MVWsOvCXHRNBur4jHcdikX6wQ19WNTJwxezI3ja91
BG/8QwQA66ypXA4qHpNb61DjhI4nHe5PI2ou3DcmzhzAMKgG9Wwsqr1D+zqCxUsCVfg/MimM9xoW
6XpdMIqEaxXx1CzCL5CFL8bRscmjSdGjcNWcmgCQ7ki1/1mg5bYknQ/+yhvjv/nhr3Rn/Hh9BXam
w5+GvfUihQnz2QFPW7I0tWYdms87dAgpgzoPyovGjrVo8hxiidQD8IWSxa96mKi0mZONGaxbKNLD
mOHcvFflKbHiOT3foABaU0rmEWaRv+zsItY98+9BNy8VlPeSn6xusr/zlFAmT2429selvle7g/to
7axNzJwz6tR7tNOImt+F582mr0479d6M0leefzDlzHjy+3EA5lnR3VAJgI57d3gF/FdiH54loAHq
Uyss5oAvm7xK3jzzaHMP35M3b7Cw9nkVKofPbmg0jWKDr+0ms4NrtOWJN6YgYJEFn4X32/RJmqVL
3KKUyWlJlwcCDrxD/K3nULnCS7puk8kNotGdx7qUgExMBBN3QaFYzJwvCDLBoHo/5vUT4lm6BIzt
lwv4y79+5Pa6YshnxqtXQlfh129CvLkp+GWdA0X59aqN0kUuqL4NPIlkqL5S8illNCzfAUl8tQK7
NB14ZR9m0v048lKsiCmnxfFslubdm75HrkiXKIijoHU9AfdUx+peIcDMpRwXm6Ct4IY+lLMQrAMo
8JphqYpa0IF0WycyU2UQpnuY7uDIZlBCA1Y51c9XnU9ShyfqlQy7Rt8BVkqXUg0YRIUQEdsxH1JJ
8nYoR4fdck2KTtQnHsGBfBrKLS0O8WTur17wc6mSo9eLcd1+pipe8LE83Xktl9YPhaJaC4r8WC+p
X/UYcqRyings0d4QYR4BDf8jWADhNnx/arrN8D3QMKb5DZdyTDq/CxP2lE3DbKVpUTpvpG+seIdF
dGiDPXvkIXdqwgWgAkWSEYQUiWojojX2af1nV2+EL3OsL3cC7lkj5qE1dobbHJ9pY+UJsrMOQN4K
MbH3skSyf4pV4cJWIonQMMyRaBuhA8Fb7NrdymKgcX3fdB9seemp2e3TmeDurq6qc/UweK2jReQx
vyGZyrQSCqct/Mn4jpoU6TpuX1uKBD2zfnaiXMriGnklpP67QPObd3XXd92TAdn0JwKc28LtPZ9c
SWBdZSDL3w0QfnGSvSklpSbdIlj9S7qC2MSAgppcY9z4ZYTAi1zDh/iHdtZDDu0DSPN9NAlnPp/n
BaTLBecuU/aeWJf4GXik7walEXd8D4n0PyDkdPXZ9kgVbzGPZ9sWFnyyM5/wSLe4NhKFZWPMeV+W
etv0MVkwZFqzzVz9ngRZCFPdxGotKBo4JFe3BQBqRSZPjN0zewUa77MatGUn4VZNR5XO5w3qgrbV
BRoCcIbM5oAYSSvEY4nXviGdrP5JOJ8GIL4DPAoiAgRr+ARlMpCf9u8xUZahuDzuQbpEcgBHdPUv
2WQy2r2BaXn5ip8zB9Fq4iVtYLKOIT8uz3gDAodfTWnHrYIJX2Hd60JAMln2vF8iuxtLAnb9FmGu
O9dBpSFO0UpJMglcyW8a/sf9AzDWZYk2Kj7X0wZd2q4cUf3mcDF790IZWX2K1NN1dGqE2Sh85Nr8
C6u63XWZxajFj4kfj5GCYCXw9ccHX41eQLIDHkxbvKpcstRcathuRfS1cut06sLi4oBKpOil60q9
A9X+U+lpGsQiNkrlHqBOZEuNo+8PqFBhp2HcUUky/vgHPdTnhMvToXRaP69QHKC+ribnsIs9c4I5
RrNdlgDEEHIEinEf0cdvT1KWCaXIYpeyNdWavEmK6FAkxrH6UJsWYfoVsWgi8pgHk1oVkCYmto14
y0408FG7CRgggvmht38fXqTWxbylvmVo15BAye3dXDzdDvPsUOK5oDCQMb233g7TLKlkpOSvFZ3C
yULZv9Ai8IjkXSzGkL9H80W1fBY1UeIQdfnMJQ6vbdAxv3j6N5gSmNtNlbBV0Zc92RTl2Jndkk0+
sBp4gvBAsDSSPFEyTINOzSZSLWEjdtwoXWOpEtvVfEw2VORbDMvXUkQj0BUjquuHo+ea6LkB6K+C
sNZ4CLmTEcldXlmspa5/Mw+sEHobw6ODvT11KEkHY55VM9YnO67aZMlDrt7iDHiDwCGMiGbQRkYn
9aj3gBuiRX9YwewyxLKUlGKwN4QS1xJNWS7TdtiuHau01MTZe52V+zAQ9ZHxcuczPDtMTCNUqVgE
O7yZf5ydym0C5+OgP3mbzm/c9Vkeml1p3k2TqF72l/fvaalyWlDZynojJCR4GBMP05YLAZsyr1eP
tkjxkpnBzePPKalAS7Xk+VRrz4s7mdXkOPRqZZPnWvZe8E5ulepf1GQHL698IbGUvckJgheFHD3L
9jx94VoqO0C8lEPKof51rvFWEO23noRwEYJGJxGZUhcc6aOETMi3sDsZCOI+b7BlTgCkjLzg0z++
To/Hnr0dFCa0vG4fwUSG/neOsG8pm2UEmxbBjWjs3x/B2+MCP5NGbfYGn1znx05scZWH8z4EGJRp
uTar5WNN0c3UwyOkULFdQzypcPFlDWfCfqz5+UtFuTw50jfTIVYrvD6hp6lAhuqYIX462ubrQO3e
wDKUxaKw39+H09lG4VvMSUdBuyNheC/4vpwvSIV00n7m1jEC/POHwUra1+Mcqlhulm0mfIya7fBX
gOGUZjN/8EQQaWheojC8J80q5lctPSq2sc0gL3Q5qMVwZGh6c6pW/SHqZtRmme8Rb4aPJ2M/UViy
wP0VB0J5Eu7usJ1xrouebpwZ7tPSiprtMWurQgGaynC10Tnjf3rdL7PoSBct3OGTQ2OxGctJVOyc
9EIWRQqBwAhAFP0UfnpuVMHby91rAXYChIeSuReyg6In7z2Mw+P1fagkU+YvKqK8lU85nsdY9vz0
GwPoiFBAA8UKUqDArI81jcreGKM0FsZpxIXfu4q9bVWsGijmvurCursyV9//pWlR9sc8swN4Rre6
kZpjIPiXnprbeHnN9Am3a4I32YGqqE+8xezGedVJw1PtSUISg4yU6w+iHZ7Yz6ZFGoY1YAHT7ThW
hKh2MHGA+xUAgJn+5bfBy3iVde2b8xdxYJCi7EvB7l5vPK5qB7/nkDQnMx7nKRJCyMFBk7c+T0gn
d/jutj/akfeVaZOZeCQdADys37Mtvob+pPvNRtXTICu+dcgxZeV95FLuE6mCtbos59onoVsx9oNS
q1IUE0RXrvSfANDyr7pwMDmafVNqVlKWMp5SPLvEJMxNbpbWLOhvcJURbjCwc91Ai3UZ+OLddpQX
Xmtv5A3bxo3x67m5kw7l3OtZurKp/jYo/khpJV3xVD3rwB7lTQ+/Ek+y+/FakAXwAoSPx/sK63un
GuxmmozDdvkAjBoM11vdC3EPDQ41y+8prxLYFX1Tgr5Q2/05catHiWsQsBtPZKcV1/dphNs4NF3G
84IgSygdentV9K3/bwHwGauVtPs5g+CPKCph8fo/yvf3Rqcoc6tPTmFCWINMEtNyQtlehpuB07be
OfdyfZfnCi3qpGD7RzWrTpiGETfrcAdv+lcy6hygx60xA3WlGntI50iETlXGINf24th0gkts+9XI
yo3L15dk4ReGmCgQKWiui7/5ios1WjXqAsZXO7Nbau063URS9t72yiFH8DmEci5BbYT3k6nHDUxH
wMBPh/aT7qx2P4+Id2RF/ABn/Grm0fpwSvuX65GN4mOWBsbTN+OBMw0Qxy6Cp129Kpq0jzGs6JuD
VBZ48UzVdAKyCdH5dglMLBrNLZoC4YSG8FWwMfWyO67MklgIykxQOwJtqOMCLcMluwTwoqKvmxy1
Px+oMRQ6ROmlQsfwLv6A45Io9bjZvTdJ0b8l36cEQV4US0BqcJ8g+qfB3c6hBgOBZVIGRL+wkCFZ
ALfLR8SUypm0JwcpgMp13xziOupZ/aaVPN3d8rSXaqSee40qU6vpILDdgDPYVpa+0dJ9hN+cgyod
WrIsFovVM8n2LhJnCEkZ5X9jZOA94xw5ndHK+faYurY1UFqAo9s4nn4NTVmk9WFs/PSeECv2Dde2
Ykz00vo9as8jZBuPhbpYpSzRI5dmS9YzncVyHze36STiEnjUeImbRcc1/DP98Br9ob9womwrf6+a
9UtAjOERE8yOGt2U6FG7PKWnbyp3AXkS5xiaItU6pDiGGCcQQqU47+YqaR7TJsNvF9yMBj1y66i6
JVHVyO08vTOBks6G7lL+lRV3xHRkFQjorBvwOlU94qGotW6W2kxbY/xNIoDfSk9AavsYLj6R41cR
TsCpNOIFtII2n+8BbRi0MpsUAQHmdtT1PyzhPXdWSS+8Z77OoTzJh6KXuz+bUs9MIBjYEKoMfxjD
hYbSrW50NchauLmoHS3sIzmkqdukgR1QTITkX1GpqvoGldx99t8/IPirDley1geOt7hA6LjBnzhs
f+FNce75ActgjnDUJbRsc3d0Hii8oPYGQ8GsU3FPdJwUn4JceCu3ml/g40XlHD8z4HYPTJ+vdzRQ
uZoxeejOrQg1Jzg9UFipMBOV377wFvoWtreIRkQ255/H34bucqiRU8HQPNQcBxWnTY4xrj5GizWr
AXL+8XYEhfS8Y2muaC2Ti0tAqCK87oPxF4GypRsgpAkIurcLJph1eaTKDySM2NdwmbNpIF0f2J8l
83m5ReFQJovx/nEmkEplvCBLLHFxngyjG2ew6rju9KIrCRcz8f3aU2FNdeKflS7o2OP1qXXBeU9V
JobpU2eN4WaNEUVcCc2eEaXYDyDy7C3K/2x5oO983+FhpumZxPXsNIozjfF/khf/sPrLI/B8AccX
29xde4R0hGGXQI2yc23rA9KfgOP1sidWc2/PyIWOssfbtIhkZpNrsb8tYjkAvZXMx/I38xHHwlGz
+Dk7eMMeXcqojp4ow80GYI/7SSBDj1uqPWpTzl0Xcts6yxtsUpF80DgL/BQXj3Gu3RoskRAmOptG
eSqgwWglp6uqb1VV/v15tUyzdpE2g9F8MUXnVPqAF4v/E/nPpUQEYjFOzgQNoLDF1KC6QHgiNsql
JT0srTSLNHqUDGwKLUoOHxn1uA3he7t88x17sdmoNbAN2iKt8d36prQf5H4XWFaSqG87M7WHdbjh
zP2vRK4ym3Hh3uv55d/ppW5/BZziCvgn9dGw51RA097tvN6mIzNyV7fWXJVesYuiQbdClKP84/YW
mYsI2J2SoF6UfW0D/jVJ2JwioTzK0qrHqgKX5fI+k2mj1DQbnpSB/kGXqT/04657V0fh1ZVRsvN5
meJhoZhmuclhR0C9qIQYBK0axDQw6Sh6pPvWvhHeUjmT/JtEnku0ZnFqSh6SQb0QUz7g3qT1BD2f
oXPd06RLXrkzzM4CLboM6VK34dmW9dVE4w3oC0rZrooCzUIcvlR9vDGuyQQLNnXvw9a15wRfVKSp
DtexQ0nGk99nzmcTy7XxirnYgpUwYA1947yKnlmPTEbmPHB7mlhV23bx1hg0Iik7UV0O3XC+ZZNg
KvML921EwYHVzUPIpAmSpnRhEiHbyjCLpuhRij+iNJoYsgife7b4CXjKMJofSq0p0RmrY5eWa8+z
+J72sVzvCN2x/uN+SRlAh1VIJEob4gPTOuyxMa1J2kIYcGFGcMJHgy+Ou7AzFKMZ7FJya6yq/VuD
NMNU57X2ZBY7a/+zVRWaN50TiG/5TZ1xmERQkEGAh8nGSq2EX96q321uQSQQDLiBpTRjoK8xZyn6
YAR7J8kRH/kKs3QzfqaqSH40co6Ti2dXlw27SYFRi5v7zq28RX93+BhsIbYiM5DAZcR4zAej9SZ0
yuyyjwdafdrPDYnZRksO8WPlIfibznGDMqZbc9AfIcodjXR56b09yUsnp00AmoaIjy5L7l3Jsi0V
wg1wybDPIS4Ewe6g5blrhrG083hZFI4F6/Vb++HKuM22ngYsp2kvzdY4F2VsAJDAlNkdvkEJMC1o
sPjpq0zgaTK4UIiQGGstQPO3cww+l0utr0KEY+X1KVP2hH4OHYt5t68Xb3VCT9qLlUahvehXWVaV
LZvF5fC7ry/OHmi76N6V1c+Z2zXa3vopFygMmDpHNhb64B+PJYwLCLMbnS5qzdYHg9VN3lWjqaAt
lioVomd96yMhY5Fa5jmZRvkz5nWlr7euIwaXWFVGZz5fxUbB2QwmYLCwSzbcU7KGBm+UH+eyBxEm
0zdguUn/+KhH1l/7Dsbw3oeXv08fB4rAnwAbxhXnNhxM6Q37FHDRhFAJEANj/mhE/DNvCN4gaMjJ
qZEverpQORl7Wc5IYAI0GvsEnFkiIIxEEVzjMYBza6G5bJGzivjdFaMmMcn3mOAMn51k1aSiF0/n
D/I9eH4EL8N+vrREw5PL0bCvnts9zmO79Js9aVHWMAbfIA58XdQfn79RCGe5J948Rr+C4uwBQiby
+LcbjTHW0mjdIQOS9TuxksGhaabZrcturu66tXvRmMR2951yBihXakMzSVcIoygpTW0JKtRTZw6P
8sXxNb6VFrgvB7ZM2gGZkNpbslRIH+4/8pVtX6Z0O7qEOZxbQgb5crPZliX0HkADyV8gsKyM2R2m
zJrbsB8+7cwyID+RZ8AcNYoJQaxohFfAUSTej/E8v3ycP86H+L5QhprNQg83v/r+QFdGkEJ8Eao0
vTfutV7bp5XXEdeJUjqY57PrujtP1WevQ+osUz4t9L/BVL5NAlMqMlxnPUZE4Hm1aalvoY0jR38r
G/xQlrsAQ6JqkFF2CsxBblrFPyhzPCXD39nN0DApFj0vDLDQpCo+aO0zMJDWp3FIcLgGShZ+xrD4
EuS7NUP1/ZDvg80Uk5F8wBQ5KFpZCfOMZa7EAgrORhb9eo4f0prlXwYnmNt/mMoKixUadyu0DLrm
lXHclgp4aJI86DNgzubu03QiI8UtWYjhZ06QVEzN9d5jxRP7TP3il63c99dHHYp/3/aRVWhi2J/w
CP5vyVJhJ67ZNwXD3kBY011itJqWYJrDmQWGZgjoEXFqhBcss+1B4o6pSNvD1149uNJp6CkAb6Ig
vmcsOGOi4BXH61PnLOOT5WvI89OB+MGwVFmTHUyHEukSQBEDAj0FGJ67gCkSjkH0/xItaDlq+o/I
b/FXUpef8JxXUVopLdaR88nBQv5ynb4vLcO04h35NO/XfTxubEAsUW/GO4cjqsDjHDK1kNlvFB0r
8Dcdl4i8veVsCGx3iPoGm5GmFXpZ1fuXvFH2hWD3ou1mcfR+cIUiF4p+6O4fVv54QylR8Bs/lPGx
/NX6BkN7GiRakhBxGrtLIJpLt4aRkP8t9b9vRyNX8ev9BHH4NNdkDJ0JsCxR4ZKnPVcZMrSpDW2v
0sEHe5gUVTw1nCVKkMKW1/iYl+gE1yzXn5oqFzCZvnefTf8HbadtOIFbvX2BnVuwgaTjbbfmC1J+
KnNhCn0YdU2dGaB5WSQxMwzjtEX0BPyjb8Wv7YZx32LyWsV4iPG2fhGj5BMgthrw+hyoZYbWHXkP
Tb6QnqLC+mqVGppubybTE7pMvyI8+dTPJ234Da6fXTfUXRgeoAmR7HhWXMjw8sZwPBRHId+myk0V
GIR9/PV/Z/kdJH1tQtk8e6mgD+ur+ODpoSudZxrEVgeBCV5/PzVAe6bvBA1v2bgj2MTuPXNNYd+G
GDFddfnUNSE/t3Q2AhLYeXVITM6r0CuYyEKKNbVmSHunJeWDE+f4DSDgRg4glneUXqhWVOMsqiqT
432kMFMJotkyoev3S+hm04uIVyruUNn7D3iBzvGGSL53cdKSJwOg1skdayOLoowLNFJsIX823zTw
UcIscU25oM1RMgHxt5J4fvclES69GmdK3InBGsgpHA+1jY3dAaqiEGmIESfArQ4xk3g6aJEM9Ppx
s2rkxQNfhjHniPaiIaq2RWfW+WWLCl5nPxI5ZkyJBfGYJHaCSlkU8qKpFsturO7hFPgXAtOCuyMX
lyLqtEb0fCGncmiBGMGrk3WZUbm7K2NdvKWPVWKkgBK9QLQi+tmGkZVXAkCq9bUh/0F6nK/KZc1i
C0+Tl/ZeVIC7aeRvj943ipGRHQVXJ754cSkVwCvYtw8ddaFaccS8UqW48LJ3RNsLJWXylQaoaceO
Z7/ZZDTjX4Bm4mwHgKzlX1U5l4rOcmVWzazdRQtPQJ2Vm8trkGUe0ISj+VRdsHVDAvf9JSeYC5h1
0MTqxCBx82Uuy/VUCnYV+hHH8lgx3rHipxx6LHBR7VjJ+f8wWRW4Qv8x3c1VxMsPQgjH3Bp0iLFd
Dab9CtaLL0JpQbbTv6p5KVwQe4YCwiMW6ywgifPRiLM8k8PrR49lzkpNow4AvWDvOMKYf2xCmJBs
AQ888XdbeShFItebFgpeCyCNfAYk5aakCULAsz8D1ZtoT/niHMIjGJoC1ENDiDGyEofS9dNUjZU8
k8LlzZALrtWxAq8+S29gXB6dC2jyB7+bLarYau9BkiVz49ziO7kkfPFJt8bWoymZzlWERIzqUgt8
OO6LIIGwSXvPVhcMZfLsu+lVfmAlN7UxDbVEU51ruzFJHfe2MxBRdaYbB1NJikBZRUly4suhkE3G
Hv+nk16N393rkeQNq4TC/fHlmc+T/eMqBtWVk3F3zHMa0wsPQmahS3wS64k/PpZo/MqYWATb6PD6
xYNUJJcVmFU9+yZXNvIrvXGJ8j6Vgc3aPB10K8MzdQZ/wqhvNex9u9ImSPrfgypMSZFgaAdXG4Sv
S/1pbulc0jc73HmyGfYQ/4CvR1qtZaEOFd75gx/upDXcdqWlI5bXS0JxzRCWFpGBvYC7IW5NGhy/
By1sWBvHmD/goLPyUdqWQHtSLPMn2k61ua2TpiWbAxPNQDcUVaoAjKsvIicf9fsJJhO+HaoOh6CT
8ryj+cNxoJPbELabXNdYQ6dOy83vEq+ybRCSAA2RWWxZqGwU+QboZCEnM78tm3pFaMBETkefV11P
iCaAJWO/TiL4t7vjCZhsOI0EdgfIrecVKRE/HNrMx+2FiZluUfW1cGZg2QTnjpIkJRq6V+vJNYZs
7QXytvsduPB1Y8/LMkiGueYxDvotYwAC/XfnQLvNDD4twJm4gAv/xIDMhsXsYexqCqfsn591CX3r
0UIfTZeg8bzr0Q9hf6Y95JIXdNk51hNvwsKHPUKoFROxsP0x6C5lCUh+EpB5lrmMzEZKUcYa+aAg
E7r64Ywa9TS0N2t0qZdseBRUQo7sq9gfwGDKHzkOpMSQgCE1u2YPjM4ogA0GaLziPbUEgRaKWJny
kAAEVN3RzAimLER2ZvdPgZ8ltNsZ5Af4JEMlyQIrwQra4hCJ65GpRVfkpWDG34kc+FOUqnuVvTr4
DnRLmyDZ3gxbIiQ+IkqYVss3VzwFuWOctcqy5KWFp5qxw3QTIWs/+WIXjF6hfasHiqYSy14SqreM
vxqsHYSZSHdaiEaJvSICbWi476ZyI84aJc5BiCXT5O1Av5dvbmWP8bbrXZmlhunHX+hUqQAPkRBg
hQQdBZK3mrzB/1Gx47TIUKCxxWlIX0Q2hnkrrDG/e6Oz3Mra+2AfeZDj1CCwS7TFmMxWNxaEEi1B
egjtLhZlSEidGf5VEf3qjkXrkpLDQl9unJhazKRxGVG79YRDH0xB3PwWgJKOzoh5jeqiGDhuuFze
3Bxmld5IHZGuBolNdlSj8iLxFWr8FE/U4UOLPsf9qlP+20kwyMq4t7Img9/y8JWRT7Ly9VlE2Fxg
3Be53DbaJ+hwq//cvb8yMn/PYvYVNQ3a6JE4753O1rQoAtNBk72XiGJHyFt95a/ZCCDOoHmWFhBq
pvNjZpkspOTBg1pUsuLRBjAmPg5esQKq5TPmzVbC5uZZ8RoZi4FmrfR+AVH2uhY98OpfyhSptlNX
cP2ww1p0RByDHthgKLGebW3ku1Tu5kUdI+zqcZvpkssuTuZzMFCWUN0BzMG5CPYD2UeYE6aOoXbq
ms5nJ0xTGmt1IOekpJKid9JsPUQBQOT18s4aqC1kI2stH2ckhYvYYLF5XWXTPrTqVPpzHDb26r6X
xeug8UqI1ewC2uadxLv51eA/VgLBxwmnMW+B6HpglBNqPqrApMSG0nKAgQCeJnFgC6tX4YujQppe
L64e80S/I91utKWZv0LjxdBlS9vG35DZHr5LMKbNtdKV59Au4UW879lezCwezAsCHnhXEYO5fSm0
v+hm7oO9Xq/a0VYkojBIaIKEH4PDvScJI5WhuReletlzfVP3Vw2rtLKi0YYxU3RPauuj12+8RNqv
nQg/+es4Z4+xjmJpQfmMuwH/EVtBkOLOR4RUVa1FjrmfiMxhdiSIzQjrCZRE+UiIb6kdYeznF074
Cmd8a4z+xPDEL2Y9ACUZo9N2LPWia4j79/d/BDIBMOZ2CNTr6OO0usGRIYPLfl7UBzjuIQ7TxxT/
SjO3yhlGwuHYZwUSpXRI6tsUrsGktUvC2puhbo7lLSrM0QhvCYOeI0MqaPk6wxx9rkI2aYKvJ/vW
9sZN1ZmXb1SyLlE2FgtaNEdBw3M8FCQu9N1bQK18g5piElcVZDqc3DJv+OjIGAgBoYlY6Fe+11pI
hIwqxh5JPMREtHM+CNTO/h+xwTIzjfkKI4cDy9UFWswWAgZ1oyPpY31hnw0D7EDnYPpq3wnUz3JO
wXPhNDs/0KQy79VGkKCH6UTaTYeQdo5tg4TZDBWSnpVUre4pq4QUuXTLs8MtYRsJ3GUcQKZRrwhz
Ka1QVasR8g9hccApPnf2ifry38o9gkv0o1nlz8Att7f/SV+AMzkVblp17bqhcwLmSow6UvkTVebp
XUI4vaXSz7ay4b5x1U0WxWbSX111C+Wm+B1lMN4N/oBZOed/XBuxqNERE+TxBolMGba7fvJu50Lx
NwP350O6vlMp3YykVpmjyMINgUdJbSyQVPmBOdmaqjCGZSunidg9ySZzKUXqvDx7dhmcz7rz9g6u
msdPgkifjEPdCNtcl/C2N4i3uhedH6IgKMzym+nSwsRCpYjr9LTP6zmtbNl31BwpmImX/LUJ0Jaq
N7tUsS5pTRpMVJ1MkgWu088/6zdTrPpvM4dndA59/XX40fv1lsudC5gmIkp2rjvNJCUY6tpODTCx
n6/6y7oSbANk22qh9jpjBnIEdspM9xkIZWxkG+QAFBJpxaD/gpf4p1fGP3Xz2Zu4E0V+OAa9xTwc
7x7qZuUiAHesxdvZxA6rhsHQuGCjSdA0aAf6hGiB2GAkaceHBUhhIndlyxEZwbW2ofk70nJsBO4n
OixKlFKhxBzjhK/zHYiosqUytmjUtAhQswMfw5h/Ze26OriXdMSEgfT4Hh1hU0XU5XnR4hlaXeX2
ZBcGsazc7dlIp32H7eAzhOZU/CRVEcCeEsBMrG8rwxRt7ObmiDxKJy4Fk1D19xjOdagJcmzHRHGw
FNr890EaMv9aaG3lpfmL5d0ez5/bcpbF/C05x50B5CTVRnIvYpw0/6NETfF6B0Kk8Fni3EtOVjYK
4zHOUiPeWfxyWbt5RBVUY9HMtu2oOTg+2+bA3dNXMLKcqXZkzrszVSfPubxm4rr2jYNuhuPb+pz0
zAcE1cHodFPrBgW1/lqc0XTaDe1d/SOh/EUGFYlNrGQ4Nx+lBxJ3dRhOntspAsKUo29nCeauGV1x
reQDt569O64SkJAM5otJc89rAsPeHvjTU8rEyDQVz5dcBWq+iLEy/3VfPRmGnOX2BxoeTA1RONnR
UZLqVclQebHH26sAHkY/MqGunGMIMrcO+rvoFZatyZIO+c/rN2dI911MsvAh7bQGttEfteF8/H8Y
NqGU2wIH2VOJXsAG/JYDNQQzYZ9KQ1XMK5+K9pnlO4COMr9KJ3d+891S/40SLVuwJbP0c9fAgtyU
u48HT7iDY+9X4RSKD0hUnlZgcqNpdgd1lc/1IxAZ6Ay1IRXHW5NsjoZ190mvYWIVCJ4ljx49/obv
u7coD2A09CHc3W1ki3MJoQyayay5kOkR2sxxngDdrgw4RPBrl4OXgpU0sp/MRoM4xHqvACfOzHm4
cXJ+ptbB5LneVSyK3CcWLKGJh4/WcoRTgUxGJ/Rpe1R8lliq8+ddBGUlpu/irzpWumi9GVpIDk4K
3xvVFKOKJSR/OJUC/T7Q7n22dI3/GtpR/vRkitjGoN4ZzznPqL6htPyFyxePxSRiBGv2FL8xcwH/
fpwFZkEQ5/Q5+ICX/kg03Kvj1zSI25aDMNFdWTt/UHdTk4KuBzVbX2YadzS3L92yeI8vCS1izbxT
VQ+xg+RNMjwVPA90ihc1zIzZ/mggE2uEmrMMgjS7fcfT/PBhfQXFuHUQVr0/1Ej8ULop9x8gY2JY
4I4RLU6XIdey3xgMpN/TACmg4vdjIBWJYyFvvLWOWj2v9ALSAJKDh5EPlpUuP9WO6kDa5W+yz3Zu
eKCboRL3I/4tm3eUUUdpSyHAj4uvFVirp/RP/iPWqmd1X6pPvSJFTipyaYDK1sMEuLsPf70NkDpL
TW9GuaxqHWoIHVs0kCuzudXLYELNahayGzmGlKsUq41ygpr2NmGWuz5qruTde7mu9J1+17qcrUlj
/Tq0jVSigQAENcaIv6P+GbyCr37VUxIdp5B0RJ9FK3wTsuRHr0eKEXi+xFx6tmpwOz5B+H/1Fyyh
kOmAt1XntXFK6IkgPVtEVOhbKWGd2d2JZp+Ik+egEnnrrXH7c/9arvE4tdJw/MZTvh/icx2gVShG
bV/M1LHg+sknsmCyHu3ytkaoDndWPs5kX7SGgHOeFEaD5w4NNJ7MrskPagVCZ6I/4sGCfuOI7XjH
QBhFg9HO4pf9UAGjrOOxPvJ9mBfJGtxUEil+x3itT4+aHmf+mBtqZlPNPvNl6pna2GnUQoHaN0ag
uTFlda5VjXZpkvaQHMdYsbyevj+0ExHjko6dZGlOlvrPwEdpUMOhca8YcPqEgf34V11tlDc/4Lcm
w/e8juVtscNik18ichhUXttM5uONjfhxfq0faTIbflQEYsJ4mkmvYCkCGH9PoufwNeb/K9X3PuYN
D0UMBzzOpm8Kc+HcZFNy0XAz1i3F71hqcD/eItZf6KZYf8SrFvocl0rR4v3XHwxBbmqL0iHHs91b
lgWEu8NYg/dzfLE84CH83HNIZ/BSTHVIKY0v4nhfUg7YSUuAzPhOA1xVktP0mUC92tB2gLPf5bGW
+8vMyd+ESk/FVVzk3G38aKbRQB60J5lsoPxYyh+gfVpJpusnQUNOM2tHZYmfVS7+TSQWU1nNH/Yy
z9Z5shkZ+OiEH9DVCa0HiFJWZVLkTMTBY3AtljLU2Ef1fBa1Bv83MZXScB37bfUc8S+TX3H5Yltl
Tt32JyA2ILJQyHRV21X9oOltnHpoG6H9KX87UpTCPgMPK7iRiTSLk1AvkqT4l6z7W7j9wlSEi2aM
T9qsnz8iW8JS+OmBvcP1JShLokuzUBMgW4C4WuBatZPKqZGa0sW6fZCV9OWZvM6GSqq23vRakOWm
7mekFoj4UkuhZ36iva02siTQ2LakY+o+j0uRPfxGzoYkuVRMbNaP/9OFIimkDU3umtzzgbKMM8xL
+Dx6oi2JCISUD0YYUQG7O9/b+vnpRdPNyXoDPrSWifP9ktyzuQeR4XPmZ7YMrCbvKKyeliYgFbOq
WyqcwJqjBgYnpQKuNrwUu8t2b1Lx78t8V0PMYoearaJP1NGrnd/qZWmhdO5vkkAogx1RN2gQ340l
+5tOAxJyXOQeaDRK+F9puZx3c2SWJQa0dsTGbptascYBdyZZE8KN9etmVNIphSpMZ08gJZ366gCz
SJOjoPQqN9GJD02QiI8To76lMI/VXL4ggtceN4h3C4a+Y77sxGiDT22uVZ+K+yufCQvXedvQxS7C
bYiYQs5tftTEauLBZBjcjd+dcQUdeiYzAJHndo3iDbUD3k/34XP/0FOBm0ACVKytG3k4rXrC+tRz
S0byEpM6PtIl5Z97wQ5hqE6GzZZcSqamcRWQ0M/cScRlPimqbjTMF1PH0Aq0ZLLDKoKr8vgB1t/z
KhOFuc8OdUWSH9jKdljFnv5M4bX/Ti+6r/S9kAXCfn8XkwF1poeoZzznPBon7k4uUKDGl1VmhIT8
fOaq16alNTalKRav2BdD7CXSe6ggRXqsX6pxGywxwDFybgcJFVKrpeHnlxsRwFQNuuDQnw5WJSOE
Aq1wzhF0xNxSGP387vjDjs0iTTr2yuIfawdkmDb0cFmAYKlpOSXBuMpYJTO9uiZCviOllsVRjLRl
D+/EdJn/Z7Kvcmyxlefqvx8cmxBgE7bhKQtsm7hn9d36scT3hMtiIYwy7owTfrJzHGf603tPFTvZ
l25A/Z6PZRg2MeB3xlYW6ISlZz+kfvGqtosbsWtJJhIRgV35zJvUngiv5iL2FY5vp0hxrOkCDxDJ
Dlmp3LRnRYxBPy3oYWlFm6Ayr//x8n0r6qHZvsqOL7pz8U/9bL4mpgJDa8zMz1VmF2lCKwuPc5Xf
ZWdC9igHksyssvoQFLptaJw3QwKNBJhFFQhBuiKBC6hoosbzkzYNzvwxJLiFgfknWyB+rtk//Awd
rCIESoKGvSTZeAPqH/faonAiF6nn/B78dZDUZNziP4+utjzFb7s4P0foDSv4PerPyWVzXuM2etSR
ycqDEKFp63ds44hn3YasGG2RR1HGGYApkWIl9BdZGm1WCj15wIkUAp9O7HKwQvUHq3xhYTrG0+2y
WiHGkwRVd5of//cRMHn2J7GKnTCJZ4gBuJ2kteYD2n/OAWXeJV1xy4d6/0R4C0Wx9/YKCToOLthN
Q3XT1Q0t1tOa31fXrLLcsOxNCrbWGpx4IWnfSkU4bAFzcVL0S9BYpDoIttUD4ESM+R2DmNscS7eI
YHFYdkY0HXWEEM96uF54o9RosLL2WB4n/M/fxUjV2v8qB86hljjS/Pq2DSDrVj7K/uQudmbcc/Wn
V5Pc/9dVZ248c/2G/KWrD8pwLC1xuVadbCraNhMxbIv/MArBS6pomKTjqxXkel4nucpEVnbgOVxh
+7emAf9qNK7ltgM4BeO07YP585WjtQbrHaZnTTkknk1kwfmWt9j90om5ttxbFvxJc/8GquL6LaoG
mpo84TuCDCf4dQI+ub73twnoCIWM9w2r4nFzxv/P4helRzbf/Rr6s33TJJGCBJdL8BQWai3jy0nY
XfYvdNHVRRhfJa+QEeUpDCSsWvWsH1pyTvcv+4jYDLxMKsxsEG+Cdh078B9DBAp9H3sVWBauc83A
8MvIF1MEr81/Lw+5WwK565mEXsT1oacUV2mmWZMt0N17YKrADDg6ugr29R53f1Xy+AtB9GlJIwFQ
HHkrkDFhtg+72fqhLouqVgeKZruwaTZL0v4aIxcc14XTKbo9ERAaDlTcAp+xpZLdPPlnhSiSkZxR
PW2MoEL5Uj/L5SxYPRNow1TGMCKNIZDHmOLwRxWUvQlbnPhg05CD4muKzv3r2Vnqr8wdoeujHunP
Troaa2dJWuW6oHlU6MwGQW9bLMgTmRjvBiheHf0zKEPOrvLWDQm+BK1KnX+ock4cbeBR6ISWXT4t
LTYy/CyYOtuXukL11aJ4uB9/PY4AVjuw4WO3uttIM2eefUcaYkd23eCB5x16O0u/VyPCHSprNB3G
6EGX/AbHzvcWXhRAQKZft7Y9XV/+Mgi37jdarApHh9biExl5Pq8UhN0F+rRHhOrZVuxhlGBiYtai
l5mT4BkhjbfHA4XjRc/JEu/WAti28TWUqlyTbTEHRC6rMiRKOTBd4FFgl7RHqG1Jn65uE/1NwHF7
5NEYPhPmfYaGBI7DS20FUgo3JIVMU/63WQCjIwXgHPnWlBV4Uix8ZN2pe7pRRDFtUm7QfargduW6
xc5Lmi2hysUx/SYEy/BtKu8hg9G2p0sD365I72bOFBsYXZjcGKmMOyWO6rrvRGadO+FmBhmuJmGx
fx1sh6v2zujOnZ34BokRLEByYraAlM4AxPqIbUREo7eap05lo7NpQ7A+wMm4/Mv7p9ifECczE3Ah
66qS1m7aUw74VwSYps/37dEtWtuvLkKTxXbxJaZPRBlqlUyenImmpKNbzZEPNS0gAQhLMlqnwmb9
rRuPgNR8FHb0osL303lArBQaUBIygEPlKopVxvVdUvfsFNUbie7TXVn49tkOO7/Px70y5RO7dXtr
x8bsURvwAz9gp4km+i6t2/2KcA6iJuCiF0XZ66UsIQZlKOkHfc11zZ4SghXnfRe2RNrYzxlV9b+H
ZWDBEFFeHTB/Da+coEAp49Svjsc4zdyIz3TYtXrN2aDsZYAGGpHmlsac3QRt9Cs/Y7mHnH0wT3/D
HnViXTRWON21FmQ2ZKqPtUKCbDM9mOsMc/Jog1Q8xTOihe2VbsvQEwwxgy+HK0L4iZKHGWnIgQA2
OpznqVPvu37POXIPpa7CAFHsRO8//gX6EbmgkVhajKaz0TsMPjTrsO8y6LtQBS+nSbN+lqueCis9
QTxv6TrFKrW17va3yIzuCYWXgQqayXmn4k2yiz+i+fg2nhLbJP9DqOhEJWLShInGOjPfot3++k3f
CJ5G6MkpGfK1NutVxlTZ/dtHnhioFvjmYzb7+0+AyZyA28rAgIe2ct+MEQuNd/uUWk5ufqT7Rm6+
EpwG1xXWKpvw/RsieU120EqiE0eoZ41aGKkElUOMQRGxEo7eF9+t4Q42N/q45GRq47NI7GyjNCfA
XqNwodVZdgSsPqmSKWHLWNMHo1zieVfuFnXZi8CV4paoqBWhiPb+Ugg/5yotomDpxQ9wg9KZU6w9
ukg/ftvwpDgEJQrs9UwCHpXO9EFJRO0xj0xk4EsUSiPUoYqJoMnPAHocNOQZA65j9UzIg/idtSCU
V0WfXmc6ETOTtIliYzXaWWM9zI8yhQsXJQtv0hDQ5k6KfS067YHEQ2g4kvEvdTKZzORxvvLtIA6c
tyXodNXlBVKZ4MSncWLLeYs4wSSmXSuQAoc/lxVTYQQXNMQagycGIAWn0Wi44p04m07vUaZcKoWg
qoMAATI19GH+W4nvPpQv2EI1COy1GAHBZJe2Lxrb/3AAyWqXHhFNhji3YMwVthmC3epcdqsVDwa8
5AG6U7yvZ14rv314souTylTf4qZDEv9enePg4uUew0Vgesw+hFJInG/5CsRt55I0zeloFms7yUNz
YMsIv0DNcc80nRy+Pv5xXbHhD9aexZA50LJSaKUuvlQKiZzh3GD5P1U9fVeMQ5mL0p2ckaE6ZiZT
Byi738gQbcVj362sJ8VHRrfNj6M1ZcAy0MqBCjqnYC3/tqzxhxP7/M3KSSwFtnO6DycqjZR54+NW
AR6PeS8/28CgGYoomzHT0xvSQcQvKHc7eSVG1mdHibX6uGqNH3qxjc5W8SmAdG7ipBQ1UAKQnk8n
W55IB9Ce740onTd60wAXQIordRjwTK1s/ZOk5GFMlCQstARCHFbebQ4I10qsrJMJ/KVJN8H/oG1Z
e8osnJoT9RW3xu4urv2Wfw2dF339w45UPzFIfZBpZnwig5+KpO6ServbHE6ijSsVqDxTaiXUCjkb
UIKlywu4HWm5Skf0m0x6WlnSXrP5sZpJw53Jt6SO2TYXIyNBnWB+n5QSdjDoqlMcUxLNoBW0RhDf
8kK9fSHWSnehXm62IISzu49fcf6pG8XwGxkEf3d27aIMGomihoNq1IJxuP6Al9AgzTDuSd2z4KOS
Pd+JxNg9IVXzm3bFOwVFS6nPFWot+7yv4Hbe4fgLBBukdCsPYYHpbIyKq8nKCAp0U4hxFaDSLM9O
hJraddgEDoi6+1NwEkqMp6TjmrcDublOfenJhBf5aTxIeuG3fZN0xiEGnlr1wbUhpLvIq5qr6e4y
Bwfy20rq8vJ6o4DbXUsVEiraLq69oZLXDvZ5fwVMbaUHoYcq/5IMcv8Lhji2BkXrYFf3d5Onbubf
iAFta9mNtpggzFQA999QPU0OKEajlsGACGo788OZwP5dDwzMtH9fmoadh6wazqu9lmq79oAhV3GK
k8sdIYq/E1CtFKK4fncYY4C45GpIyw0G0cO46Pi00GQtFSwLrKr2VY+0IFHKhTdqQWMBSpvqhfS6
7Cs5W1F7j5oX5vQ1x8+l7n2lHjSpNlQGz9dnxZB1tTqTNrkePs0J5DMj5ux0B98F13sOAIfJ1WHi
Ahwfw+SZWWgqPE00g6+nsTabtiFBvdQ8P5VYGGgvpeg+5bgvU3rRkNm/LXzJEvVElCQYMrdRcx8L
1nxdO3BznSefpQeCxPu+gm1CSXBEnRhO7HO6BUbbqndzuCBn7GmEuxxa/3cGTwU8WrGL89BL+i3j
2wQSSCN4tZz8ho8SgeljgDqUmgUQTzt6cOSsxzcy1o04zWB2sojFV/x5jLFCujLmq1zguwW1PS2z
q5ryGtqBf211IJHNne4K3yEWajb8raK3JgrjmcCLA8S2wRcrRDNEIr/3r+R5R5wVN6ygVrGknpTn
M23esWhIWihkI+xe54teCs88+44bKsuMUkUh15o1/ZChodYohzcGsyXnQjPCZT8e/gsRgViUCk0f
EvabzIeLQMTa1xfqHNIs6pHbdu4lIoiLObW2eoZ65yo81oe0yyAQDxLPnUMrL6KosLT6+Ab2rmqm
y8odXbMlTLjX+FSCMKr4HZOQL5pcuphC+A0tcfwMlSUIpFZEnkL0RSWD0J9vrbzr6jjBpOTYJlZr
1d++k9pR65q6eVMXstzW6tIYdVYVfG37u27PqAWkuND3mgHUM+sMythDATVPqsazXJVU9iStwtRC
muJTLW2GYMHYzW7AX3Goe7CM+g9K+kOoOTJMpOEG7Welck50hGiFsl+PvqVa846I8LrKRr24HzlL
+QQiW5oq+QeHeWKlpP6KRzmSeoNyH5Y3ecFMiONvPqAcrLr1fM+cRYfPo4zygb+wZjbJChpHCd4Q
CWdNT2TYJl0VE17jroaiKOLu1tXyH/R7Pr9YYxDy6pzI/7gqygk9/mF48MVq9oGu4ZHeR8LHlgh6
Q31ff8Qw7e8UBuHoSgnKIOhrpH5kGUiIiiC4U0tY2LR44Gzxn71cwDNNejF9skbtHLSjvILZwfM/
qtIcwg2dQ/lPw+6rTA90ZOyYw9kw/agLEWQPCA9Zkl40sBFlZoXT3MBMBfoTTJElroISuS+FfXVU
uF+BUynMhTCdHwvDxg6HOtac74XKRBr/nU/I4z8tUD4WwvgtoG5YpeMe2iPrvVX+sPFLo0WIYXo9
+CViP5TEGIA8FzAgBijWRjS2bIoQVfaPXweQmd2WbfwulWTOfR4AD6+PZUAr7/evGqvCkmv0aZvJ
7A8qfWiTIWdSSfgkI2m/E1YDMx1Q4F+ufOWZ4/oeFLJgsEEANOrDGXF/w3pT9ni+ygF6nvf28vlH
7IbdxrDHHHSEY2GQT815xh9D3rJ586lC/uDG3oPbe1ABZpC5YThzBPAZv5X0kbtlIpvKHVVlQX8J
60BYpvOuL0wi6Zn99jKyq3yqwUiUvVVDL+8kdlKgJbrViSWiniRDfrfrIDBX6bE2aa6+8Jn3/CuP
DKkoSKyby22Sl33NyDFT1R2wU4xov3yUuPdLmbQyrBEEEExwZ0L0HVH0o2zSEcx0Jvs8f7kxMW/H
IBFj23PudKqYhXhwe82c2b/KJIJpKlyQLSXqmTgqmSx590u6Jha8euxFwMneaoTsEiyub7Zid91g
T/gRYORToh+MYVoWhrytTLhzE+Abzdyf0e09Bkt2M0eGFPpbLU642QTvIg1nRB29gjvaXhlmBaxK
8JMMD6sfMIDjhagLo8To4ay63qYRbmG3/LcZLFDBQci1XHYucAGehlGpWUnIUFjSUWYX6DZGcF/n
V1MfYObqBMkTbbd71nFdyptPWUf96b+ujjPZJ0Pn4ly0PxQ3YarugobqutHaC1aItLUt508MCQ18
YmJK4Q2cYvL3V7WGfgSG5n+tiBckonJmA+7/MqZMFyOyWW403CyiG2sdRngSxhNj9kbEwJgc6xbF
R0n68bHXRoAuyoPGgZUY/7PBRUvhMZ+6SQMm1nGuKqhPUCONoJJx6nucdLRmhb0fqSIR2/0jiqta
no0cyH/gzr3Nm1qLYeyl3AgjCjNEP9HJ2Wf4Ccb2gqD1hC2evdVt+SC+IUnZLNfVMiQ2JfPkg4jc
K7R3T2VRAfWGsW86k6kjaVDN5TzhJSLo+aCaRU+KyjXJz8CuOOrZLA9bL0Yk+lgthhew2rQ4R/EP
4fPaVdRatL7BFpNplLdN5VnEL+hWrS7ZjPBsbV9RlC+M01ngHhDjDhQnY/vMyq1U438MfgCDGDRD
je+mlxmEfh0Fkpspk7QM6+7gE9+Fbs2Pgy5ckbAUNbVEG1Mq1DMV+APc8onUFbuzfiPzHFV4decA
/7fLKnzqFT+BEM/lsPQOwfI5+tFOqC+aO70ar2OShzMDH58Shd8Au1KOr9rKUFM5p9UokKDBSwsL
TqbynfOl7TetHZUxmH6r2ICXJeQ4qqVAM3Yk12fzZ2G+AqNfRiXCQjm/MnMBAncjdXEU8cVAkS2Y
kxaV1WrQ5+DYhADSWJp8mZGCe8y1OIKaOmYeQ0S8auLiejlZ94wxCvyYwOnO9s91JqYxnYkbewXO
/MxCkI52739Iaeibiv+XpX1iYQjt3g2XPuOorDufsF8CKENxrDmHdq6ihAJ9cvFDoRFBYIlheZWU
E4Fk0jIcVBnFVfZxk2ecdgpyghxGAcCNagSPNQnrD/kwH/LuWJQrP0gSwPuDop5iBQBxmm3TszZU
LnDoVnc9IGcqhhJFhQejzmThX6t0iTizcdbXuHMD60n/oW2E4qVUcwKANOp5eQTNJPzaGnZkC70g
VoMyzXIcnucQjItHFMs9FXmIdatonjFcVzTXsGGdOfRNgKthon9U74CgjNCBPazAPd5220hZS8gg
0+GimEBoR5ljmm+fBGBPhP8xC7vh6LiouJatbpaf2U1mJPBBBL4sEedXfJnnwnOa03PGbjOjvsvK
BhxYNf9eupLK8lemy60HlKa90ItdYurhpJ1QJBaxVVsfIsfloC+gJFYZgJ48kKQWD1ILG4NLYiDf
vjHb5TBTCUNFiPCQSKUVIYG4EAQ1dIVoBJqjR2kJP+h3voC2qGM2KxZIu9a42w5USn4c22UzFI3Y
iS4O6TPxSe5sECBdoRNBD/NioxKXncvGPQMNVd5QE95f8LX5UhGP3Ma5Lh7V92F4063Oj4r4bAdU
uqA1QPR616c3hpY/ScWMUL+3H+f4wXaHUBy9ReojZogZ3B1pk0FSmGq9onJlw4pqQvVY0R6xEwG6
EiKkZdh1dK9P0Lsl8WwyJ3eQ/lBTD5eiA1Q4ZBWFyfXLDJHdCz8dJEY8vvuAirdjJX5ilWqyXGZg
E4JVuF2zhn6j9hi2fYFlfoKyq5S6NdqK48adNOo/0venK1YuI4DV8wwKzz7bh57fRlYRldrErGko
Nn+5xSHI2lD4XuctxcgGquHsZJOw7Es+Ub+OjeZlGJz98t3l8bDOl889rkVSQwli2HyVMVC5j3yv
0vyHohSaVV6S7TEdZTZsTLWU6VyYzWFK+DWc11J9VVPU2iFUPL3z8k8W8NR8C+DZ7+2wk5Vz13K9
0aAns9M1DlrJRHqBKXEka8ydTaUqv2xG/B4nYmVVBnEWoDx7fQmJhSRxDIBk0fhB+yrKyRz/kQXM
yJmLTqjRnb+mTKb4gAt666XF1gxazWHQCuDTt7n1SThfBCDOAZgCNGIyL8lrfVJAHN1VBVeQNqAK
1L2sHUa2GRKzEjpO28HIdqlAn2Mha3DbrqcqzNlnTvMC0lg84Y6ubYRbFZV22AiumA8FLkfDUxFl
LvqmGqiRY7RNS2KegCNGlh/zMwV1vD7Ph33apX3MHP0wbZtUqbw3uqsmmmSb5zrbaf0Izyxrdp0E
G70EmCDObWa2gQS5avtAdAKZ2tRz8P/lMVVe+2ogIWfpQ4f1QndaOnpq5K9VPdWuSreSaNfFqWH5
JkOPeQ8y1VoLuieXkqu6vmiQ/zWxkeJkUbnb81VhifMnhmgumP+JLaeBweq9qkPNGoBl6bqhoiqc
s8sdwq/NQPrOR+MK88gBbzHx4CwVROPN9p+0EQ3WVU/Nyjvn/7mxufA716GvOwFq/skK6wAlwp2+
5gJyde88SegtHoa5LAZnu50h7etL9njacbBjoD1+EvxQp1T7v3RxkHf6EzrzLYTj0KxJZvDuP/q/
ksZR6/gKrQaPV0JMy8YzorSvHq78iVtO30K/yFKPA4C35jRJRKUb+YMQUmzabvnEP0u8uSe67s7C
zSl9ihn0xJ6RXRem4fBEURrmsVxD+G+uC89MNXWe5M1+PAmzAjaqygTNCzk48TSiqLuxOAfJ76aA
rft1pT4KpWMDi+cCLMLhfs/FvmH8yqdqLkA7xmV9k1B8oQZmR4nK5di0FFLmfrTMFO3GafjxDdee
2nWh7s3+gEN45j+cDzXsVOJ5N8O8l460R8WxtrFRwXcRW6gSSVEbEM+pqEHmWFRaiYyADcBY6vZv
+nv8lafXaAu41m2QNgRfcQ10Pjq7AVjbNkl2DagAIqgh9khELic+bvg4GgKwn/oO5RvLXEVPgYvi
ao5v/6oiBzgk332zMsQ3HRXTHQc5K0JVJ7VrVuga3Q/saHSVbsBRU52HZg9DgRzy6qCpr6VSIH+9
mALdnlVx4kjUuoZQDavnmq/yDMFbmH3ld32pMF639IAM2WFdDWk7duJnP4b05UELg4GzF9BY+ghY
AG7/xslUJ1MtH4gaa8t9KrSEyRvZevh3UpwjVaR1bYiOEFkwHz81jB0+9FLaLAjEGwiSIjekBp0X
/2sAj/ZMEf/BdmgxbKl+8yTOod6TohX02vSizVA1yK09m6ndGsmXg/P800+k+Tz9Ia8IU40DYWDI
nBRtKSE+TAqEVedf51ybp/dTzYyaMrymO38I3BSwYiX0hVTY45B5Kgy4d8LeCkBiVbxUdDA3tpfF
0CokzRYzsLYVFek1t4jm8PbpKJbcZr9fqbdwiCe32LH2namZ16SbN9KeuNVYPZHAE+IzhnA0JJCK
k7YttHW5qQ1/Yr87h9HTFf0TRZAWNUl85rwKzj/XqkUZm+9KmuX0APuvct59KjARzZIRQeiVQEbZ
GMROxR8Is9NlfuwBeBqMdTYm/0YkEaFmI2j0nVfQMzlXXKzKsFB83Tj8t7JAtNQRF7KyqXBsgmA7
uWdYdeE1JC2YiZ8NrDRorw2wEIeTTCg7LoJXF3hL1cZ1tiQ3gn6Bk/t7UroTmoSxdBhAlhYitAuG
hci43q6nxYvojxKHvKFORMMpfL6tinzxuzq9jxASSQleb5HGMW8CIlj8V94l3ng14liF/iRg0t53
qYT6vDkF6xak5gl3t32W8MhgGfyDOi/14jcqukqa2A3Ksx0jx3YO/fcvn8PRQsSet7EJ1Px/Qvph
Z6QUaEwhPx6TUpCmYrjJpx9LNqj60RKVxZPeUf+V9UKFc/F9ruL3ff32lNg0QSNjM19Fj4RQPGH+
7G7j0q4cMHlc4W0kTkTtWHNMKANylglUkK6B2L8DGLRBsPfG/22nTP26Fq/DKOhZDuVNlo0kWi/+
UvzNujEIWeOMx08mA0D/TxiRqLBh9dzLNR/jRtksLbeoYBuhXsR6uBkO1RNvttWCqizv7qZ2+DTl
j/p5/FdzjVqk7wbf2fm3fKHiLWUq1kJiUffP5CSNaEuip5G3arQsDkoBo51H+LpzWptaw2aSEfNd
Nsk0nGZImb9kPtHqkY21+hcKr4DIk8yAGJGSWv6ho+TkVFfQ/wtwSLxibKeD1eTr/zw0ypOpMJGd
3onXAFSvrNdDs+JUiDwP/uPZbTzzy4fKq+eDdvHBNfkkweyyfCJuDXyJaj1LP7d7/S9aIXefe/f8
NUpzKJJXycjubvlXMNvnb4SUa6fABBPH2+DpW9VhnN5GAjPZPxKwiMmWhLD2huvVb4u7Ct3r+yHd
V9/SXRuwt6Br3ds13NaysS28RNpbJ7FA0x5IEIRu07otcq/bTmtLpg8vFZAgXzc1oWVF15fTOwZo
QSCe++h6j9vFNEOq2bRhlKehVRkn4lunDU/s+Icx/ZJB7NkGQ7X1q3jWUoaUqhMMK0YtpE7BspvY
FY9MKJBbhMy2vT8naf4ivq2NatZ6MI45uTgVhFLxHyHMYBs/e6044rOAQqwZzMzfUj3+GSar/Pzl
fHzr+q+MNaYzc6cQi25IWKD5V5azEp7lX2Fx3SUABFDjoIHdUkYsHzvERFYNlxLz0/IooW6/PuVR
PEDJtZJyvcoYHXmMedCcGrGAa9WWZHR/6czNW50t3qEruDVSvlb3SEOwf14x7VV2hez6j7NrDntf
I7xximaw+hCWGiLJGAhkQTQ7dNfyzpFi69ej12fnHheK+LzLl1g14GNTa7Ghk5m6ZivMrIwI1Nle
Xwz+CDyw+fd08murXkHr12Mw9q4ja+6L0MrDHWoKGQ0Wna6MwoXKWltvA+k+oioDF9x47AO0AiZQ
ggGB8iU4LqfZb9lsKy2sVSYkQhH91RpWykuObqmLFOHySQ+hGblF5CfKRFoPUre2CEaL0d0dzRG5
vWw7CcRelpx7HU70MkyZ4UhHIcUgyYKeeRwA0qMsehVVJ1M80sRhUD8GG2gVhYqxj7DCT/mx0YoT
0HPsTR9dBv6OAV7Tw92YhMzJreUPHrvP/9D9Ow/UkgU76GRneHEDQWcoiIUzAhmNQvj6gklLdaS5
nvacvNrtrzzo0QR2kBY2chD+bvXJ0us0pPKInATw0rdABe/TFifZ8MgQXHvulXo/nBqUSYTL3p1d
9h9LQcA9C4Zk6tkXx3J/JZ0T0veOBqrmlnJjRZfZsON8KME82mPEMuiZfM5HW53OZIMualxPz/FB
7oCpc80WAWpPR/Jir0shC5ZhQCK9EDqqe8YxG+xo9m7NnueHuzIWaKtV5dRCv6vzOtFnJntDb21v
IjoVPv9nRAyS9muN4lfI2D1k4HL1KHyd1lFOSjvYzyLaIs91hc1BaDYZOHZggG0HpUiHo0GP9chR
aVL1AESWdbKudBhmXFSLbD1CpyMqIy2oIybtZv6RIVHo/WMjj7+b7wGl1Bk/qzWsp0xLSDETavr+
Ha63uBDuAaV+IZRvfAt4sEkslVppYgIEyKwSNg4xsJTufYKEBp9qje0eF1xd6iFwFBL7WczgXlA/
DfxkhOZ/EgejI/BTIBe3KTGgRac6SQXfbrKvkS0el9jd4Ai4rvtx6l/J/mclofCGRR+tx+C11wUd
gwqDQ1gMsx9GoaE9gpJtsPPghkjndEPprkZ7LuZjB1T6oPXeNrJtLLTLyc6Ggva2+AMZEdNMnrMh
bB3L+IIW9wQmegvgJBiQV9tU14Ml+vBba/eMqXZjjU0vCzM5b92RUsIvhBZyps1kEkXptWVbr9kt
iluUQmVn1RSlBRoxqlDFl61A7OjbOfESsVaQ2QpBA29FYShod1LCni3uwWl4fy/JOYbjTVq2Z9CL
00is5HSAxyNPTjinTRjeUKEagFuPpOWYCjXuIPxoq5fT5gPzxsomgrCd51DLSqdypSHgpGmbSll+
PhsqunXecJ6qqA4ecqxgC2PMvtO0RlAx+oUsN2aj29org4A5g8qw6nMNkn01FV7P6D3AZ+dfg3Y3
D8EB2BGuN7z+oTEedJDfarx3aiNNmUeYvMXAlzZGnYA5ynEulOzk90IoI/AOdlC9n85VC7z8irBQ
Gc/mqW5QeQe7t9JMXVk1SF5PR+lVwDOHQPw+KyauhmYCNx6r/dYTw5iaY9eT0/Fd1NBESu7pueDs
kAoKO58oLS0TepGECzJeNu9TNyys87hVzzSK/kB0TWBj3Iynas/sgm1QzM4eWDXeYBGr2rpsMNnj
EevcK8TdAgqZbI0+pYq/fJs7OWlUBCfjPvP3UDNfTxa0SIES1BWTqMHAk2JJCuYe+ou0OSyPiC+g
y8+Oy5s3G1WAUR3ythJvSVdSr24pK0SBOZ48694zRlecd27l5awIZpWtmdAj10oVEOFzcP5zgp+1
lHOWB9VdSDN+yWhB9DBwa5sMp+yuiCkox/iW50cF8kr+70rq8G1FfngLQChzAN8ZH6cjf5md0EAG
3MXk47et5hCtoarDTqBt9fsXLOEKoO7HZ/3739ojQJ7lkGCZ0zGsuOEDTaXum9NJSe4p53DxsooV
adX8FZH2wybEZuU4j74Sp/Tc5W7W7AnqQkTzsxiU20AV2eiDIR8VqlJMun7W/0KrnGjwOkTf9mm4
2u8y/vmFtSrGKOB50vIF2eW7mX/fooOhFWMtv0ujyT7DLO8V23m+WScFuMeczg6BEMn+7lSnj1e/
bK9Aig0k0eI37DuvduI3fEN6v+2oAsgmrrKMpJ/uAZV/KqZw0g0obtZ2qwvcMmdTavQ2Et/n5Jr4
j3tAdF3aCrqt371EHTBILPprv3Q739rfIs8lkR8dKOJ4FNGkxtnE1VkhSqbSpfD5gP+jjOSrLUtU
wIN5rEWFy6VxwNVspPjoWSzsSo5nlPTwbUnzJpuct17XcTVAP7L+pFbPd6roZRljvhQbq8h0TRNK
o9qYEV2+CudkxJziFiS5n5EkAkB5CozBMXQ7cssjayQAwWXbgNxn6q4qBvGzx1Y4RQT0ntDctxVS
RMXlnl1sAtxYEePThAZc2xcXLrA2zlXK/sOxVKPMjaSICVBfssfBDoj6jaEj+5o52LwmyVQm5WEs
bjqXJlWxuRvw1p5oJI0A6uE40JPxD/lC1ahuBNPvS7QllbwyV+WN1PHJrnqfdzTu2N3+t+W+Fuoi
Yanamtc+lt397Urcska4EbwyT0MhGwU2g+ZR+wGfMlMVEbASw3x5/EHBQavch+NNSxfCAP0lpdi1
S8MEjov6359xOAwxwJjE/wspQpm+MGKXKb5rwabBUT+3bGN5j7be5RpD3KOluPlISZEPFopJRj6i
7nzXzBXvDqkFNFP1x/2SdBoxvoY07HGRUn36BSN6gYP/Eh81+0tdY5iHVF8MA3dNKxh4byq6fJSp
vxMkwkmprWlCHmxKphDdjvMUlz9O0pQ49AZy8hNO/7KPDm9IUinoGEV0uKFNFdtyhIn4vcMO7Z2a
7722R2pEy7SaO1Q2wUr3251iN5fYYjUPgc3w61i9GBURtRvZ0KdvKePiV8DjQ3uHl8eVptsrrkTO
kcDjEFlR84cv3mdt4KOgs4sEu1vFvLx3SPos4cLyffelXuEfjPgoYwiqiVG4enPs+aJylWzqIobC
1tK1sjcvlYkblSj4Rjsvb29Ha8x/ZKsl19yarF8l2skAAv8Jf+aCJoDV8GSItQ/5cFDLCPzERWV7
ZXY5KT/7RHhKnC7bvAYc0G3oSsXK0r7potDsHvkXwuo5SPjNJZUkHnf9qFZmYbv1k3S5qZAT46UO
jtfnOdM83iJFePCZq71VBC5C5ZgS2DmYS3glUJAcbnN9iPYdjnSlBeuJ2K0y3ztiuunLhrk6PG26
i23giBWJhn1HmYdY7i5p+zpG7TQo9Efe/H5OdDdj/NBwfbclupROT0rUNNgOSiRs84w/woRtN0q0
jL20D8alJ5jT2BQXbJxtcRYurBjlVFjrkf8njuLP4tjR3tcursoNHI6qRZ2dutqTKts0KgDQtgQS
/T2SPlvTs0rB/1a28Kg1w3RMHGFTAMkbQJbukRv+TsEV46Txy3ZBuIXQA3TJ87tiGHUmP4LpWaC0
V59X4DzEsDWgjcstyARun2VIoOcVjcOCPynbxOo98mf7hGchcEVYzwSTKPxYBt816qUqPMeFu3/L
ROXso9omJvxt+P68ZYEYhnykJPiAW63IMnnXHblKZBjLUZoT3zUZQj9zgIeNWYy1AHjCBd+OUPQ9
SMCCCGR5w/M5MB97yDofrZQEdXzY0M2L2aOCCSOFunWAaNOgXJ13PtNZD0jopYCR8uHrX8vGMh9Q
k036I7n09g743lYSxMvBVenm16v93EJ69oNQ6LI96IzHiHWJGqotg4iHPc/AzKIqoFXIibj68SfW
r4CIfbJQDaeQMf9itbCd/VAzUt2fRwN9RzWmDUYOanPzplGGqZQOkwxHVxun5aCHv+OSMLxn246G
BMUW5dFvrwGSJ8ajX0ObM0AV7g/eCThl15v6nO71urCwiFJFbVLyi8tBIfezZMd4dj1ZbWhipalm
CRtH/PaeSIl2jIWbXuw5mFuZTCPMocdNN+ex9OsJK8zyWpt+M0jiQtbu95OfUbpOYYvQB/7M8+9X
mv3/A5vhBo9AGPrBBEjUmqQ/kEdAXVWS0tKn3c6sIjg9Sj1nq/jYx6XK049uBH4cYQIJQIpDjMnT
0OaktBFf41T/9HS3TSahX/8KC+bImUeojzNSetiO37S8nuAD91sWgK2xPxnq2avz8L1RMv0fq53j
N1LUWQNQ7MDjb8f0lipNZPSS6qy2e/qD8S0d5PWwk7Gq6O4ai0uQSiKuPlVMwtu1gvZ5oEnRmxpG
rBFh6c2VgAKrnvMnUcz8o3sylPrNBY5YdzRPZoGTXthqwWV45htHCBLBwJfVV0SBS7qS2EoHXO4Q
VW0H/vIMPsScss8i5QSri0jVvMTENxVeK0y6RIbfeDlcuw2/7PFrlifbGWvq9AcQjYgCqrDpM/60
Khkzc06e0br/OHhJ/C8klUVKNH54vPzNUmzur1hgRe8gszFAydS8TrFqy8S0q/2HoXPmQGMi18XL
5j/pDUHIl8fzIXXRa1TcrgKU8/WoaYFJHfyU+kZaMR5PzPYnP2gk5OYfyazEPdrPyQ/p1wVDmx3X
1Qqfvhg9j//MNGXpLgVGA/0e0iU4aWG8dbhNylGm7/swoPN80Ru2tG+U70/OQew1t8bU628q7DBj
Gb+DWGz5RqJzzMLeUW9Eb6UVbCKWrdcJdtoGMpWIqZ7tlOuKK1pQ8/aOMuDlW6pe+/P8t2YrY90J
jeXgFu4aN+dkYcqT258LLqko8PneADKCQjJD4akK7TN8FjqECSbz1my2eFlKniCq2Rxfs0s0s3Yf
r7uBRECPynCzk0oarTjQ2k6EEOn1OcAtXiPleRuxthyyQieZ5WUgVt4EPP+kITjCPq5aVI/6hHO5
nvYFQlSJuyOlQcOBFvYzpVhOe1FogH3ED3s18a6yI412H04PisnPHptAOrTM5xLeN249UUu94uSp
vWa2UyXnHoPVFtO6KsEu9WaG/V0Uy9YEMReFvDlJ9z4AX1yViZbZBg+QmVRBuOthbrTAcGOdxdq3
7vapY6MkKXNVcNZNdQfQfdwdkhh/1lmxrUhx4G+eW/i9z9/9RsWwnH6hIHaIZBurnPMGBs01WLyo
xP/XZsWJzEOcvi7vQlvXWir4gxUFQrBC3ZYSyplgKwxegUcRNKlAezZx/kb07gPHyuquOnSwwS1F
js07ccVczau0Zt5z1S96HWIHjfS1914fyFE7WgduoGPhsJwwMzfSVXITP3t3OmcPJ2CjHIffoC7b
cOlpJgpMNW20lZJDoUGv9lRBwp0BJttSszFyZxNEebN6LFIAPLNJQYHhy0V1iSz+Dgpc6Wn9bevu
daZXRAMT6/rfIuWFVfoC4LjF2gl0Jg91Pp8ik6MdIRNs7yWqn1JnP198I73uAiwjz5RhxULlNRSg
XlT5gzlCGyurtJD6IPnWOyNTUgISiuDad63IqY8MGgvRINH7x1wYw9dF7b5FOL1kgk7l9fsQ8SDS
11GOx7qqE/78JkBC6+2W1xwaWWZr3Oqmt0MnQMXhKx7JCVuG6EFnrUVWqCkE3F5i/qOwtzTfwk8c
njykWaIB8Cdv7Yly+FmWIvS0sqTrTdYmJYcM1IROWm4fIDZxGB7HVcIBHyNDo4gGN4Rf9A88URzs
HSAyzFQdsoD/6/HAI+9YS1LDJ9vLkn+7mLEWe5VcOxh0gEp0TewB422NYg79rFIEI6ahq6xLMY4J
N4HqaBzPCW3RhU2Ej7+cHNL7d6/dIIms1TNVERdmp0TMCub+km7Ko09/8hjnX9MwqU3bdTivx3xs
+DdNvVYv12Xv5YQQMIjxJx+r6w/hyklGKqfqmcJNUkg52XCngvfkonsg54jq4GZdBxnqEOb37Htv
k2kAEM/JaA3AN6eaB01JegySVlcVW+n5sJ/bOhnZ8lQPpw272xUYyUjPoFyviY1ysTd+KbwmvqU0
zOQnDeiSaP8HLgwsGOkjpeLhpbUYo93zwQODdOVq4tSqyO/8DwEGvCVOu+Cah6fQokfQbYAEknmZ
IeideYG3WACBykiTqA4g7P5uSMNuvWbhSAyYNNO1olpEtbcGq1P+Hz1pkTJsvBBX/CXb90FoyE8e
lvdZzLzX6e7O5fkljUN9xYRxMQ9oB0y0aH3wIaMyqFwWEVlK2YFYZqNzOtLVH6yS3IIcpUI2es4w
19WbiY7zUjwJpf9ZfxwBwGh9V8IxpZgWht5TJzCLzt5aQBhDZIV8gJE7AeBYJETUJp4+GJJ3QUx/
7fUj3Jg/2B3ppesV+zq0GViU/cfj2L+OrKwqF6C0u/q5EqndBw4KXUqxdy3x9FYqXhMoJymU8VVY
sMqQxniF/L1pRFOBVY3b9TqDDk+b0VESBueJ/1RfyF5tI9uOoNIlyB0koZ+Y2GM5JqY7iE71TQfC
C/90wt5ShjdLuCG/n2K8zNaTGYDvZcHDhHNeVQLCOkIbOn1Jg7uzXaAnLznlHv3zsaUdIsESjS13
QPkGV8w/UPDcVp1CzVnaIVV/CytYEsUg67GgTDYGEQFO530GNvu4sMH9uKVAdzsqgIVTTRHjUDRv
mnRzgJRToJ3L0EwB2anQTvfjZjf5JO17DKuEwfPPwTYs0i4YYMaFcf7Ofg8Ld5WDg0heLA9SScdp
PRlshLa/I7v3/waJiykcPwlXXhfoBn1AbKcfflnrQXI8nkaGcPHQKlX3z9P5SIAf3LsWhBVNfU/4
5GvMu/1Pi3zY0l6n7eb4+3y12JhWdHLrx2kqWtgnD1ICMgK7oijTre1aq6sOiW7eJPrvZMkl6jlL
TuSK1gpYMej/oKhs8Ld2EB8VVSKq3OszZqp43alMdhnC5YTmVsb+HmCkHQCUC9Zwkk0A0V1FVI1o
hvxVucVTYXSnpOYt6Z/YqDaRnrrMYJ2tJlTbrSLlvq5W31zQtrKyI5Z0tILO/mjq6jA9oI2DvXTM
fDnzvrIPlZUfYyN72Z4Cr7PxIUIQAHCIaZUifQ0JfF2uqRs/m3UjVWy9IQxEvv/1VPAXPTmN0CDD
22OECGDgDNputg3nK3z1aPW70F4xJ8k1dUeGM7piiKnbZLjqAtc6fA9p+mDy0HerUVxh1z0JIy8K
K9nOnj0OcWwjU0U3w3jkOh5oNjPV3R+TaWQaGayeitBGzqsHSbI4XAWWyTZSpnMhfJ9oid8C2fRp
9syUksVmTvRcSr94iW3pLXi7DskuFrozvB8hiqLl95LWOLuEWhYXyYiS67ofWe80AyzNYCalUeEh
VZmpzf2Yw+osCr/yFo+fzHUUXydxVbGeIeGbQYHUhrhDl+VrjP6e9WW3t+isGsdNrFcWzP6I0wiy
G5FdVyLsxUIqqfMufaNNXZ+6WQiFxpPMee2jX68TZt9rLdz86Oxz2X+FEY0QXmq4H8Zu5bhlAqgc
hyLqjlXHrJkRueNIO/GPY7esUyAiEMjnxU2hOj6HyguGykrhcxXlVtzGzm7iN17rhr9nIU4o2T46
6ZrsixFFFlzj9hmbqV9HYbNMCOlnqt+m+6dvGd2jo6j0SJcVEgfgfFze8zI+8xMCaLWO3hyhLpyX
b8uq8kTe8yYMp5gswo0Mp4/RwbRrd0XiBFqpq0bisNgQiMfSo65ptQLP3bXAqcmBWQGhb/rF4c8e
HYX01zte3TJGv2jovhBz/Sk7/pqvUw1L0sjZPtoH7PQcZM7V4+unw4OOaaJGXypwFqMz3T4VJVPM
+LEzKVkaOeqkBnWlNgWUaaYvya76rw84j1AgCPSLx1EID5hcad16HlK/boE+vPqd03ynRc9ciUN+
QPazQkLJFGu6XgwWFVDdfzzXlTMoPSctbfvLiYozrrLQfaXt9CgMW6QnLHGB1S0nEazk/thTpB2P
VrJNF/KvD/ZOvprkZWP4RVvPMc6EegoPizBr5WZuhD3r37b9F4hPK6OiNXZco+hUOh5z4fivcjIe
pDh2Rkn434MY1VUOBG721O4b4OtEv/oLNS+cOXXOUP7H7Hmqiv4m7uqMAENxqfMTqo9FQzRGa/Yn
IMtwBEzs3HRYfJ3F5WyQtp7Sg+5GhJn61E82/0+qOAjfo5bhphjFlBOq5cBNFmMfhw6E17YRbYHU
H4l9QaR2+3hzpYwBINSf0vMBrZAjmC0qOTN28kakZj5Woqn4HL4F8OUegWBrpSSNUyrxteT20B8h
sRI25vwwKRbV7JcbC7saNq043totcF2Ae7nt6E/hmRkyBECiW7k6AakgPpw0VAYqnVOGoiXnp/yY
bstvIX96S+Zw7I7y5+/YWyRDds1aNRYyd1mFGjNW9NVyBJoHQiDaVPtYRdV4tGta2vux9iUdXRyn
Hh/3PvQF/1IuqmOWEwlxrZWmA4p3W2z2Crth9hofiwDAAluVmBEkd7CiifJYXk8TxmRJ3HdtdIrb
cjhbw0AqXk8HpuiRXVDJiee7T847r9eVAULN2vfXi+fswYw6j2duCEGdzX9BwK3J9TcKxFZ5da7f
6WBd8RB6ZzyPWanc5hZCgRuw1iGFR07zOJJJuT4E4CLmYb1Bfv8HExinc4A4tNd9lybGwOP9tml4
vuop0NurFBWikFuyU2T91OjfxlW5yHEqNFXHp+hieOhT+JSAoEiMAFOHJywMy9LaUq5VSIA77dj2
UtqKsFxhX9WK3MQGYQ6EWD5TtvITnd0b+aWPqqz/n64vZh9fnOxUtKAPHoMm3oITrraQWJBcao02
ufNEPGRYiISDWNEGSuqvADrg8GNKk0WzNk+Qi0FVCNVTplXe1db4L0l7fB37yIDGex5gUKJ/lIcQ
4VHF6XCI3QKPIDGfm324bZtzqg6AS+Rel5Nj1y+cW5B6z6tjXlia91IBVA9MQFDrH+5474FaTm8B
VlRMPdZqSSN+flwW6DE26gJhRbNXAxKtTj+G5sENbS7N1SqQT+/rS3RWMYPj/7xvStFlqaPwN4O4
SXdU+9AgKe7VVLOCBVcDvbk/Dh/DeD+gcfJM82s3m90+VGaTwDqt/xITFwVe0Ti3Hk8431HROD+V
pfvqKlMQ/YWrSs7ZaXaj6Vpyy+cQ2w13L5sDgHNtJA5P0Dzk59MQqYkolY8/z9dcU3UGaJJ+04gM
MtRx9X0wtqB41SpgdW5ObsnrNW9n5nU5BB27GrNA6sVh8eP2XjWNCJs5UtNV2uYxNh3tEbOkn1sl
lHO2+Lud63M6xj5FHDVx+d69Uu0Hb7tHVeW9E9sos1DHIEWIa5SGU5z1IIfk1LMUYmkiBY3nSza8
Tzw20DE9A0o0oLyzvGHvtLVyHZuEZ6ClZEChA+9Cod6Xj8Cx6i9FFXpoM+XUJv5DZp5NvNzXOzqH
UH8W8fM5NLsXH6GP2Fk6mt2LZMXCGN/JfgjC1c/RKKhnFsdhLCLgJuPuQ6NG7Pmc77kTos5po7On
Dv6eNIsaLaEoahhhC045+wUxMKF83E3AD+zzs8M7rarONhvJnJ//OYt1ezldKJiXBQVmxdZZ88gE
5+fGucE3P6z2aCK3qqWAlI1zIoO9TWuitKU0OUjWUDHpPgs6eMs/WbRvrW+M8UlbIVE7C3Xr2s+t
noczd3VBu5kcHXNQWtHfrUyzQgu0AuffEwkCTBKSxoPVQiNTheYwOlJh0wOIf3fEgEwHdXG3N4d7
Je8TnyRomlCv0bzX6Y//tHVxTWxE2KWRVIjKEP8LxX89TFyHRsni6X/UCjXaJ+wB9Su7eRkM4UNi
ELwohYyXKZo4Gjlg73QPcz3+aiyV1ljGyxON9mjb0tR6VSuiWNTX11uAARNOqgaue8aoDprTpR4+
9dH42puOvWfr8WDk2vEhmGTW2bTkx7AhsSkehCyNTMPu1unn2lVz4P7bwVXvfgfpB3xwrnxQ+rCk
/KjT0aYxhexWLU0ZAxEXBT3zR8VMqzbN4Ke3B4PC7taYAXfrG4hLJUiFmfWq34RItCGj/CKFsucG
JPa592b0f8zCLF4d1Q8vxGgeHFGh5ni5YXT2GzAL5IiE54dBzpEo2T5dqYEwdfHtU3wp0WORRXCf
3OhTNzI8K0sQeqZr/xDnv6sW1wcUYPk7dIN0N7ekXN8bIh9CIwWOAMgdgzg3Rl8HPkw4Ace2/WqQ
jxjEnef08HMwYijOA18wSkB344B5HKaWhYjjVkpu3vlqtTzwPELXPz3nsnVaJI6+h9glQ2FPNMhr
LJoBQyJFvC+kFEVhMjrVOE2N1bzTxAppdYgWQ5vco7QspT+qHYpbtQDwLrNJaTjt+h+6nehZshOz
NF8+O/1erFjsZcucYCaaQRMkAjOK4t2RYZej4uQePRrWx8QfJhy9I7cg1rz7KKRAv/9RsVczgdiy
MIC2P19rVNX6aPKpr9HvuT4jNqmuyUNGO1/0a5A6WEmBF/JZYu24jOU0Ta2/tbJezfrpLgwf4c4K
6PlJ15mSI1WA4E/VHAjj4zAc8wUOzoBs27NYc4q0pWfaovq3GeXXGaCtrGhHFoi6n2dO5TGV6LTq
bO7qBklM56L3THob3VDy890z5qlt90B3K/0cnPUaMFEfBiq3I4VocXDXgSGYjR1nGGOqGsw2SWrb
MLqcJjr5w+rJEJzHBB/62tChftkuQZR1FqUGMcwDatzfs6HADt1t8b3M4jRYqHNMX/jKBh3wgVHd
ZcIznfm+5zigLmiJJbe+qqlOlEMdajBLJJz+ZpHA3jQmnEyRrpLuDEOAjv6Q2esG82nlZbwnLLAp
cSLodrclouoN9/vIEhH4ebO92CSwhl4tFzM4Uw75DJ9K8JlDZl3y5NgFgT6Q1pKftqgJVlai5GN4
Yl8rN8DvhN567Gv3jD8KT2ZEshhSJgrM4ChOey38eNVBzC6rEmI6P8I6xTNs5y4NcyHZKXpxzeaw
LPz5pfkhhFXCBsjlAEl5af527mMq70ODIN4PiBygbDBQKFPmtFMR9g/YVkDNqOnb1ZWOlip3xGPN
ppcQgXWvKdIyhSZG16V72cPLUkQwqkYOtyV5vccS42vdMVUDzbcMrTCsBZFr5me+PoOSKN9KzQ+0
QB6eA7B0ScNSrM1OkHnhqz5QzJTwZreIdqRCOj/bE7ijqkGZ5bsCsepMWnydfUwv6mrgxzCpKFB4
Eh+EOsDqq9468tycNAQBMCYkvnk62F2ET/c+s1JqhkVHZDlyEvl/MX568RAQEi39SW789KqfJ96K
2QmO9vgVQjqJLIjHuigrjn6jKvxVYBgvLoBIewKRLewgeoOircHJ98KOIPl2zdbJ+5JDsq+aAR+r
3FzbdnfQOD4+NtmphrFyvyYqWlWSN39bGR9phncpgE8U3hPiSyV349oDggUdQHXjwXthgD8BAw4J
QUmFClrEQ1qFEWlC31yaV7u2eMKV+pGnRutPvkK8+fpN2dIvCrze8KcEdvMltWGCDUPwWr4Y6sUq
fFFgQ1w3Ivqs0hnjdf5iYfeiapv7S9Otr6JRV+sdJhMA+UAEF5ntPmqzRJMIscBy16n2xBugl0gB
idwgZ5+XD54QS8PisvB63cX5WnShcBSoGhZLsWGjooaZ32gEEcXhUWw5Mc5ggsHe876Qh5N/V4lr
3InvdM73YTB5Xl5z8kVkkJBdxetjNJwfWxtJ6ddJ7DhDdAqwdSY6euvKhqbPAtKh8NfcRGAZdimD
YO4Hxof9EehqYbAnL8kzV388ywIwvJM6Kn/XV9ebuJvlo6vsLaZkjHe4CMrHE1UYYnQKq38yNXDa
Eq5aBAdPVTv+7tE7/Td4mprmD75utmTdiI9WC0+Q6ymsXDQHSkoGejYIQnoVkccyLD6kE3BFBQA8
HROBBBP5iPZMe7kJTpc3224O1x5oKD33L9JQqC6RraQ+k2d97dlPLNFyb38ENQdXlE42aNQOr8JZ
XaEdvblUVNXw65XtIh9Rmn6Wl9jl+cGlsSCkfZ4cK5C5RqU3jxCy0m2NA/SUdnFZqF3EHrjq9l6N
s9M6jZmXKzFk65xOeMkXNYNMWPW2zNxu70oERpZy+WDBQGNrmIXFxPxQyIHaRF4JHRwuA7JWnqip
AXUAxr/9GKSfIuO6tblo/CkTmD71KalFPo5AE5/3GJKDJ+wun5LfIS/fVYMCG8MjTMxqm7gNEdMF
fdU14mbsZqtrb2iqJnzKyEMA+693rzYcu+5Z+tfLybMq2/D013QFj30t+uXdh4vwKFyt/06M5654
JGx90bPcB1Y7R2vIHP+WUAPvDcqBbaGAMc2rME9mCg/8fGKkLOzr/ZwmCQcxxkL12dWgap5qux0u
bk1HLkjxx/B0n75Z8pBTgV7M42d+JjCGb4b/l8G3Z6mcWdj/urcZ2HsuyuHeXZtrgriV7Dmwx4Fk
3y1NlRrKRhiXA9MvNOsQDs/iDHdjDGo/jfjCM4zpIowHp7afVIqRZmzI5fI58Mn1aYIx3UzClqv2
YatQkHS8ujc+YQpea5mleUK2dcDOPsITx1VdeV7YpTs5NvnhVSNgd7VEpbi7nRjHQY+ZPOLE5H6S
P5JSzCR3Vp4C1YykETTUeIeqJI33EUIlFCavOcBpCTjBkLZLIFgv5hy1i2hrv6F7iYEzOjmLq7KT
uN/jNjQDsEVYSMg1ZaFs60dkri9eySIEN3vaXuVx01ENylI52Ajc54JXRHNHx4B+vtdfTOva2drG
VoSOc6VdBsGJlqmZ5vY3txogS/mnO2e9pI5lAZhk+zOflHkXfo4bKHWUBMFywouEpjlQbf/DfaqH
OLgH/07SfewV/5BEhZaPuT0gz0d5yPCroFYDoUVxm2QxZEr1hPBdJUgs3Dph1iOoNjesg2hsnmDU
bWFuvAdfVU1PyspfQnJWBVUT210rc1X4UFPrzk+/6y4yLdq6NLBzuj6jt8n7xti3NIrUvfogC2AY
uB0OlXAQJXHSLCybhkiUgnaXKWzyYb9D8HQU4WBux1VMsRa6cROw4G7XW3ZbvCQyl84db7655o8n
Vzhfd9Q4wK5TfbMZhQnzII2qT4voLomrO2pxY4V6UFAVVMkD/pcMrS0B9otXUtPD7Gl7AzbqxMYT
wONbWIw9C3vOpaq0lV0i8CDQrfGhs5a96eSyhkoQYrAmL3zlODDsC86tqNnWXwfn+xsrlkOivti3
IbsiRbAm/wVF7QvlqS+QhFRXiWtT8AB56lSJ3cLKHVwZPECDCHtmzKuqGappbRqwj3lF6D/dWjH2
m3+GgUxS7Ru3f5r1GDoKs4LSjxFQaZJfxQHtMhaREMekrIZHhBKlEcDCDlCAdCUjOWakbwBIhFAX
aHueGbQbat1+jyWjr58iEzYZRd3yAuc/ue53Thjz9b5i0b4q1g2frkCJe2Ok+V4jQKAYu2vgDCwQ
K0BXIqWZ2W7ucCJVJ8c0xMb88sdlOkX5JyHrYUb5h/fFpjrn3eeBjVF1TgdhOvDR1Md8vfycXF4k
PXHPa2yJPM8KHlsULXElph6T6jqvJPQvMyOVhkM1mcmCLvr0w7h0w8Bf6UZD1OzwobmbG2JahOWP
JfZEIDwTw0sALlqpltGrnRJWLrjXksrqh/EWo/t9G6+xnIz/7tw/kESwbDn+FR8Pm2h6c3fgROOg
BuPa6FHl3qGOVq0Kar7xyYhz6x1WrKO61FbKCISZFxdcOZGianQRNS8eNTEtDoU/+hMnH74FpfDM
s6iOSNFzSOkPvXVGo4rapg/t1Lp+0ebOCqEi9ZvzwWfHOrkZn3sW9WIOE6mLPrIapkxXSzu02Zm7
pB7Q5MegZSgArnh1TKDPXXk7E4eHtCPaGhxwLcQBxrD2NAeregHpw7qE4k20869qQ6qmg9VZ0pxl
+0p2RcnskFFy+iYggnsA67ovbHmGrHF1Keyh/TnpnCRNCdSyu96KijgAhQVmH7Eke/ZbSZIVEpmE
YGG+2JzZs+s5h0pth8OX9hCPWIqfFGGIr/uJYU/UYX5tR9BAKcQ98wZuFJu1FfgxAu9EL9o9IfJD
+oYrj7Hh7nLUOSlZ7+19Ync6/TMpSnXss1+sB+6hFFOlkemb53GwlHIopzZj6TZw4Xv5hUQgfrai
owZ7w8QMrYzUoFFBl/2CMhcZCWLiT4c01fqliPcSfepU8KdNr5+0QZfxfh7Z57U6TDbxYJD36Pdd
331LxG2L88kwoR4zZCiKAB9wkxBHhrNuYLlHeNYWQm7+qLIF0cGoghhP3u6Z6MYptDWAkb7sFywS
ILHfxrsG8nlJtaT46/LHY0S1N9TNbzfUqZEDqKwooXq2Vcog/LFmr71Z8vsNeuw7iYfY1QYnK7Hw
N42w84NmLV1KeOPKVovs4orxKwvfK7RhMgs03Mbv3UcL9QtGRGMUGBKC+aUs3HAmNOqLeUH9JPN6
CSzA5BZ5NRcLWcd7byMIM9xtBcWKv8owqryQymG5tRLY8j6AfoC5bIB9bmWKIoNKNICibb9SIs3D
pJC0yYt4QtDUYT+C5SFY4+wyFLz/y5AbmbqxVIAlPtqKJxqcqHHRIiF6tZlkZ+2Q6C8mIG2iP5od
7mHuBZY5sLn6tpn9/j3NheVnuqH618aT2K/uDN2COYVz64365jjTyKFoukp5yyxyWLL1ZYB/v6TT
TskMwSgMYuLkd9exSI/Q4ufSVcHnRFcQObIsMofjKviGAP3TZ3HpRyl1n1it+btBsFH9zRh+gQiz
Nl4jMAt6hHBM3s4pxeURG4rErEYrnBzG7AxnMMuc+rIOug0Y+e4j4u0WO//c7g7Abgh3imgn3QVu
O0uPcDRN1RCsIdNDnj76QCnC2/MNj7Wne8t6Ow1ZJmMJzJCRQq72OHDbLFKPaX0VgaPZyN2TIxhA
OpU+3PTUzCm5B0AOF/CDeyISM2eg+YqiWil1NaCsF0XJnqvEoynVdZpCasv7lBlMQz4M6ba+H2Lu
WKNwgiXco4ou84B5TQhpGqgPKgaiCbUGHgqcdEzcMKxMRtgv2DjTILVsQBPICYut+i4rG//8hRma
AoKXeDBzOC8RROPeBheUbk6ZDXdWEcsCDyu3ES4xd74RyRYYhmosgQRPbVMI4GoRARCpHCUymki1
JCtvL61Y+gP8S5RAzXAUS/PR1ESK1iasDVFEguu13AGEnddTpTKU7laeI9kPgjYZpkjJdJuRObg4
bPrJjy1WoKlbUTcMSnoiSvaJM+2/1WdmxSkZppy2ho+5Ule4Yuumd98OHPwZmZ+geg+04H8r6bhn
TWYCANwrVFwN0ckckHquXbdYzANsyLmwcBEZ8j0jLCVxkdh1465ox+sLMovR/eq6AbUTmVTRQSX6
yOq0Qyb4fPaU3sr9U0AblVSBNBGXuoKjMz/EnrHYByCYRv0zHFfQL1JcAN5AlkfQPu+QAr3DcqHc
IofoLKg85wfHSQRnh1IWjt1lmQJ/kcUvynseAZzwRn6ZzZ/A1E3OqJ1C2mDRrbyghH+fFASD81ya
lG/zxlzS1emK7a+EryqtytGBLA6IDLUkCIM8QkyQo/NN9qYVFrnIaS2MyOrDHxgyaNDMzouFK9JI
j/NJyAZHr8ZLyrRMNgE3tvnTJ4zhKq4Ocd2mXGUC3sjSdnJfKEROrffrxnvtcgWqfqFRzcTnky9O
sgRHhowA6I0Ng0crjDniTAq5LhC183tzGvb6Gdn2F7jzYb6PAg6pm66Vzozb/Jk2OleeBa5hRIGx
mdzI0vkC1714n056hm0LRSuvnEuNCU1wc+507amusWV77QHbLLw1Nyig8MbfccdjWO2kJCLkHP5w
x78six/9hF32/C5jBh6qxFBOG1yO6x8CP66vbAutchZplm9vuf3MLlCzylYWtSb3mC09q/9/cyRa
MgVSJdB1OLSdqRaCl3p3nz/V6xxhGk3W/16wEM/ohxFporNF6PlwtCMOONP6WYHS20P+vOUXZVAK
pmWB57f4ogIN7biQzqFAsFWUXKwM+daOTu+pBmWoe/L40ukDhet4pQ5QR5zyk6P3352AAdWpZGML
i6+1keDE4P5GNM7vw3r5eTOaG3hxpvwQt2wl/GFaVZHblirgcE9AMSw0LL36Jy++drhwvEOSe89F
pEOVkx/DPM9rsdiPmL4T8qvl8p8AK5VZMB6DqO1zk/FTsUMTKVN9+hL22UyBfyFIaRStb1PLTBLH
H+nJxczp/Cjk37MzzslTwiJbI0EjpdELzTby6UL4YOIfhd2Vc31I+mk3F6T6yLJeY3WGZl3CPIxL
PdCrZ8iLQ/jmrL4sq/uREHrR1LB1leMwSpBOg1asHoXtcNGm/QGQJS6EPLosxtN5Qcp1lf/tqw4z
PdPrYeifwuSwcKng2hqBJDji3jxGTyvGLFtMaDxcpow/AC6n3Pqfm9UtHvUOBa8coIfSFKCqWDYJ
ZmxvB0He37/vwYpmgm5uSujIKvv7a6WG/fHGRViA2z7yqSXb+/8y/INq1QJuwd+NBs3TEeU4YNkw
vzg0JNKUVgxloEFpSDqA4e8lhl2hNoHBavpnDztZhvdBb0wVRQ9IAAF1HKNes6KzA/EzGRMORHlv
tmv1L7NdZMfPvV4zDgosqSUyfYIV/G2KUXfHi6JatpAE5byuPmrGRsish13v+nEqLqwAZk8WRE1D
955Hju+02o1GQIX64sOlwnPzh60pZivYFLNEGOhbmsLA/930+jflcoy8fqAsjHPfjB80RFH+R4Al
t3BiOJbXfWZZ86s4ADRqVCs/eWqg3+R1ogmDs2T3rE7jr8M9NttlEY/fy2epYOJyPPJlv7fsSWih
B1WdjHPd0mm0nPervdLs2AnslkR/SoMMWqnyGtDz3YEW04eUMcEOHHwnhRyohzcboxSpDpKME3zQ
azWBHK+PjjtneS3DeaVlHHt4nsHu+Ci4UYsWEdbZ6GXM8ksyMOIHgtXWWfuxMIfDnq6vtjmjv1ox
a2bzXAAQGZtvifxnRwiIQoyToiXRKCdcQGUDivuqX+ZOXiwbMzwcKDnLfgyCXrXW7LVz54pqQWY9
zh33g+5NxRtfNY+3j/ZLQCJVfi1GEWGwRO3r5o2HBBJykKvf88u02Zr5zkkwt9OZ1/29rn6win97
DrUaCwWXyYRjUzkP0Zk6bh3mhndiN4Qpvt1lvB2B8z+0Kog4TNRZdiOZJdZHzxMcoHhJo/Q/Jodi
i2QzJuHTq/rSKkw5/YUoEE5YJ+6a5HpGnQaTX1YggCDNzk4ief3LviXEF7+WJgSbewNQ1xuJbE87
EDMZhTq2wnB6A4ACGn/zIV9+nAFmIq2ZFZIiAQvkpS2xtb8Q+chjWtDw66OPQUjZaC62LBgXBTJC
hGnCWexB0ee9muVXtntfuyD2qxLs6DTNp0BHi3Mh6dHUH2lt9iAMsL0FXoyZqVdev5+lKuIxKkgz
QCgDHvgwAHNI1xAheCxIFTjNN2FsjX4jk7i6YyZO6U8T+0smyGCPs3WlCgAKqe4LZMyuuC/0Jk+C
yy/ahkGQ/Jwwbb166XW1AXCe9cg2f4S94JP2PcLNijDTJ8mAO6Rb7m+gkP4zn/+69c+GITd4Fpq1
+qmdAIelzccdzaDQvIWQsjnUMiynjr0v393vhG0ivvf/l4VJoWPKtVn0E9HFJzgJVn3J8dv4FQwe
OrWV60+5svXasg5wpXRvEsFx2z67p6LqqXI6wfxke2RO/1u2R/X42HqwYa6X4u9iNNT1r1hAOfyk
HhQkD0GWtUaQ0UQVAZ65Ug3b6Wnhfld/yfCo+XNJdWPBt92tXx0Cd5VL9FZNOAsC2x6Zh8gpEyxH
HOkIeF7ehpORpeG7aA70zdQRfNATZnST9a6u+NqUMsL5iInY8zxA4cjdlcA7Daujr5cuUOEeg1gi
2DxJT1tMTlWxBnzjo3Z2p6bFscwWVyWd1A6dl7aOB4gcD4uBZs8dabW0fFmPCOzKh0pfgkb0RgJj
rSP77BYC+zDoisV86r9jz0Q9kE5l8RKvIcc9XnArjZfQ8j6V4NfB7MfqmiGNvHd0xeWaatMFzxOp
U24mjeVfMsGux4H17JqZ33sn0gUc/mY9LnIi4l2tnFc8tAlyTfFQJuZIS9TsP+GpZv5sMk0TtFWZ
PWOe1sZYh2lyx+OGbnGLrkvEmkCnk3BbvoQK1gsf+qq3t0rylai9J3zy1z55CgkLPxjjSpLt2tJw
ATUbCFRzLIEIOMR3v20EJQseDxPyiG+2uqT8bJ0CC9nsMVuij02awRNEdOrGOh/eYuBJhoyZHT22
CxsS35/vvE5OhK3MUzVNlzmh2YQVSFO8wdbXMACWGW/EscY76d7QbZ4/NU0pm/IIQiQoN1geNcD3
mCEqKsulRxW+e9UAzmFBnW5eCg6iPxVtgzFQhfw3Ws6x1J9fA31UK91IEtXXVXwfPt210+f6YkXL
403fhzbq9ZlbCN08TNOyHhVIw1bxQGB7EL4zLaKAM6yd4en1jrMw61U4AamcBX4SPEYL0EiM8gfq
9UreEY7kYOBySFy9tgnRdIXzOkH4d9Ex3oT3MSepCfxRjdS8bHBa4NqamKEwj7pHIvm+alvTEh/a
Y8DJ6iNZQ/2avbzcfjE99GjqjQlavzN0XKgT7EKLhWhktd2RQb/c2/gcLIhJFPLp9P5tunkDLh+P
N5vsjp406TGBId/kmlgGT6ufJutnU0zhyWRHQx3UF8yDABiH4GzGb640JhPKAo9+7Qq5slCvUKHQ
BQMc0zAW85qG3ladCVWH1HM3GhR8KRZqZy285DrGCCVtvJkAczj7OMWDbbyCYI+iEhzJ7TDO9XZk
0pZWTpvaNxupb4E73jM+aMvUHfEw50cQi9u3QvOIoOp25aT/QFoI+6U17VYaImBPr32xOG+uMcHa
13cjlO1mQZ9vsFhgh+ML8UBEB+oxngTlZl2FkBHDdgZ/0WPOaQYZMvC2oBDfaroOPXY9bK8Quvtp
sSgMpxr556X7vP8dSKoJkOH1hLDHCTFSKITk22N40g4/+bhsYAIdsbWgC4+MtkpKDNdCfNID1lsj
LL3LS23RzvK/UXBUoBJ/mGrFqMBQwPccLRaQZx6oQHr6U3hm/DSxRqClrMmC3k7h0ZhYGekDWAuF
eJ+jLwWKaJ/cy+zsORFBqRvtqZ8POUI8aiby0N0hdfenza2illOud8CLie+ejwg/UavOtxithtRv
dz95wKgrQd7s6q2d2gP8SP7btTDAHDCM4Msd42oK+EAKAKfgvgjOMnnXYOPChKtHPLhvO8ShjLAC
rCapHY9pCAIQFchoCIaGErYLBovcDj4V2ZryZAMlo3huy1WQvCSM5itgSHyps3sl9hmDdnYoD5oM
5BzTuycdycskP5pgezJuxQv5orAJPHQwmrQTX+z2re66rSVnp+xQ4x5Q8BIQS+JE7bh5AEgGNyXj
taJphT+UnTqsLBrfos1UvsLyxsHRIlwBUfFCDq/6fBeFR4+PA3PSUodgP01s0ZZl5RCcmwfQBt4C
yz+b827OAof72XUv3QuCWWcF1RnXg332Ok+RcGqJsKFEmebqOnTF2QA2jHT83KKCpQlF5oPxBA+Y
9RRNzzo54IUMMWvCiO1Ya2mh9L1/OdL1LbPvJD/FcbaewHOYqr0bRA1ku2Qe6aN9+7TmW3GaA5CL
dF9vhEc7B/rgO9Jb7wjJZ+KAT+L+9ca8giXMC5VkumEDcx6KcyvlFgKxgecRx0TwR+1InUjKBtr7
5RyUEFrD4nKUabYBmcSsCCBNCI3sKKIl1bmtEsdhX1Om1spPcKOmZQpeujacPlg/n5H2qztQmsT+
MuTlQMs+c+etrpaSg+dDSp1u1Er0fff1Xm/FQEVnY9SrmP3/odJB2HacZdo66iCizCIAL8AjIf14
nWtfPdkvTAlbsnzX8R9z8fK3r+tREUO7qb4uVe1V/bsYstNnU3D39LQU2g/uz35OtnoT+raBoDz/
UTQYSsqQEduW83B4Hk49APQE0NMtvxGjzXAo2f8tfymHZGYk5I8/LqwdpGzNWQ0JTG6nYIcLciQ1
dAnMYhNUaaFgl18mJ6LGdpArhZtRLLJJOuThpqrXhlvt0QeAVd5v8TqDHThB/2P4DHS2mc9rFReJ
iVxm1FJB8gbPTgSqcpIY0ainow+kpBIPudLNpIfuNM4SK2M8G3sk1arzM/TuCPDxU4T4IX9ZWfgt
gU76NTvQCt+Ho2S0SSNBnGJLZnogvSCrwnQPp2Z2mW/piKrXYmWELoLr80RR+XBg52qawELLiB8p
zv5PzmliSfPzxfN13xyR1e8zQOnMknjW+OM6RfsoWE916PC633vPJDlUW4OCSpeZzMFaeR5VTuOs
HTjYlT8DLMlFcJYw1p+Et23imVadDCiHFcK/pifPUlm95RfOSEuOQSGmsM85+a3pyHku5ufhC9r+
o+hVa+qMJBPxRDtlBbTr2Ta7X7d2SdgoKSAlWf0ET59l735vwceUiiRrzHtqk+SNJvcWKcvQ+ong
GAXG54UM6Q249oMv27PUVicWFoMHykKaRLK8mBysrewsr6MskGkueHWayJSmcauLuf+bVeMXCOGG
ggoNqx64AAsqNP0SwFeHx9hYFo5fNxWC9oCW9YsNvwVmvZt7vtgXLs1DSTu8wlp1EjA9/TzTdlLw
WbpnP4UVRrPFTQzZ6qxRU+NC4a9U/kX/vfTfFGEOYmpWpRfoZabD8bng3xTy5psmQeY6PQmThhhY
QAPkLvuTGHdV0Dr2MulTc+93wxW5f0eK8se1uh9PjmaFxEf+9lAqc0tlGdPLcx4g5pFGnTM21s0s
dBcZQ3uGRzzQAn2xBI+6d3BXgjvgWnllcJbahOWfyGrspNjna6bcj0q6ebjQVcTMNCXASQC8j6KS
BgO7wTGoEWcdWEWpgm+bKdlr1gVyn//ljwF+lvr1KdAx+vX7dNfANXXhKwuxvvd8xyBs7fXF15Bx
snll+D7HDVvPq55dc4F421T/1oisZL/pOmGJNdwDLfDLmzptFhkEa2Cne+wQmr2DG4AaPQLzPBeH
+V6m3hqiZH164O6nfZ1uL+V2VTY19S05sk5nCQ0/adQJvH4n5bID2XFwRfVKwS33y3BqgyepAjtK
RIDG4d2OAFz1T78m+s71YDKgWB9ikclsMXrTEK7DhJja6r0XC0LAu+QYn7QWwdK0/Y59l+gue52m
SH8JExZbitQHEnnuKwDtJvlXMr4aoeRnGjQFlhHmkagGtYCA/MyHHS8j6T63LAcU1E9sA+ITPGGg
kVSPgEwOlklxm8pLRaGPS74w9AS3lDjIdYsOB6REIdX2hpXKAJ7/2148S2rhB2pildPbgMnws7PQ
a8B6JLd0n2SEISPZFVzcgGq7wmBwfHMY+Y3ShDJN83HQOqOKRJ2MrRlZH6br3+OfPGASzsJL3860
J+A9HnwkKZvVN4c0hoFUvK/f3s3O6/MGol4j1BukHrixy8nfBVVwPURr6DijpYq0wVzf5Bs6MtGv
EMHZwLsTfRySBLY2n+fqUkt1u4+DtrpBnKl/27jLPRh03kdeQ0NSHZxsrau+Lr73zaaH3vi2uHAC
tFV0axXU1guUUPq8Dj3pkRF9EVkAbgGhxlaARdm2uZ1V4AElyNlCyRmxjUte3HkVP7+mG35i3LFb
wwunJQxR0tpT0s1XYDmR3xT5g/PzhhNGURlxPb3QB7JsXjiG18PB/F/M/MYHHSZm9TGECzarI24z
Z8ZPN2c0l5ilev4ZZxm0YHg7Ml1Nxdr2QVgNwhP7/7bleJ3qgxq8D1S9zBY6XZsOXIRDNidQ7XDN
KCDCbi5jncJDkFpupe2J0ZqXlmE43YfLWcNtIs2pm09hZxplrU82p7Wv41eTTNraDkL39esF252E
6NMEzpqEviLA9ZYic/4nXebiRk1QZwoMZrv1/xvE6929nIl84OUN/nF9vCe9cKXLPWbHTke/6sql
2MgHV7Nth+9eZEIKzkCakWwRgERbO57GsCWvfxV167Hn8mAzZHbJhJZ1o8Dv+uGWP6WF7JnAcGBB
+IxMig/d8PBcZl2/J/DnRAVSmVb/HTY9H5Rz8l6GEJzhhrY89z5I7vCJQAewp7ws0wRI4+iGOGT9
48bnw8DigL7wJeq5fQwEZ4aUV2YCULyTRB5NX5FbcDYSjyuZ/YTGZiskfNgq8H4NySFJtsRBhLhN
tXtkV/c+W1hb69bmc5lLqfuqOFqM3voTl+GhP9WNML6BL3cYLemy3m6MkH5uBFGkbLuw5qhRivOX
pHqBsmUibSWhEBdsptHEcKpV3vkH+4qO0IHApw3X9SJQgJ1xcBGfB+7y8v7NJD8Yc6J0m4bUiIyU
pmaWK+xJq495nAiRk1nl4Fv6iq9HSNr1Z9sRj6ZN+2YkkqtrVmK/oxwEF/1yMF6kZYdAZUn8gHcO
uYqF7Zgvsb6UoGzsH25LBfKOocs55sIFb1LrvJZZlVn9tkLC9bzxHoqjg45s2C5Ysc533PmLunIY
wN/B6kux60qAewduV4L+thKUhFp8qqWrGcQ2N/wk5EHRVSmFq+AV8LegbtBWst9M7dq4eFYASlbm
CIW9idPxqZQevyQU1FXdnWDrcKTfmXvYuzV6StgGUbUOEdiY72HYyr3zo/WIX2iDC+YB7Bx7YyLa
U6ndzfmsaUVAcXkfYPMJhRZ9T992/Guz36lqaVycg9j3V3fnPM3eotxt8Vulyl3bY5nS84p0zBXq
/M/e+IMfy3u8wJeAwz6AO3cpegKeC71aoMAHn6Gv50sBJoYgghhMmG8RW3pBQvUXFdno07FXhq6U
iR5SgO9jKHsRnx3XAfzRAmuDoM+kiDV/Lu4DMwyeAQI17VzP9RDqGEz6N96CrA/3M0eNRco6lSpU
CcvAohVT4JmhWFKsFO7WiKT5AhlOjPWGXyFrN7qQUQYef9uEnFM9xekHmZ4dRNxlEfzjbkXnzUEg
JE2scnW7tpumFMEVdNRxK8Mqpk0kBzB91Ocr0Fp2gBHyUeYC8SDwqHls80tLyseszOqPnBA8y1HT
2zTYhUxa50FLDhdcXMMskurj27B4NHv4pIuO3orMRjYHVgFefRL5U7qmZQ4vCphUqF84b17qIPco
7qDCU65X0CixYxmTsZ8qj5m0B6dXc0EJ19MjfOICiOI3VAGuhWsvohbnutLnw1EXFo8Du0wIEKXI
diOjGfI6PpSuYRPurVzMhGrFiEUoPiXL2nWuQ0Pi6ZxSqf0/mNsukqLoY3aoMBPRDuv7uZD8lbMA
NRL8/Onu/OJiibGqJ91vMdSS5lYpDuO4gLI5dBWH1y2tcux0lF3aYk1gumVKPgJaljix5yCp2lEb
EFQa2Q+zesgYbKWwjMxQrV4YDar0Vs0WWuEff4/YTNq/9TjzWnkNe8E42S/llXW9bx/rwj9ZfGey
q4i3QlAv7T7QBqoYtZQnPCjRDQO5Uhy/hOtBCz2pNeWR2f4oZRdJr9n9gg59aPbJLceX0X6jqm6K
jnoltc/S2N/7dVaXdnJjYy6yLFZkVA3kZbLN5DUfJln2TGjcOrTt99JFiMDoE6pPKWPw8SNtddAM
VUXJv0/jFTw5s3wY0ZaD20QBJdTcnsLuevQKUF8XVOAx7fp5al5RBiRsHkNw2Pzi2/Ltg+uM2SXT
/HPhX7YTKSm3JCJbFQxu32iLt8C8KvbKR92HrVlLb6z8qMZBBZ+yxp4Stu99l4qyb+/FQoW6+pbb
wG82IcgLCtnwMMca9G8jUf0IayunE6yxQSKZhlYiu9wcHzBhyfWDSSxAUGQsMLcQ6m7b4BJpX8i+
15pKQ1ltG1/JO5Oh3i81S+xtevfLUnY/SKlGFp/t3ZkziZ+mgweRRLVsScsS7+YF8CLUw6FJoNUy
siTaFhz5k3/kcwJQ//i5ah1lip/nTAgPdrNiq4Gro5d/KUCrwPvW5RCSRN4ChbssXsmyeWTl54Y8
8xCcYAjU552GZgh6bQyjXP1dSWDJNqjPkUc3iTPuFPDIlWQ5CZjasJFu/NXHiNbcFFzlbeCcF/xy
83k/toj2QH5lvjsKZ+bjd3ppk8xwTxXLJfSb5xlH2AoGoELPBtI4xNwNIihVtYJ9KDdciSBvV0RF
dnd9HEALnF84vlib7AR2w+/NBwG5iS6ZrDeP3bpFfogy0vR2RDOecH7+hvBZ/mHoO4i0k4u3E4FH
rCLUNMqf2ZkqkbvW7OCXDgBqXpcKHnoUOErpeSKGRSYCDPBeXQIWoGPCa2boKgpurdrf7cT9fbog
vMqz4SYXifT7l0879qbdMVysIY2PoHRyYHEAl+HAToVG1uzP11xhbZQJT7o/qjWg3ewEVtGAs7yp
Q2SIzcVautMBpI9E4TOgqmWsYahpXYQWxPSCrY3PZlAdQKjZaLiz5EfHH575m85jeCkqPy6hB3ZC
gGLNTuycFqkyNJvrCZfeyrixADvs2TOhUDRyOBzUazFyrqdD9UxKMwua7HQfqCTGdqA4/tgqv//V
I9L7JU9iLPp8CEJPno4rfCpOrP5vMSfj5ZyDnNzG07wcTVAJwm4d+R8axkCzzJKqilQd5pSGHpiS
2e4hZxAcH/3UtsioQe44PgQA9tUtNdbLUaIual1BDb1aFyamSyZuoCPNJpZhUiFvWoM0AwDbgprh
OB+NSDcvAOQ+lxyQ97eHRWmpp0H+4aeHRvzAw/GBLRAbhoZCnwLGfFSfHy6ZNcwGnxSFRhBAM78M
ZKe2mfWKCWPVHGIuuPwcPep4hSZHaf9hoaUev2bWhGurAAFG9yYucxQFRxMgisnLhkKk9nk4+j4w
uw1lXAxJjXSD0X1o2CXyKHLH05sdye8kyRyQfaje2/UOyEO8z2wF/o/utWDgtQ7AMPy3MaJVhAjU
AiAoD1kyCqFmbCGrt56FRNpPS3+yxxTRvn3CrBD6hH51A1NJSAixCyx739Ii1G0P3aNWa6VhsxiT
KKhOtWxbOYxWa2YZ36rMCecNYRUxOjmMvvYqY676+mJzyGnCG9CYYIcdEWxRvSeeEg1GudOIUHUe
Kfa76qyG5WvrY8vGWhaxG/Hx4Ab1hiGyxTB+JN4RQGQ8JnNs1+pRQEnDZ/XMY5NbdIDOr5NOxG4j
5WTNdizCiA6iiLAMsTJs87wMNC+rhHnf1y6a9T9+oZFFpRrFqKjJVhCNUKm6JM6LoL6CnTNpQCej
6TL2bsDSHOb6R+KYT3ZbcZ4c0XQ+OmZTvuGjojXaYGY+Q9IICyctG+zPOSrzrLke6JSpZqnnvx6U
398m0gU4G1N8EJqS/B/+N1U4+teMW3p9bLhDtPJHRqY8zfN6ZaWIxJJ/MjAY1q35S2eDb2SS1h7o
uiYTM+lwiz8zFfuYpkb1Cw/+bx6dGcNjykds1gxCgEfzMutYcvfsdQl1E2pgec65ueAJVKo6DaOX
YNzWZwM/U+b7c4fiY6/jM0AwZ3O49LoDoYQTx32B5ZK59RuKDT+JWVReS2hHmFxHpAuQAHeWc42/
8LyfdqXUwhSbmqzHdZ3Q3j8mhmPauZJBlNDzwCj8UbOrYY5BMd733knac12zSF4V5zCbGdFN9uaC
vIH5jRbyrMLhqKQhPZKmusnJpTI5YaIIJbH50iXolm/g0tRqrVQ6aG1MZ+mNZ5KtxJvXmqVYvyoV
cXPXCJDFm+MSyPObbdm6byz5dCCAKHH9+KFKRd36gROsC8aOP19XDsLx5inKDrGyp1MKsWJkeZXr
xBAXH7u78juhfFGoEMnfem2JrRQ4cKVJqJVeifM2nAQc/ATWusScI5jtrSWHO9aKqAURsfKQ3Zoy
o9/qUxE6JqPYWhREOrx+nWVmaRcYC/qxQySJKdVrTKkMCqPb722MkJQvF/C/goZB4grSKZRQaBqU
Jv0hsf7QYXdfMeLrwbDd/9qIQHxVUZ9KjPOqSqg0ih9PbHUexD6JehgF98Gt6adCrnDHg6pKk9wB
HcpkkaFEglutDG7J3mTe8/Iba6hbnkXJmbsluwoMvrKEAT6sHZOXrNJCAeefUcpEev+TNXdJ9XAh
HfYwfVldMmPOnw7h+S5JD4Cr4Q73wBSlr7MaRBb0MPl/540DU7YYjqLJ1UpiFXPHBJK/nlRkmLz7
oM1tYBjIDh7Dvby3mVhQOngTcp91sJfLLmaWNxrF5iGUO/KEvj2z7ZjmvVyqKOhrQkRKztbVep7h
UkByitfmgqhJ6xPvvQENoCDmzEcY5v07NkMslSsdwtXPTvC11vK0wcGdi4pTyqSGdlxIzaY447nt
hhpFReKoNtBIfo1rMiF97jGvJCi5o6ACi+x+z4i+S3oZY8Em9gMMxAjCp+L0L6Eo11RFIADOl6mZ
YHICaCpPJ8ulYMVCoaO40SSUblKOwbCIVq9tmKuaQjVUEOejN4VNIBpNxXXuV7WO3cWy+751bt2r
NtpTsyhuWZgH1YxZM10vuYBN/snjMhy/dnc7+K5CGbFGafokfzUb5c1ZRNmdeeQopDWfPlhASf8P
cu1rOFKEP59BWmG36VELgUvnWRFfXc1474TjAUNHWpteW7WzLmTjIbKb0UXbP3S2sR5Tfx2/3EAO
/TXqL3Dp4hFTtkNCleSkYdUPADW2cFzDQD2KhQIZM9NzBQT7yEUdh9kmVtu+NCq/D+NZ9wOBDQJ+
sULa5l+My4KATi5r/abA8/+BxzEJx/o1f2a5RZiQM7XdV5FSzyHlXCQzFBLQLYSgi+jcCOEJg9pQ
8zav+9fkNoX/AceLFO/vITYe8IVOiXXjEhZs01qvO/4TdF36fulG7lYy+hav/xSX89tiNtwgOICF
aL7hUuma7uP4u88CF7HSCe9xl0qWO1MJNMnxMRpL+Uz0/M5d3IPrGeqFb6+Im46bBO6W69MrI8mt
qeXcdDH+GSpsxmpWg3yu5oMJFsl0HFkQp/8PSb0kial9jKAy7LwNPVGyvaSc/sXfZoEf93FeqIqK
Y2rRl9KburmA3mBnEyiwca4epQ7sCmekoKDlDHorIEZ3YWyGrMoyMyM+YQwSAPbAquidBYNYpFE+
CRIH+sYa9Jm2k3KcsBuS7mqFHlMRpiYJAsTqRV+6Ng6n9LUSIvebmpP+3PcOkOjFy9/pZsVC+aWi
L1Abp7S2MC67gjxlbwjoal7RUuJUckQxguUXRHXN10WliyOn2xAJ3d4ym9+mvmha1XYeyiAY2RrC
siDYT+98rly3Lwbf3BRpj2hTwzQh71eCb9wiTxZYPEaX4YMP4kymUDb5o82gdCA05gbb7AgMH64B
/PBSnoNwcQjiFTaG9U/AN/z3NE2SYIKukZ56WZ8ZrmFmwJSk9TrTAoRm5t7eemOLSMWkRC5OwEFK
gSZkoPuLBuCAUH0kWgec6EL6nrLEWEKj0/q1nYTVCQRs6glvn9sq7DJaKim0rRwfAc2VCX5jDvE3
AsewPPTKxP8tIcPj1oVdytZuhNgsF63GhsYz1w7FTTrlOQAKQwlu/5v714Iz9YRLo5Zr0JBr6aAH
EQZMBWXDPL6AeTlGmWID2Ffv0J2yz/5sB1fu9roZP+PT0yl2kMS+QV1wpa8XsSYr7RrHn7/3BE4P
KuAep40migblmNeYke/q+YOOBCGoMTGhHVXzjff5w2vVctxqp16ZhH6juY6PDZlB2DFb2jsPu8j/
gGsgsBtD/gyprxNFic+UZZU05/LICsUQ7UcWECJR2sgAYp1lfSQ1W6W96dTRKA4G3MpTPGXR3r0E
G5PM9KZkkM8LyCO2faWAMnTdrfJV+dE85bkOVRKA+tnl391cc03WdXKPUqnfe5UsgNV8AFj7pjF6
oGnVieD+LHxkg6XH938G1CyZNbHpmT9yEZFq5YD2dbEFPzRSAeHij141u5iFYrISS0AMIgdWMIEG
vjE2/m5RT7GaiW1Vkfyi1fECsov21rYEWH5+ZkBUcR8dXn4ktojnKNSsg2Ca2OfiTYt44r6gBxn9
l3VWMbOZGrOrMy1wisrIP2nClJqd/eXrqus1QdwV+p0jzSi0/QyMdihMloluzuGmQu9XHnrMAfLb
1GCl+G3zL+OQCWaFJSvtJDNE/W0M8SAZ96jrMUVYjBC5yS1SGGdqPUzyI5JoE5u9hQZQHredvunk
cZC+glneCUUwKzxJARG6NBti70HZe2SnkAmoKwTyyfbClew7ZxXygTfczeBxyCTvixyupRimejia
wScp1BeMgkbeddUK1BCjD+bL7vi9ETRSN4ZRMgR/DIxqXpq/jziMVT2/uzd7aegxlvfX9XrI7gLd
gjlz6j+mLGfNZ5LUqwwI3TUKhzABK6M/1Qaws4OCdQ8O7Fhq37VBkRStt45Ek149ZlDUfBRsfdlz
wK+Z18mQ7Z6CwaoCDS8ppZO9qAcgO3uNSR4pN/1jJ6M0chzx1d9PkuS9H02b+QIZvfwTivipXRG+
5N945BjrW25xHNa8R7+Vw82RBsZJV/ymtHR9O1Vsg+SJSYXdafsUP/unsKRdd0nsbkUsYHiQ8xT/
F2UG7S2duvQOlAz7GZRbq+DvLZHCs2oU8SWQ03SNwmOQ1EcbmBRjLLjkYd8/tuApk5nN0m6uzShh
j/NcjzWmxPO1deKrul+T5rlO1/OZUQKk7Zl1VC/2AJzf5PkPlHhhaARNewjpFOu6sMzkfOasXmTZ
ajs2cSjWYJXDxs4kGAXYg9MsfXIiJSl/TS1swQuL6Mcr7/M8H0S/1l04Dfi9KN7HptlSrphgHUWZ
Cd927N0UiOzZnCcvX8Tgs6gSjmN/wr9tqLvBzOOem77WZ2w+Z+ftvYBURAmu0XNIPoarsR8LXkWr
TptNKABk0/berv2ajEehF5VMPCNOiz9Bh0sLSwIFwBH0BdgJ80lHa4xnkPO4oS5rv3ySnuqKAx8D
3LW/anUHswzclF8l5chW3Wx7Nnr/vQbL9thsKWl7yeleV0BE2COonuhs/AEiwl5Nnun1x6IT6hse
JRnSZk27cIaOBV/h8YaxlZK7fO5bme5KK3ILe42h3p+DiZqCaFKbRKVytiBGwhD1xt0sOXjx1Me+
rlmy545yFTfKXJUZJNBCsTGeDGqEDwRwOARBGTPzpSv3G0vzsE8HrrYrePOPNjbcj7yRFVW9EdvO
Zyuk7Wa9Ge/lF2GH3BEPEVSPl4GO9QyeVT4AotcFQ+89J2P73FeaF20+IeIGvB8B5yQdMYBVsAYD
ooat4ttIFXORgauVePlaGDt40t335LYpdoRuVJqDdmxPvrP03Z2ioWGWkq5u5F/77b8FqOHOcH2y
Q45qwSC8RVY9LCrIuT5QiGOnqxYvrrIW7t1AJ2DqOPZafPQ6rvDTydawuN7MLz2uWJwqH3KkkJND
i9oBPQUOITobHbkWMk5HTJqUY/OlzyloGVsI2SctvArEhtUMKrD/4V3FFG5jfvzO0pxoWgVARRH0
y+SjKS34NaPajzx8l/sebAlo33GWY77ftBxiZmPdmkAzsXGzI3jn7I+Ju4VPuldzkfwnEqEG4+4z
3hb1gYoXV1R3h6jncElGAegYSlObHSDxt/ZvY3/WpU5h5fgSTlzY3TV1FQiWuzm8jxWXhGKEKRbK
bfsX7HaHaAG+fis9Pzfj5Km7UkfdXhK7uiUKvZ1cIDEpwnYp6ivxw+l1fUzgRA/KYS+ARBB75DO1
frJLzseGWT8ucNSoZ5SzJ3G3v+zce0bALQI9T9cs3YDG3KatLJvS0qgIw2mYqrl9iTwoOE+Z0E8l
H6FfM60XjP3/drTQQFk0p71Rn2CJDPdcjDN+Fc44icmff9dUIZxSl1R3pYGd+rmMuAbo//CY4MVL
HRuryZ5/7nLCodv4WdZxYmqI5c+wTktF+8URBGKuuaTg0jqTGb+v9TvT8+9/VuJ5188Y3EzNjUwq
SlzMzkKApiJSwO6YS8ff7AflmVHpLEtEHk9UrukwYl2llnVUjTmmA8ZUwJacxgGvvAu53OxGJQiN
J32ImDL1/RUXGnh9jmBjCKYaomRtVCaY6fFsDABHoiinOnn2TujhAU4+eK1oeELwLUnfhqEMzUCL
8/2+IjcCw74hjMJRJbN8+29/tDsas2hp5RkR1t+rEH34Nilrri19EuYckRDFWoDk33G6svnepNf1
wrKi2oQp0LRS6cMJSxEqFI1cNkm3dSooPBCFNWFbnpmx4f/mKpePE9Kf2Thq2MKZiuDXE9HLMxtl
n3orAq1FpGd+3ItisWKcSvAbgOpOS/EPD2UR50j/aCdG45qINzGCfbm+667NdWHfTcynyn+uUuOM
x252a85yVv8ho2Yi4zL1evDSXz3mVqzqtpxIB4UPw1Pt8cDQ7Nyj3bA3zLTcXwU60rLk/dnf0XP4
HWRdHoDHuKpQOKe7Z5QUHqp3iQg9N+gPpbVDLCDgVvzRCdqubFRVWCw3R84H61hhaGeF/x+n82eD
qjNZgRlfzGAepuwgWiEGmNE11qZ85LPExNqg0WmFhGvTO2hizC89TIoXrJflovvd/L63QVFMI4yL
AA8qdvk7YisgIAuGfqH5pUfRrR2G9MfpXzZHVeH8qEPxZ6v4nm/IMX2Dh5w6IbIcaRiJSqVpzxsi
ozSHaymEnf1hFk2h8FjMdW5WXbRUNS7nfZIoxEN8Nog7eb/XemED9gJDhLPbdhtK4BAe/VVBOUgF
338r8id6QUlgrayJU1nIvzM8TPmvErUv/ipS9ezm6zpK+SRTY1lsk7Z+oQr3+st2ist0FMT9A4nG
OubSVgYJvAS54MVmcQQwcXAGXl1hy0QlID9VyESfAbBDJTCeq/at34+T9WrxTOTK9Bh4SFAdqjVU
UanuO95HurYGqy1G/LdRJCrWIPLo34b1vWg4W7wMV8N2Key4PQeAsR4GZZ1dGqMMJAOj/rQ/YKGS
Amzw0nrlwUfau3/1DedVoCVad7+4eVxCss3YODVxaqumwFAY0+0kGTlY57snJjzQmmVmgRH0i91F
q+wBa/67+0OOBNkwkoxQqBcOLTkKpnFw/nomuqHw/RkI8cjyJn6NP+13c3wn0cVzrwwKYsVa10Hf
RWymQgOv9rLW9V9oNrkmKQktbH2Ji7DHBiGfsiz7RfzVf3wRJaO3fE3IBTCDmnL0nfP2URYBMq6q
/ECc3GC7KQyuP1Wy6f1RDRc2BxSxFE5/N44XfW+9O9mkforoqJULAgt4JI7bPLMNbqgpvHLZGBdY
+SZyx+VkIkM31/q9JBzoGgrxoJd8sq5yL4zSWdFWQvCahtIH2u1+7yi95qBNynEPODxrzAprJOGY
JeclN9DqJoRdYb+5Xf62vcIbrSdPEreT1zh1L0MxBDakeBRmEjAAvpapOpdzmk4QDJT9JfGY8dp3
AyiozZ9eZQJ1FLWJfTqYhAl0T/WiLiNcrzr/WsKzBMzPi3yTP/jcma8Q6kLnf3JkbG2iNOdx1JLX
FyMay3BsPgmajYJsXulX8cGl0ouG5TbHS/Csu/YD/Kze5jBBEwBJxHT23K/WFAI/HrJsGsmU64ed
stinbJyVpqRd0oSwPkKZPp+1x1dImgJJYwoedWP8dBR3jYK2UFQlEbRO5MnLzR5l42uCreXKzmBY
QtDQJML5Itaugm/b6FvQpE7290DeRaxkgVCtWBFW+Ei4oe8luZyvUvtDfdFA/XNQLOL3lJzkCmoe
6y2pHxkWELpVKDYzTJEypncqChlXrIy1KYQAXxvlZC7Jzttr2qo5FQAGH9U3WDOdcKWDpO2IY0sD
dMtJqKPZp+lmJbocbbD2a+RErKPx9ENlvGG6ABJ32K3UwEOeGeQROyvYnfGobCcNohXZWxfS7K5o
I8zJXrTEV6/k0mxBi3Row6HL7kPvb7IGjR+kZhSQ0oIsa5H0FMfxrNnowdBsf7Sk5H5sl448ikeV
n8dSsOYRrKpgkKrBxcjiGW56uFkY+FpIBgHGHN9rwi30zB5pkXklXcg5OPbGSZta0GghtGCzy4Pa
aV2lQMDhVnrIczacTbSw5zmN7GZpWHOB4MQ/UGyL0px/RDJ3088nkpN8RHzSPwBBV0fVMMRNRVZR
+CH8yF+uT99p0Y8pWLIiy+zaJvRfzQrxMu7FwD1FvzNH3/RXNbj1G/JjzIaApAIgAbuVY166lIWV
zKi0qEFR5vgxdI4K6cNkKqJ2u1kyjjnTgUo4SHQizBBo9Ce9ewRM2YPDMiOIqZeAlbw7a9t63Yn9
mVBwrDEM5dZQgIEv5THCdDjxH6kuH6YysBvIaajqrLLLen4Ae8n0KjttqRn6RjaK9FRkjt0Yk0ba
/l79SzOsC8mRIIFIdqI8Nly/yJlFuLziTrbTbanG5atl2Gi7dtD9U+B0hheIHvKmBeTysQZWKs5W
q2neOsjiKfVaQlNQ664jXBg7ClrFoxnhq8HrVHw875Duf5HngNFWAv+h/bk0eYqQt/7LbO4Z8I+R
UudR6L99eV9+rzNL7oDyUhFS/R4tnte0lavDZ2I4/jJuN6G4+aWQGwylBnmnV0jTg9mvNiu9bxtr
4YnApUje5iV3/rr2pxQvsOiQktR7XIRtw5JDBQezfKpPgICzLg6ERowye/l5p7DDTMg53zggNKmT
1Zluj0FIjOVXnJjKsKd36h+3wyC1KOJ40pmWtaQV+AEzax3id6AkUhxm2BJfJwwdJ9PPBxVv+ieu
CntOW4ttSlmq1rWBZnshhG0fLpFzqcB+TjgsymDhNaCgURrSYHGmu1OJCDuU0xev6N/Vx/x+r+vH
Y/gsvlLP6NzCGaoRCnu3UqegwKA2J6BDrzO9hov0+Rm8OidprBAvQv2WfMOq1cMfjbbzyUwTYp3o
sKAJa9HbxRD3RWLl17MNVNPayW3MazmsS5QES5ruFeuH4hK1Qo3ulAuz1pCOzDak5job7HmKkmFh
X+WxoIQmagm1U6Y+3OG/TsUBITFYEEYkOk0tTKn+4093dJ5/cE5gTSDErimbgoYx7hE2kzWAgQ+4
yXm3/B7cPhATMN7C6x5kTfG1vzkSc1mr3Fywm1glatuSX8CMXn/5fb8tbMggLgk1GQ8saRS7GIp7
OwoEgLpZ4N/l2KdasBzTXXZOtV/bb4ssIsONDmXCtP/KBfoH0bQzqEkKd+F84e7TTwb/AH6fNZdp
InIAH58sAv/Z1yoxHNNRZaeZNmBp+ewVEBD2eXB1iWpBj4yKxZrISV2qIiR4XAs7i/tNfR0Cc+OE
AciZ0tFPrbk9CnAhDOX+D4M7HBnburcxXhzHtt89AowCVDuStGR5bJs6ru2Ect6wu24XJ1kui1Wc
1qgyqZ3zgJEsk/AJX1RjzMfhkXqSRHmm234RwBdZNVOBmSDCNwE/NSesWotsZqUODkDdgqk8wC5Q
El3IMHAct/lqseB6WMumrQdsT/2X3D190NDQ4yEN1oT2nImXLmZ0ftjG1kZdT9DVCM3lMS1Fhcj1
Y/vm+linItn0bmkpiiBNRAV+lH/x2PNqYFvEtzNIQ0Hnrb9XITcKLf357mdKuB1Q0IZjHcVgszBb
sJtt9BhLukqXgLAQWmuO9a5zi8mvRKnP/8+VGbrKOXmxq6bTu8S3VuyDnKcqv30UExq0hOQGVi59
gYEbsvh02wefRSj4YqdgzaDWs4sNjBDhO1wZk6RPyNnk5zP0uYyHuKUK52Xc8TXAYTWDBMqCe7d1
0RbCnCGcxcrxOCEnqXqsotnAujXn9fdmqaPS0YuP6BDTmo4bossWSOZMKV1TW6UVt9vPW8VExf1V
q4fW0OpEkBMp+vj49hUJH4KIx7USNx+NvTGVhJvZBA+r+8NDcEc63bX6henST/+fBthhZNaWm0EL
XRZAfjALYATEaeKpOfyzXFUPDKJIn/zPe3uj3QgBAVy4ayCmgbr386JK4VIJ861QUDuMPnii7HJ6
Yf8ZVin0e9OGIcdFRn4anlVw2rV71VYl/yI5rTXOenO88PesLMur3AyuLZ6hPTygLIisp+OGqdaK
szX2df4TX0mIErNBNG9zSM1+cOgnXtcRbR1xeTnSjWp75lk3i4vTmVkYZyXoj8cmfaUvg7oFrSR1
8r1XqQYnINxHr+LLDgkdBPuAR7ys46eWdqXLne9dKu9XxQIxajWeGxBNhMM6JTB1EWACDJqTL+DI
QrKgrUArdH0ujdAR5lj8BPBs62jZNcaKD945HQyRG24DhM+uJe3dd/XXvaYdTt8GFGhWsuDA+kin
xizGntgIKoBSrHgXCZxnk8WgnysQxoucXaRJomIXB2Lxp0ALkYuRBB2c2x0S0F/zDwQqhzayOqTR
Yj6e6R8bry861aOvfDH71B+AW1n2QCTdBrpQ1s3p6/WtDsgaQLZLygsVdEV01x+Q5KOi6xT9gsUL
VEnAcbu5kg4HE21fu2iNLbcDKiNXB0Q2LbX/+jXgptsfsNaynRpPuss6QBHDMs7aV37fLy+7gJqj
fj8nhcjO+CKiXBF3GqGvSETva9xjmAx3MvENunzHvp5uBJUfZAnMPiFWTMVwgF6X8dXhvcMc+l2u
DrPAZLHxlKMoI+5PXVDr47pkn7YYiLC1Uus9R7JcUBBriC8GWNwir1h14mz64LvrKoeNQ/k+PPIA
Xo0Qxn5JEbHz7GLjYAKND29Ji6odWLSuPfuydL/HTftKdr5Uivgt2aftc/hFoeWcIXVjcC8jFS2k
sNyqshOTJC2SV1ORsZvjpIHPzHcpXf3m8Y3aR16E6V/4tt56ataERffHsIoaDq3rYpm+RjQkC3y2
N+hylPAJhcObYYYH1tOPpAe3nJLx9qzwF9TwKxul3u2hZxLxrq8l5qV9Z7h5UJIGyzZQsepXcm16
YARLtv7jcAmvtJSGh2RDNR7PXjCG2mjA/7kYXWqScq6Aj9MnVUMunbKoVXaEGrK4PJ6nfPkByzRO
dLQhi9IF/UU71jfeDORAgbiaZKH2VgsnLfu35AT7BCt3WiKqZ3EtG+/9cxPwIzWlLBMkIUIzeaBT
tGJHqRzvon5aNUHL9dZV9tNwDxAg5aKNtce2WxArD1FZhQfcicjMgXCg2cyCYW1oswmbvG2ZzcFl
D5hAt0Q/x89Ruw0RCHvc5lPUAHOCEF/Cl+pXf9WeZlJMsrMHsnHe2c4idToyUrv1KhYZi1xayDZQ
MBjwJmuZ0vZLU/1zAZHdVmLcya6mHwWh3dSPcfQFvl/3W/i0JObxoOtZIiVjaSb/3rUhCD0k1pe8
Znxj/6OxyhhLz4oGZxYBrjgG0TW4Of44d06SZ3aWtySg6psstRvV5UMrh4ux5mbVD6YEcZ39BbK9
g8URbO9fqLfGRVnBqgQiRULsXMJpvbvIr6DWKFJRFKjZ+Hr1OH8XRWnLEX2hopQARYY6mdTZGB78
d2HMzJuy9TwPQaNTBm5RYTmaiDhgnjCtVw033nGa+ULvHZ8vgyK429WMEJJYO1bSjz8dGgGl34X/
y7EGNg9zpcM2MahHJ0qBcbJigz9lgYo4ljTbnV+cJw+Q78RV92qiWu85YTDgOcj5XHWLPNV8cEtt
x5IH+DWTUeNj6uVuJK10HzPID6h3Ip6ntoEF1EMcXr4cteKAti+pLd6DQvocmsuNDrPgu1UJBr7K
N4L+Cp4RvRwuvUreM8mXAKRv2IkTRaGBfD8H56QBiHg8bw8PP6ejXJsHFIOdD7Ed3OTGR+8cHJd3
HVzECtCYLrCu1Z2fl5QzsWOqVsdIiiH1/jtspctUQp1hXQAf4GaD5n3OF1XItBAsiVGvGee76CAn
NonVHZsZDs3erH0MOxWzfpXOByduD3GAsSbxy5QcnU3cpA4jbxNaGZhP23maR63BvJ1GtKodYjA2
k39rUc56mGt0yNkNWkceqMoO5ukIVL78Cv1u3WUOaRpAD2t/MmZ2LJyATG27KgyclOZYh8tk/Cbm
yiVRPUao7w45H4AyTpARNYHeZQlVRf7KCT0njI62Ok+wp4nhqi4dChjrfsrrObv96MO/mwgZ+s9b
Wu5geYZNbUNCVSac8migbWXNB1RJ+gr0et4eBZLkDggUUKdn/tEb0Bz7HS6xNzNm3tTWNBl19OfP
6OYGLdnZT0Od7q5YFLfwMLlhr5pHjiEfwdzA8kAOOvICCrl3hJ0WGyKuqh8cbYQunx2nZS7zZBEe
bzEtkRhObaaaJnilIsBoRGVG5sHKQorqE4wkiCOEdcsYG1Uu+sPg6oKMA34pNiVFPEMgmTj9AKk7
NvUMIg43gdPhKzGQ6oMHVRn3ly/VVgP39T+TNiHy7EoOhMUX9ZTPDSN7WFV7sTwKD6v97G6Ch37j
j7xoS555ZHG8i4xC1rMaBwNYeGGkoOPEw58YU6+RIdQXV8vSVbwiD6At8xrTiCJVwscjzCMV6uCD
aZZtthSNN9xhY6Om49kw2f4Jaeww40sXU2ksU7AFUSqC0LoQhFqEPIyGp1AMHdbtZnSYWqbvaVs8
UScuEQBOz6msXG6EI3a+OPI9Ace4GZE50T4oBib+NTReFVxUoKIq7J34R0pj/RAdVTvVygk5DeTK
ARXiyF0ZvuxIKCWoNgxSSHj4n2nIDvrKf67WVDstVozL5StZbL/sZvp+0hLBJzgthRP41vx2RzFT
FX8oBVBYEzq9iAa4/Wo7epd3qJS0R4kEpjeBevvvdap3Deqv1xdnepFFblC6UAv3r4SmBy+PHyHO
jFUDSCxEsrUHU0FJtHhoch0+zw6aNMSqrrPVV3xvEGi6vPYrVQjhNHj4w6o10W9gZ4oIZgqbKhJ0
JCyEWQw1NHDGB+CM2o8VkXlxcPdmaxFKhH+VH/r+g+qPV0EJmi9oRJs8144YVNWGvmshcF66DDiP
wbaNSkJE7JP1EyItAE+GF8A1UTbRYCnKvgVcypIBat65ewgX60IaLeY01pLJ/6Iil0/urNi14gYx
49/wqHJhcV0cmzZuH21dwRsgInkral8QrWUOERZ6MQQbKdFDi9EgtzDMeSZciihJ8jrasFxs3uz0
+o8cgVzsxlsdKV7X2p52uemfMurb94uYIz74Vngd4H28ptSmgT1ZuVSHvzh9NlFdD1U5LkTpGiFl
YKlKonOjbpcjppYHER9plBHoRImBXGDFiqoIgha/K+wZk88t3DXbfPsibx7iYIXTuge9X4uQ2ANN
lc/n30o0yBLd7A9hZs7jeUtKJRzeWH3uU01F/H8yfwhk7LJzVtI8jkxjNEm/PzLmRMmpXCIrog9e
Z2CdK8hIDUCxTm4QGmFmI5x55IcB66Z7A95Z+gwH2DZxCT1tRjFO4O2C+aQ/SCcwcuOoxH3FCCfk
2f/EOaP7kwEtiobe8Owu7PsWLecnacckjFvDsATSRaqN6klXOTDHfwe04pbk7GUjiBQ/PyLpeLZF
8VUVYMaqD4fYLZ7bmhrinK9nU/Id4gQpDgTSc+tRAmqcPUcBKpNpD04aNaJzMnvTvkLIPdHMljNx
wgzq3JYooYg5kgGTCP561C8oc40MOGahAFix0nT8d7adq7qDdGG7HO4zzFnDcDE5s6u0hUYlrhlj
l7JkBlmJMkLb/HmY7Lhm6t/xPnMQrr4PbosGlwRg8phRHQ4WKoBQwdfrunidnn+xdOpckhnKaHgQ
cUAbctt+3GE8HNSt7JJYKZzI4wcHpY16ize3nkvBDAazmukM+fTR9+tn1mJ+QD8wGP26Lxcz9COA
GN7NGmeH2b71ytOAs3gqabWZRIFArq9V/YXQd14DuJ84HyGltIzVbN+e/3JgWXJmS1KCwb/vXU8p
eUOUoKz/PFBoi/MxQ+vu9UcKAEcB8IEVORpzpUeniQpJT459lVO0GQhhOlwlR2PM4JVoB38gN0Rc
yVIcU/WDVsE/nffGBWGBAUwo48SOAIyDzX36FRTCBKWvUA9A6IRBHTAucGFQRGfRowQ80lbuPl+e
qCLiV/ukiVTY0o2L/kYMOd3Ce0BoEH8AcYn3508F52/C4auDrCixyHBfYCCVl4j7gIyfA76iA0Gv
I4Qf6zvIUMG+Lgl0qId2EDUPGB9Q/p5JL1Ejjta7OOIkuidbJWZ9qB/VZNDRgAdeMf7CQpwXUWvi
6MouMDOpy64208fnFtUUT2V/J9Px8dsSUMdHQCCwhy31utEkHXLccTYUv+fraxlWezquglv65XJ6
pwADFOOHWf7WhKqHPf+f0wDmuH4R0XDuvx+m7wtmO4KsSWXCQ5oqQ7PU47rcAeDEvM8+OLE2eP/e
Cs7FAeEw4tki8N0NZamtVCnuK0K+ncWxCMj4RtAPgHp6As87SFg2Z99+J0PmEQJp54hGW3Fe3WWn
Lq2DHtvh24ZvGZ+IRvUOpcT+oP9AfaOAMUxU2SJDkXde0dd9n9V1kWYUlWrHCcYNKML5Zx98c9LV
6jLXvFguEu+yHONHc4pHo6GB4Vhc9KYoAyNI8UrnsM07S4lgQ7mJmdcEj0wcvlj468da+fjb9H26
3SCe95Mjrny0KJo9NV5iWmEqYZCJmQYAXVyzytYuIk3EHe+33JVl6nxilbIH6D7ZfcIbrRBSf5v8
qtNFEIfaDtpazIC7rwDBcJGlCW3BULfNJ6mdgLLfu7wgcstULTUzcBZ7KAcLHSoLymcIezi7UqOu
5ZJHxuqdcfB312gpcm7wlWCK1bIOPaJLMaYLVEfgUps+4/Jnr7bnWVSfEf0mkk6wwGukWUOSC+bF
hFLkf2i9oVgaoZ64FsbWjjRXXCIU5bC5zIugzYTTNuTilFk7E5I6PppU26to2fCaBMr8+cxq9PbL
KCJ2tznJgPy/4XH3yWdf4ccYO+PyOs2kblTHNfS3uIEx7YXHPDt8sgU60YeKOEoJGRrJ53zz+Cim
GLoYL0ph1HUqon9gnPX/PPH9pyC7JqZPIja+XO2IlAL6bvNqvlxc4U61Ggfk6Dv5OVs9fZckJo+8
IGlLzlQv9JVxA+UUJWGE/YvOrRHFBtu9W+TXnyoUVUw/pRob5Fkfo039Y0prH7jlMWkGdsE0Y3T1
OCrC24yrJ+dx/Mg09W4ZfbbgMlYY3NzQr5jxxiZ5pudpWX1wARQCkbrScU0cpWmncA/io8TismYJ
xzPpURfYWo5U9fSE7h/T8ljpgoBDSRqnhSy+alsfPve/+iS505Hrg86K5IvyEVO+grJxKghsyi0d
rJQFgPvAKzX3dUbvO2BqAlLLJ1lKvOcnEgVJo0syLJ4D74cf8WERrVhlOtesExArIAzDLjJbymLu
hmKvelOoMCIqt/z0fagntYT1hB0D2NB3a30E17fwxwnyY2HMaEPum6sGqyACLsgc4FpJKvAFxP8G
w2VZNrsFrpeQrSTRHJtehoFUPIJAe4F2E97L2q1ZaaOL4qS9QC2V5+X6c7bm7bpBcnaNteRorBIZ
OagQxNB9kEFC2PkYgWEkAjQg4VjxE423fRRsToiJuN2sYfwqQUYuB77wfvqsCP608VNYtmo7j2jT
Hdw9rvE3nsqsQxD4ioMkY7zvMH2TZkiSxR7GukGk/S69GnypkbKmJ1fnlWRqGDIW+3pECZR5SaZ2
HZgpdpe92SSvkba5uZZZZaZOtanEhfoEJDIFNTUjEdUuapYVeufWOJUgXedjgUnh/+qQ9rYVB+mq
beBI/ugroWukmnOY4PKkjpAml6z8h3pkG0c6Ab2Wb2m4F+8tIeLTZB89uZ4SI/Oa2rtwuoRIB8Px
G8g7XsLe+zUcj6+sOo8O7p2zNfZLyf64hYsEc4XNRklgR535DnSHjz6NR2Bm7x6zq4wE56dXpwe6
sHaA/mH76HeKIgB2ijTYc1erj2WAH4kKJvhUQ8bqMUf2vbOqg9ZYefJrIQ4q9wUTyGYDnuQ3nfIE
P30Ehf/Bt1SCZ7yvyHScjtHgOvLiXJPB9FMCh6tPlFvtjgE/YgEXj2CS80l1Y4TorFSbDZDgx9nb
sN6dzIRPR0jRc1+bVJEjWwL/i97SXDvtd6afu98l2xlR2BsVaUaIEGdS+1PmA2POGnnI879pRj02
5G4yGPQAMWlirXXCLw0W4dUETy42TQy1sQpXUIENDuL3TCXrfM8cDtsbEx0ZgIYOvWxC7SLrKEV1
QwCsjGHv4yvmNWYMnks7usx6f8KHMIEwBaplEkMMZUsv9PF4O/qqDJcWvaVdz1ScjbNYdZDobLlq
gw9YCwZKJy2IkFA3KfO4iSRMhJnUUch/QkOvg/DR4dMcCz3wEK5b4lhodt3G/yDVYkyYcag2b7Nr
wCdbDfQWck7uhIsi/SiGXyq4AaIta530HHZhZryGkA6zLieQrpoT0JofBuheDgdipHIkP8b+PHNL
Yf0LUMdp2NJHN982s6cOt3EvlEOeLJSIdBOXEH0+ep5wqtrR9eYQ3iZXlQgX5M7/AuTfd5l/7GEO
lq+cuKx2ouwPl3o2xh93wLR6+W2vTWLPcXCKcHr7Ap0f0OhFJFzF0C0K80ACMagN9kk2IuXloLc9
f/8f6b8p9aqZVEZXUzXFu6d50mkYjoDry1dJTeINCgcCG5GUwbf4VLqw1MHxP+uZJqt3peu3DeGi
pR0Ijbeb7i+DqaJOll+3ROgSIPAlyGj7mFKT9xpmdG3FaiJa0ePQf3qEqYBqLpEm+XPghZYPKajs
krAss31oi4cstPNALvRheTrw4P+366dtxJZLznKYbW07wjzKial+6OjuFTqps1ewRR9reSjZf9OZ
9iEeOe67keR6JAM8Ela6Jl33+aCTiYBJPjoEkdb/wZcXugwnnkNvw7FCcoAEo8MgbgAfz13mxB9x
ghymrTURxWpx1m6opDrinqwjEzJkt9PW2XTDxMdRL4nt7L5rz91i64TB1SZhqLMwTnseITXLR0Za
/c9+zuzr/HVxFLm/vf6H6WyCam4L2HaSCaSuq3g3aw4AdJ+81UpR0FhjkhLtZaeNGUH3FiOtnHxc
5wDYwFwYPzuoSA0PgWxYJOTPZrYEP9ynugV2R1jSxoxFi4AGlKVqVK+6R7e7V1bzN3wlIZzqnO3s
2Ae9AAIzDgQqdSgnMuYv1jsYWyh/v2iINe12HG3lv9L4p6uq4F4Qb4KA5t7XN0NLcZTrqLh1holP
sqqXY6tXrKCT0258HwS1lkmGZLiyP26qiNl29ZhWiwnRSHaNQWDV5FmRUAOiXb5vt+rqC8Q3kAB3
h2bY0NFAHM7AGakv7zt70wOqfCoQJeR7CUx++yAFWJ25JS3keyTv7fhRvOgSdSlKMosMAVn7ZADn
ldKS+7xd1yLUBoJ0zvonWosUx0qSkvu8zOzgJna/5p8tGJxgl94KzLr/TCBy2uicoJS/xxhkUp+L
PwzPUoZsN8U2vS/4CxZqfYgz2xejabxblpU313zDwbZiexpSMOEL6OcKCeOICNcctnQdycoQprXD
UjjL9wqV8RFS2wo1PNGvGgsxjwPQdb6WH0FmXxSrA6EaQpMT1a79eRiZ80jQgHG2qQW5QDTdbE9Q
rl0gmkqELS4xEvvET3YJlCmR/a8WcfN8a/HfmC/povw0Am9P0mPpKWwFuBfgoLXf1WBSFV2sMZBO
4CFwiAFHP2qdY/buu8GriSvN2C5xm1Rx66gfNUvfpvfHKU8yOVlrU7xLZkVh/cRnmJteH4rIL7AX
1s+Bp9/A1/qP3AWTZrWDhorcjBdkhAVKb+6CAWa/CmSSPctXvVYD5OlYiT64kx/8xYHLTMoqQm/+
NLsEHfzA+HnFHKyXOSYZavl81o/Du/NUnXKx3HXs1xFOJMA2MNpc4m+mqZHfTlT1iCvLdjg9rc8U
dJYpxoeD8hze78Nqzbx7yZY/hGwwn+52IQNWh4Gi2oGPR8HhORgQIqFaXvv0azafh1iS2Uo0EIvr
DP11c5zdOb4jRwqdcCFVaIX+Qx2t/+ujlkATnT4OfX6CfsLpP1Ijjtr7V3eAooeUINAx27Fy83C/
wCPOKybYoidoELAAC4ccd0ser0L3q2Wq4BwP1Bnmppoyte9vObRIcCVpSXissc6/1uNrKKutkqtd
/1w5/nfCNjrDQyOtzzm3PtcyU8N9rEauuDYpHosmj1/SEat0POBk273OhY0Ls8dzFjHU2HoJRzvF
MMAkmzjhALQlnZaFBG/E8j16gF+7e4mRBg8apoOOGjZg6nP7CWZLS0reAiJpjffg32VihHKElQyk
5BfjV5a4WNmxQ+tCke1uJxiJYquRybXumJm2EuEaAXS9VX0x0fe5jGqESJQ1QNrHUBVQZuj2f6hN
UVVBFNh+a4P19o/QtteQFLgR/tFrKqtpjlHslVcqV5X8WxxoMkSEG5tYJ+g661h/85AA0wnunqrF
mkpBE8iaXb/haUFHuJTWW8/WQ/tXEx8vesKEJWQJYsPfHVDIl84rXDWRlD/Iiz2b+/m3ZhX/yIst
w4Yv3QWbec71hY0VQW3n8reV0FnN6r4f2gC048PSwqpJGG/QRIDrWnmNf3E5jU3OOy9PrxDH3gJV
Dts8Khri8jyPdcPACY/Ntg/hDrzFd7fVpnqlhQmo2/eHwpTyaV8MfOalwVeSXc0hRT2myG6wtvK4
DkyN24LUjqbqvQUM8nNByKmHkPHtIeJDk9p3e+21/ppb6ZGIh0I6/2qAZCqghd5HoAxB4MwSfgff
GE98bo4ZVrvTPHF8Y953uHteukVGpBIev6faB7dQ8TPXXylKcP9nqpBuQffUYHZZ2FC7pZ1cWtEn
Vn75gd1sSHbMGunUnkn9/vzplKwX/5m6R35WTQtHTnCQ8AvWML+wCDkLQ3SMsoJwBMVUiLKHGWce
Sx+KZObdYgUmPNvEaLlPViMt/jqKBsR2ADnYIEvEvfNRfm3wDbRGBQ2zCclx31NnhLvUSOpRc8Kg
A5xwsUjvFN2m72+cdL9QIhYI7yaO5jKYvW0bFDdMvZSo3o0pvkN/ly2mfLzEpaSY3qbl9bJtjEYN
Vdsi7LIz1VjhYzl6Og7GbAN8J/G1ZF5h9fEtdfmAORP3VMbOQZZZIXwuvr+6P+Jwm5Syjn/TDink
XB3RWvuLX5hnt4kId+0J7sW2kDq4JgOvllE2hjdHjTG9zUxHFqD2PnVsCluVicpHvoMhIqrpLA1t
jfefz1mY+1T7MVYk0GhxxnktZKA/mWTNSW195RzAoj379yj/48wctGNRtrYgCjqa8r+x8tp58YFk
vAkdp7cUdxaqbunP/4s0fQUpjFCxaoYmYj+0/PgfwokBNTOLtlKmjBDJ/IqJuGV75BNyDsZClqpa
AGQDuQBS7NfwTHztA85Q5lho85YtwQwZZb0quq/iRoPGQ8M7+AEDXTCUJJ+QHt+c2/y8Lzi8qXaH
2Ip81dmJlkUeocNkQrfdc9P03LJSO6mq0aRsSFJSMk+8ytk0fS41QpB5IxQlF0ayuIzvLecLK9PM
UYDkG0358zNv1/eFWyH2kmqqOprmEvKWf9dhAF+xhqumDolZezw1oGUXM6wGDSb93Pp/1aooGqJI
oRMfKPb06vEVI0UJEfzC3YpE6Ibfcp39PkEt4nPq6LVBnkTLzVqChrI4uFb9SRnQm4tR7TEGROMt
6hYdTiGLBzGfeoDkm4nOuZqof+lNmoenwp4KbGH4gQI1P9NMf8TtCe+6oGmzoP8WP6TebeCXuRQ+
fc8WmA+y5rtHyFFWuvLIPoqD1WwXp43OGGaGmoOyOySSJ5c7ViBGxq0EVNUsp+otOWF9RevgBioP
3sprs/SqVj3/0sQPO46kKeSaCSLS65DBu48xF0iYGGbT5jAYZtPWMOYyrw8Dt+vjsFVnXm6Li3oI
SZh/7ufwVBu5MOXz3QSYte88QRgJIihbY3P0y55CtCEGRq+KQlut/W8LRM35vXS1CXd0M9e8fQh3
tS9DW+d0hQEyymKhcbvAFMN45s8Ep4AkplJ6JmOPtHSjAjKEfAU4Oxh8FFWS/YYG+zUCzTAL/ElY
1SMJrp8gFEYemhcPP4LojSbGx68sQWRw+p3+t/h9JFFwi03T3tv6Uoxtaj6SRrhQCbUJEq7cQGXO
BOR5IU/foFHpP9KITdN+KK9XZiaRtlYBkY5xDlqp8vCChdq/IEsFidfZFbS9Nl8WDQ7d8I8Kyn1G
qD0VzAZwgsVcXnI/w069qvtTWjL5j9LaouffPL3ihQ5CYwc3+j2tlTlRX0bTSssIgua5NEV9Glx6
QdMbAcq1ppnlhXDg1zgVnxwbRCIKLdyX6Mk/0KHovd1rvNoVgfTerUtgmbEElsHjhuDpl22HMHtr
DlCGlvM3XwMJ4KTa2YQlGR0PFrU3fEfdYKxDXwV3PppwZCB6OsLsevd8K43zlazjhcQNRcjAekOb
Cttd9FMpflIa8BkHfHwpuy5E32TzOafN8C9y2r8niyc2O/frpC58EXicPbmRMAsqpdKajB9c8Hrp
xUimEG2G69idCxombCxEVEtLmL4Ba/rdSZOfJiE75bGvjLb9KKPgN4UfqEg6qwPIvPiqOvQULsuQ
0Bb3nn3MPPKDWeIoNETm/FnEjl0i4yJK1Ukj1ShJwHYa1T3N/fYFK5VZ81h6HNdZd6fPvNv2dzA3
iW3OEmQPvfMvL3SjEgVDSKOamsLfe11u3NQwqogl9k6bIxBKFyCygZonmxXiHDj+gy2kPOgOuoxH
1t2xycdwLKt79A28oRAYlNadet0CZ2H2gYonNAk6q5Ue3wJcEQouJTS5pgR/DwGsTdGxQWwwlUzg
huVvLMAO55kwgKLD+3crRcJEj+af2uS+XZx96QfKBr4QR1ntBdEU+atf54RUIK2yjvDkXEA9qJMb
cyX1o8xr4KsZHAt/NkW5mZZWlvkIRaPAJNSebpFie5V/hJ0NKms7Hex253muOhNcroi7Xkz+F74n
XbabHQL/6UPCAYtt7F5mG2sTRo2e3zFXIKytMUcaNbzmlzJD9z4V1Ss6GrbO3Z7w3rdbHUqFz91W
e5bWzjAxWGnM61JN0RUa1+g537BzL9GviyppyR4H1OSo/XpZRdRz17PIvDmfAGvr0GmtlD/QpMVd
SQ7ADlJHfXl4vS2DPvPwGtjZyVBMdH7C0YkPI8qiy/cww2DeFgk17MlW+akMMyM6EyLTrXw39eQI
SvGICmA/SKJ5w3TAhv8b8Pgz7QJCrqO4I8wX89lsMTyTyGVgue6Gi39KnXMpnmTWEuin66GHBeR/
vXA2mnacSY4RUs8Pn37/K0XI/Z9HObyjPyPiycHvY3kaDmNrFRMUg9TOdfW+knlSRvvhu8KNIzGS
qvWfZCuiqhZZf9/fqw16PuOoaI9skiAPutCBAf+/BXxN1Ql0wzM1+imovHbJottl9r2UiTt9gaer
KuBloR+Y7HyZu0lgR4ehPNNgpKTJ0rv+q8oLucQJhe/8mxI8Dmf1PrpBF1WhzeT3bU2ScgPWmq5F
l1PQkMcEWWExOuRAdfu0F7dqI1Amt9zC9WwoxDXYop0ROUzsn11RoZn/cVqfSVJN5NRI0OOz1do2
GwYkE5PLO4T3bYYTWii9zWz33L+sTmDXAqTU4pUrBfSjf+rar2BHpFNy2nPSeOXuo9pmwLQnyvwO
+QMQPxC5a/fMDID8YTQV6kBkPJ8Sx335MpN3jR6omVHhWwBeEhtshLO6YSAZnwbkujkWKqKQKFUL
bhahv4g7nbtxgW3RhWAyRgIHTnf894CuFthO6hQKa3DkYVspp+dQXspO9kkTs2LEed8JtK2XlyNN
4Ii1xzHVK7y8ab9I3q9chHSzDn255BXkwLypm0HrajcclGEFhh3+E+MMx0NAQ/gFjOV+kZQwZErz
kkL477rxlQ1CohTiX/Jo7AxIuQAhCOKdDopFHJzYaosmL/72WsV0Ml4x5jcHIGdlQtD1iOOJO+xO
AzPiYYrRc/fF2xH9nU+AQ9/hPWrCy3gkqZJErRb7UJw7BEEcmcwqnwFTY2Yq5rXEwIzS/7kJMUGF
wdJqJTS61AGBsQ7EBLjeXFCfk5KMnEH1IBGUp9r0WmX1J/G+fWe0wg5yXgJb2RhnafmXG+C9XLCS
mxg4Up1+lXsX7yp4UW2YPX524p2KyjTtZjB/7M9DTEf6y+iRLH3r1wOjwLPN0noBYt3hLEpU0N+s
zpE4fdLa5qgZHWuX1XZkarSt1RNPwCRc9uNyzVpCoUD+VCTalpvpZRoy+N6PQazivW447kfgyVqO
V/zVBjmNsl0Qp0RY72aG5Iwasy86gunhHgEjxDZenWdXbmQ6wkyjWPrjOrB34dUGvzFtoL6L17/M
CDLTtV3MRX528dAAymU4HCRGVyT0gU1DCiM0+vfR6lMnModYvvXf/GoUNQPHBPXmrD0yWcQvfB7w
vbGEA67/dje7KFtUDGsMtHZtQuNdWkxZRYwQQkuqYfzBb9I8zF9jUXu/nhDTd64VVIW0j9LkhRsF
UDxx3mXm84Iqb6ttJFjKU+jQueoN+Pi/7e7ebWhSXRkRrDfBV83LilO3GS0snkq5OO89rUtDWudN
Cmx0XSd5azlCSL8B6Vdq4aKE1Pl+PRr+uBZjaciTZyuHBewsISJ87bC1UC9Ilnl7/LxTBFOVJiCv
cVcIcfBmPQmsPyyfc2nrYmkqVhCPbDMAWfArnPhwQkhmCVGaPJWaABXDAN+uDLKFyaJOcfQNez9O
gx/8LKYMglKKk30J2AsFOJYV4A5eqRbCGSSnhXBpNw6+zfD0axDIUbX/enmyJxwzqQYSx/012ENY
4cPsdH17uQS3TqEKAMc8L86VspERY7AisF/ZMCospvRe4RMmTs78+A7v/WbmtgacJnei9iQI4ZjK
NlzvXSmxHa+Cy1k9q8FNDbSzMc3CsEEvzbc4+m6DRHC4FRH5TkSILrREdngRjoQyggUb3bJJNAB/
/bwxoXmmROvRmRMqMfiL4W060dFNgv+SD+6h7Vep/s7UNbsOTRZ4rbpNWSGdv0eLiejdWvdmXHCw
UOmRH657aQJILEGKuxyDiykjNdHu+0GQAa0IKLlO5hmh8OqAU8BmVgRiqLtbcqb1pcv5AWglc6zw
6Hza4htS68KJabaYzk1Jqos+CIMBPtiW9em3eZdRJSgmQk0uXYX+r8rRaUxBjMz7WvTzhq8nbkl1
FSaepnRHTBeLcNsDGsaKNiXw6fDbzF0bcUetWdh53SJBuo8sBcMWnWrdRYWurWQWgeNcMlw8Sj1T
IaA7K/aVnPLk8aZo1QLZsRXyKqpOQWnetbqCnM1SONwvyL6fc5+qJ7ICFovmiK146VexCaK4327r
3ejlcmbj280Y1nnu7/nU1Nwo2cQdfSFMyT0DJX4xSjgY/7NSPIruHSs8XN27afvaLULxV11IZjfO
igmjPXWWJm46QHoZ5MvNp2Aqpc5xJSmhYMseRyQZRE39ac0DcLwEZ+RR8z3jfoY6x15Bq/bDSiw9
oKvaQk3KEvW5j/567QDk8kO1U44UMrAuWeNrCYX6flaTmuPJRIRbixJEnTZ/GNnQWDsC4I3TYuE1
qMwJvD6R1UwURHtogqLar1CgIMyd8N7Ouuxkmwf1RGCMcRe3Wg+clHWpXpN582kCr2+HIFNdk/A2
bOtlfBpzm65Z33FWQEPYM0HwS6RvgN0x6+AQDcXl6N2TzFRlgYUpK7VFAXsYgRLHdYfUyCXayeqU
cyG03tVHghy/etsCywOGWXsvO1sVePbgDGHvFLXX6igrjjk/ZhBX97OJ1DWCLcFYL3MPVF8wL6Qw
QvZ072jF3psTzXjbdZVvU2VfTqRsAm99bSbxvC7145HGmlY0Ul53jFVRAJuQ/FAPTM1Tj/vz8804
L5Ba70gbfGk0AClOpTi0tQRuz2fNx3mShKQ6EuOFKls9tjwoaAbOC0MzelI84s+d5+hf3ClmXtDb
+aj0fUZvSd0vVHTD4ARJFoGZnOSNe3yn/VGgQ3p/OJAuExlw1CuWA0y1fYI3OSgov0qbvqMqPc2/
8V0enGJFn27WOiPMNZAIq36+mRpDlCV5eyu1O22eS9JQLKkxZeXS4oIxO7xORvR9VK252iyVEHUN
oSeFZgNbtkydmXVw1WcuRZ9J7agUQH9rzd/5CFieovYff8CQCEqA0+4MhXbw14tCip6vMmfIfmst
Hr/7yVikXbSAXnSUFDEl0nxBQkF+Lt+Ut21psBTSPsG87tlz07Xzmnp+vDztyAFzrGaCcBOoKoo1
B2nkkKl68WFMACRQQYpTOdeH/+qNTYQRyUCD0SQAxjqR5P8e3nh/Z7GuiQD2bKRbYIYrf8Z5DBIQ
z9/PNKhZF0BASCy8+DIXRpYF/ki8hBh4OCfxfGEbYlKeg7ab+xgNwdY+EponKoeGqs8MnMooJfHV
6k+PrXU52tHF5j2w02bqawnBNRE0PfUMqF8RdYCjgX51gt+DHBXuSllz0zw7jq3K9At354as65Pk
Dzxla6bmR7F1ohiAbYX67cdDngA108Mhotw3NmlhWzCLIHqkhv6VEo+MxlKV6Kx9RwT8Vu2A3TBF
5iOeFPMwLtHPnbh/txz1u8VJ8sPJ8vpyiZ/D0IYefddLubZAK4ZFweLVgKX0+UxsqdSjBrxIAf7U
vStTVuyoYNUf/BK3rucVU5Ji3q/++qng+JhU4MSbKmUNQPRocUijLjHbRKj6j18rKq2tZYAlTjls
QoHoIWMxihNeZQlwKOQyLrhWfXWV07IWAmZDCFlDjUSRngVctFfyP+0HrDnbp2SY1JCqA2g/dk0R
zhEFs9tMyv/pjszP6AidtD1Wmv3siaNftVjmAQ4f09puGgDHTCTzFlv+kO7bada98yVRgxHR14YL
eaP9n7AMXWPQmyON6sCdwn+Z+nPSaeweePfF2av1mCOtrePlhKca+NuPTMHGPv9s8bC+t2igQbOT
VZVFNisq9krA0paQlNm/G0FSQGmEnhUOoJx4WTKuf495vnMrum8Z0yqALZl9O8lCfyiyrK+aAB2O
frKb//Rq+P425u3Liw/HAtAVTpezCaxYbuRv81XNRf0Bvjezg24qSCNj3TJvMVgEA9J9xla8auHv
oSahcMLhM8dDIQYGUDQavQKjwz2MirhEP8xKXSVDIYDKbxvV4DJeH5Ja6hMyNSKNrRlsfuRFQCbM
Hz/9EVdOWcmgJWnxhxMuNWet9iwcD5sC/nu4f9PwSIoHy4vTLz4GZNuEiZ6bGpWQ2zZ1BVCKtWpu
pAF5DjHQqdYN9nxNCnnY7QpQFG70SrKY7ASKem2En5/Xfbf9aKNNAIra+tJPxRNjclyMLxIfspDS
NCYATGXYYtoQ6NOM4FruSQT/TWbrDF6V2Ka+p4XcIMYX02EJC/R2arbwkRpl5gIQ2V4iskgUg4Tp
inDPabHvM1rKpTkT4AXkyr2VbiM5xSB+u8Z8DxNeRJN7VWFIoXtjk9/HMuKnUy6ZF55cUYa+SJ9a
2SNcBr2KEzmRcfT4XaX8OrYREk/vP4kin7aGsR6z/AVNYDAz2jZnyPHI9h1pOTGlVToq3Z6llZha
b8kL/UiaYm00LCCn7vE54cyzqML+aIjHie+nA2n3KkwTi1NquMro7dn1myzzWOMHP0X7D3Ct2wNi
dch58ehslrIMrOIIbg1WQXAYRFOpb3hM/dqAABJseb3hakdNKG3GItXy4rOZv/FTt4EoEsr+flSg
8g/Ll/XF1U815WMgK4rdJtisijuHdn2baBuqquF9FPGSMa6rvCYMbvS0S4j0nVpRBOrSn5QBM9DP
1C9WqXmz0pdRUV9V+X60dLYOyyxm6h+LFyzJJmiKudIgKSS3PrW+ZKJYLm3IdbUFujvYOkwHi5b/
EngyczvonhOXmgc0WhOI0rhobG7RSH4LlxuLc6BsfW/qTuM4FVkBQmcQhTobcR34/aBvkc8fJMQr
pjje7x3qNMIM6baCvGhab6lA6TC5dBFrLR0NVBEaTu4ntTIyRQ3oObxlfBHob6T37hnIPNpVRxIB
Ho/05Ps6F6/1aLUJNHHGr4NU3d2iInucLeDE6FiITH5MXlst2cm5IkQXs5qY9sXnT83B8KXNSM+Q
hPkg+eUMVD2EqIN6kjTUyjEG4XK7ohi0RpnPoyGHsGZHG82Pg/CSXKIL/WkpBGTNyE+OKKY2eXI5
PpKbPg+hm7CWuhKNa7dGYHyP8DRokIR0vdcq416KqD9HgpoEJjAb+B3kN3T2R41yPtcrPtUDdy2I
rlQKIEtRxo0hkxlRW0t6yllAJjSKyCsBKHPNONz5uCJNwPRhdDEDKNchIKs9RD+L2uohXfkVvJJK
q+z/UcfypKN8oka413QqdbZsa9yjPF0jNO7hw5zjeKLzP2G7ARRqXo00nLii0k/n9XCoqylYan+V
m4PO06dhjd04ZdoC7oCerOeID33DWY0eaxjUwyQBH+zaDO4lq73HUep+DibRXYr/mTlNAh6fzoJy
mGvLS90ducRm1esdMo2wezVePEtNVfFy8atA/Afx/bBTeU35ORcRzHlci6bmKEaMSq8OH+zz8nma
lfXV2lHVTwxBoIiyVBsxgOeKgGHL6Msun7MFbl+Mz/Ud5NruJT3Am1lYF1cWtixgfPdndye/ukaZ
avxEqp03cTNDtGlwJCr4yg/lFq99eLWF/edbBk7ooi054QrrE6cLBoBKPniHxDfA5kvernsuD+Z4
b+PjuHEB1V8uomTqT/52DZgtxW7gNDuB7A/+2LzWWlZqxyaSJqBfwzv9ru3A3wSvxXDQl6Vy812T
ZWe/N7WIZRcpT4ekiUIiFp09gOdKHSgvMx33JT0Sz+IQr12C9nko0Fe7L4EhcJAAhDOQEGQAvh4c
xFQELZsSMxqxYg3rdx1i8fgeTNkIsNrnG0pcvKNjjbX3qoNtJB5+OymBVKXttiJCyI2MfEALQRBN
cCHTSXPebQCRAa3ESX0bmh0VHEVoKT/3UoK7T7q0c0OfJ4lpPFKc3Hp6QsubY/q7jnp1/BVOsMF6
pYNeWaYPvfPs4nTai2+UK0lVZ3VTvuew7AfX4JJpZQ+HZvcR01Yx70V+wUH1WJuA3LyXbl0o56GX
auIOfmKiTr0h5RrglbrhoGol5fZb3XQ7Aw/TFBnz/FoLt9iU/77srtcRnOtwyKyjK52pEMAlHYC/
TD5axs/yf0v51ta7PYrHhASG9IjbdMR5bapm4GOjF4L0BzKmd/KiJryOICtbxhGca683uvcFMt6T
MCc6BQ4C+k/G6d4aDmqbjIGKvMWGYIASgYYJVjD0+Nb+k6WgyOmH9aNciPrBYI9RE92qBbnCpM+S
0Yor9sQUKS/t+fbJNibEL9xi80/l5QLb5/zVJdXxhjO/izF3sjzRMCzK/7LKODlhtuy3C3UI6NMi
9z0zRIvuok26DMn27Cxmh9x+QkeWygYtLP61w2wtrZfvrDjtC6/TLpFaDbvn+wJWvqaYeiKZCaic
MpjgyCCe4ktfiwygVLM3EMACaaAY3hffLcbxCPN5OsyanCCnHxpQ46kdNml2zWvR92R5WMy5qXRs
8qm3fEOnHy6EGJk9UYXKr9fbSSc20xzgeuznPAZ+SCyKTopZgK3POxJquxMlUmDB0VNYaCEyIW/P
XI5fbO1D80p72D8htocBSFLH7+Gyo18X9iQxEiTyIaFc35hYxVELHnVhBclDYp31McTiqWRm5OcW
23c8pSHUcm3vm8/HnOxDcWlptNc3wcUKLOT7YMH1oEOOyNejGotD0klXm49jnGbIFz7xTbANiTFy
vF9ZUjS/SgrqbSD1vtxtAJA3ssVeca+zP8p9Hsj60TOo161+YRvvM+juVn08C8XnKm0+uwKipqmO
TYGiiWPNqLtU6XEVrwtKXP8v6i5r8GWQgEABglSAs3K3lIdGPfXNB0zSRJavAZUAlfFwSYGpSbuF
Do0xjLwaY0znNjTX0myCJHCxUnLBg+ZMVjWh88QJKrCJXhz6L4EK4rmQLErFMkygrH9LDwNK3uvV
xPR/kczf63ors5dK4LhlWhkCUsqPJ9CYUp6oBdtN4klgFMP5wvby8TRXxTSRK9kcgh722dbk/6oD
efgTw05RdV676Mf0jJc1HT6AQKfw3yo1l/lZ4VqmBjF5RG3xTs2oD0qbUBhFwbkrY90p1+EtZt/C
NBwmMwDwxtSp25VUwRYoO7K9jCvoWtJMKK0iKhyySmLhFt1eVzVd6Viekru1xzXKkQlX85AU4XLy
bLbraFT0DDGkwfDvqV371aEUyqJ3kDTYYw94oce/k9h6/cMB0zSjdPlM3tj/t/Aw19xTzIUI4qpj
WP3RBSiGVyGaNgaib3K4c9CCfKYYqAu/uHATW7CPwEJSZnRGtCnQGZ6Qv1e4zyyrx3uoKIFS+Kgx
3DlErvZriWwiMNtfrE1SITPEPL6NWpY/pXwYXhaPuzCO0+t2wPDtlIYmUzZGmr3Np8ncoyG/ozrs
ixRa2fiLS9isDzkukoIu7raL/uPqMj77YUJeLJi76Qtp5NuzrzdPN9Ajz9A+Nmj7c916W4s0NvKE
oEQUVq7mKgGzC8nXXz1AFOtJ/T9h7oyYvrUqRCmMoFlMKWCMjXW/fQaavjpPhaeOVzjwl9E444ye
91mo/REp47giPuVCBwG/QkUWhgniSrQGns4zz9jV5lmzn9qhEzlG16Y1sFl7FIDkBymLslEMx8Sv
BGo27BCcyNJDoI0ecuCz18sVlSrhS/1frxUgdIe0nm1Y0yV7YupwadP2ErYqFwJUXe2F9tlG4Guy
oS5OtRT//XeMGRk+9xYQ/jS1zs8oMyWFm6Uj5LIoEre4Wa1U2WeoM4OqUxdHCkAwkzowAuY6AUQH
moF9kMmUbRS21/l9JylxHWWAkiHo87bDNdUjaPSGam6Bqqi28qWUfjgCWB4+6r+A81tj30odhOWa
v8HeAzoddp3ckEEYw81ctW2swWrPGkpB8MUsy8kG0GRLp7T0EV7xzwC3/xR1XaL4T2b42eXVEwun
FjuvH5oPrHiKxhnrmtjuIAUYDBJih+Je2zXHEdmt0t2BZnniZ+90es4Ojgpe2S/dJjFJHyyF47Fg
03gMWaOx0DxarErMmoq0gSiOYdn0Wu3cAKb6uzBOcue0P0UkIfu/NoVAn5nMAJ9WyFMoD7pSUrS0
D4gXDvVUU11ER3+rdoxsK1Hsgjg4C3GPestZcXNFoTHuNo5JyQxBb5hKhCaXLy9sqSlvZG3o8mx2
8zuu2JV3vdUHYQLzRqOt9FuwyTI7b4numdkNOKWCZbsR2Mi+L0q4XTokQaWzXqhaW8/xDqR904e0
1SuUxbTPfcHxKATinop4CRKYhwZfDMXDLQL51nnrLkhTa6/PiEA3Qi8DEvgzEUqnIexpZx0ZlH3r
xggMQskSS88Ba+bRR1qNDd+FJJfX2jDO8B0J80R2HC8gKkP9k9hLjPsBbnzp78GRxEwnhDVBDOIj
PZ7WYPxq47McfdCDjA7abbQL4KKXv4rzC1Ij1ZhAei9vuXGGiv+CRWHWdDgUYkXkvnMxMhhNgHfM
Z7QxLayBRf+EW2b4OmlRwsMrshxSnu1aOqTZ8nnPCIz07n+hSBy90cUbxZ3/XMpfuVNLF/F3NtN2
WxmSqE1d7MXT0nN4wMKxSMaSkNzeLWxB4oiKd8oi585EFdLQBLfnb58Eere5I2M1RSHbwkPM64NP
R4K4vNyAFkCgDTHE80DMbRL895T8ZLXCGeaNwhu8VwouiZW7Zd777zLGIM9gOibAThpcFRqd4isv
9ZW7Wru1EhZ8vl5vo6K84FsVy77tLEFKlVeTSMjn+E3/lheRNbHok5jY0mJbKnhNVrc1nlJGnyOc
RcJPrOBd9CFE/ifcZgpUOArqpUROCBMkcoufump59RUAIFi60CGUGtXQyhpRwzvceocNH5WazVvD
F/bFxCn1w/K98xBuDI08PlFDpexuBE4jeJDwUu4PyxwcIbEP4XF6R/OWfBb91831u7rnLavvG2iM
k1u/0RkLcsM7v99JYo+2awF1LNz+k8713ZAeBB2vjvQVT40WC04puVx3MvkCVQsxa2HCSLK5kvnA
muYleziyd7GHboUu46Wt920NflQ/TU5IcTrDdyqM2ILutMNmoRDjOqat4z1bkLEzYxC8s2sdEJe1
0s0xfIDYR+jfuAe/KdgPVwvO5pAWfJbvUvD1VL9iX4gNaEcn3iaoOkj0cFwZUpj2jHXZwEZTvDgb
T/BkqkW/C9zB8oysKlDWYgqVlgN7uKwavaL7774W7Khwu4NfP4q5KO2GLBvCMd+g++6GAjcBBnCC
hWCQWzswslMLZDumrZOXFz3KRm/tlAj9Tlz7DGyVeME1ceAMxW2EHSR8kceVQKhbTv+u6ywrek8P
UcQ2YBHCYM6FkyzjHUmifgOHxpMHESnhsoVUomhoorRDObbkgZ0BzZ4KZwfmupzRX3hU4JbLKZdR
hXOABONxbTOsGfq8JMSB1rfR6DMS8NbGZ/go+rwUarMcaJxIqk4Q7YpbxuxpebEmlfMMpIiex+Ae
6R/sDokwUfCrUvsZ12kspMDCuMNDgBX6kEz7Kv+/F2+/wsBlJUqdyCR5d42wSXAVwZZ8nf4Nhk2Q
HS1/kv170VN9s/NT4KAFdcifxNmBFotaLWfGiMXy5Ws7+tDdO0X6d7gAuY7rXsM0JwTo5Bv9Zet9
Ur0yHdzkWc/NtHx7n1/E59zzwm/JceYKmJMpoAywWj1GR5uUinzr6e2uUQZ4qJX/ACmhbGW3WjHw
L+kCPztzhAl0873Yd929DIaHDJA5WnnjvFJCiG6VNjqfgajCa4eXRObU3OGOkImOprSAG98aMPKO
7d8gWA88sUiscavp4BtvEC0FCR2A1izjjhnaW6TMbusyuKCczu4b9v9RJeGhwalJTn+DiWV9j4Sk
W1Xla8nz/j2KoLtSBKu+AKmOQ04ffu5GWMBy+NEi4fQHk+N1RK+Uu1Nxy7KPS183Puv2MOFuKQ0x
3J3wLWWUi6XPwvRWL+LNkk9fZscKGbFTD0BJmXYHcy2lRO5dDTGdPSTP7l95z55ZAOwjcGRukXcA
OcjY7gQUOWq0eewJyTzWtjagFQ6X7YaVJoq/Ppx+Ws8oYiyrKwKdyq/wiA+rTITbqfE30eJF2Ic6
jOLXfjS5eFdvn7HO8hyD7FrDOZh0miKGbKXe56QyePP8/eJFxEBHP53CoXfn+OfiTWODnJYii3kv
X0lTrdp46s/vqO4HzJNm4cSADwYqXCcs2fHJgpVwkYAkHzaim6mTCUFU759HyMdaq2/OV25Y6rFX
2bB+Mqn3AyXg1qQCm9Db5opWEtT3eI8D9OS5p7UQMsMyQE7i8RGjtKxAU8HLjyWC/tqzeslJ1CLL
AAdoF+P4vyo8LUcxrJWKBgMFHRS5OC9abgJlOG9obkXBYjXtg8NKhTm1pFExLsmhTC8SOb70Bcwg
PFrPJtfWa6004kZJjlTfTznkeiwfSlCu1bMVu+1Y2wb8Q1T7LzOJtTJOQWw6C4Y05PnZj46elUb8
dgwcSmBCP7fj3Pz+UNVnkUsmp7w4lBpmhRAK8oO7SrnnH7zyNvMFa1+KowZAWK5wpy+g5uGFdc3R
kY50oFHNqiZhK6MQO+Lit+2pgM00SJbDeQVTo30UMRIq0u0+3DGW+lRHxdt3HK/WPvBsiN4ROO4b
RaQmECpNruy+4iYnajIL06DYgkYypjkihhAFoyIxoaT8f18Wut1lWWIq1L7SwKLXYFoJLk2ifUy2
xTw7d/M52GEyZdHL1zXCPES3Ij2WYFBW+p1EJtm1L0IVwvrRhBasWBhfSq1GN/lLjaJV9PQpnJYh
Uz09yuTN76fhHZTEmkdRTIYiaqCSSd1ryWg3jmDjaNij9w2v8/p9KYHTbEq3sum+tLDm3SHB9y+g
vwdvMJsemDhRNKR/kBvwNFYeglbUhJuzopgntRFAj8oDVmXB3BJj4z0Q/l9XC/ZjcHaxWOjNmPdB
lYn8YbLeqOACBVeXQRGSnsd8Leo2qSQSplsU6oITtmnCVSOZTlJoQv4zRDFZx8lahTDcVL3lCPAi
67GfEQtDkF5oWBlkOdzoDCJsJk8obQ5YBtVNhwkWsmHT0Zkduev+6OK9kqzcY3DKqbrGWAWpH1Iz
kuwIhyQhP2+RP9cze1tfYOPjLVxf5IJLKI9OCPNSpPUUaf7iVaLyOpVH8X0kL3TIt3rA0hKFdfXm
UVmqAkYDfByDYnLwnYiZjXg9JTvijDNwovpOKBWGQAvKHt6YcEzDE/opAespBipvNJYzD4KQusQf
EJm1n5vHxcUXnK9LIiaBWJ/pqd0SuRXkkQ9xgOhRGPok/8d2yGOc5oIXiEtuMPS5kfvehEkC6GK+
BFIMXeeu3x5enuL6CsOhibIlrUY+3Dar6AxK5sFwUw4V/hhZlC8A/NNPmi0OEbur3bc1ZUf6yKY7
HtpaRLtxTLZXjNpE2KozluEnjffiZ9hBgBqr2AYGp+bEHsyyjjGo80S95I968PDfJoUn5GVlrZOy
kQlwTtKkiafrRB6lSlBvZ/IgzBi4nPhW3DvcnjgIt5tUAloiv31KckwxfRREm4WJlV484vgYMEk3
z4iSFnxcHlCNJezS0AInu1rKes+/PVg1j3VfCVWBFNr+N2RIPquCPRYFz5faBV3vGrrRTylUMUM8
QmZxvjnemKO/ikzkU+VOOTEXVUIF8z0JM4McrzbmlbGOaw3Mr5oOFDO40zPOvadDtWPBGWmBtktM
uNQ3nc1a+DXghEBn6sH+Wr32wT/cjVI//b7lHX8Yq706usNqJKofHeJcv+evwoT5aEQGIO21g6ie
ys1zJe2g5i/jhQhcXhydEXFkPUB4MkdrJfmwRcHLUIPvOGPKCT65rJHYWbK4or3rAkRQgRiyAkLh
vehy00CO9onLH6ih41+hE2vGNl3ubwrLJ3rhzrS/0tXVH38VOuNqmrZkfdQ5BBoZ11PkVQUpKuHt
GtXAlxLXUsi/VqNT7lVQ8j40vUfkYs3HpWwnEkaWgQxKtPWU9zcxPCTwdXlLUmvy2oRA+Li8MM0u
0U6nlDkQgJOYuvrmrqmQKIeDtBP1suSJgrUQ3h3eAlwMMK0cpbBLG3tmxB+fusUR0GTcOZKNVah4
//Z/793dp5TJnvsjERtEWNOiHFEzuISEjq4aR9bRk4Z9qmcGrewPLGV1Mp3RuGsBfsS6ngyRiIYb
gwZQNkI2Vz5BJzq+N0JTV1zyNv9Rn7N+fIOKaKYhVdmZMQPcmyN8Ke+bZoKIYptWAYvcpyYcDHxf
G2FAejpYqE/jaoUjGt/jHMm4axiZV683MhwdZRZSRkUt1LWSt9DaLzkSPOdhJ20D43creevczGBK
HZ6wTgeIcxupJGAcu9/f8ySbOWLk8fsk5Jl3bm6m2CUYsckKTrYxfnLHHnvZFv8cPr8x2oXqtmm0
+YePmJNhuT1+ZSS1LeOujm0DS5kxGNHTPotL4shCM64R1biWhQKQjcOyo6ZGIK4NUKKyGEnS0Jci
FPbD/8U3rox3rEVtZfG40phxFQvtx8wBf6nP/FnSZovW3Fhn1DREJmG2xbrRpMCUFJ74A3wlD0Tv
WkIYPX6ZM1lTcvqb3eStoZfMNRbI40WjVTqZ1YuHEUnD+BiQjePHiSiRfOnnyciX50o2sLMXje/q
YXmrWNkLhTiKSRzDntAHlMB6bYIajK1SfOVnnZeCTKlALaRx/xYLPLSQk4t/4DvwgSMzH9xKorMD
hPekZ5z5ooN5KV4Ce/tho3fFZZ594RFBkFo69KLPyUu4TbnQmrQ15NB/+MEiKrz8I9Un/2bDqNy7
DIbv5Tnu2h5VZ6OQlSF3q+Aynf+iuKJSF3Okax8ww7N/wEdj/S9Upcjxh/FpQ0/6GaJGeA0ace7u
brqS6YOM9bK5j20LtwCwNwGdCAU1Lcs2EZfyYa2FjspFNuXQvP//p59Tz3Tssg+3FDNOf+K33Kze
e1dDfOaGS7D7XBPPHB6u/lnUgkkjNZJgvgpR11fSMbmsqBdWtGi33LY/93dUTh0TjhWDBeinfVWA
U7pSTSIfoewp8xmEYJmCRX3BMFkTTRESNQvKf84qdaP6LK7J7rWKRtBPdURlYq3boHt7TOnhElel
/BmSXCk5rRtqKphGil1P0pIaQDVXQ2mdwaxLpFCyVr6mc6zbxeTuM2RxOWNiIedDGhJznuJJUjy3
Xn+xhyq/9HTY5smA8TagfW1rshqm2n6xadrGjNG5EfKGhBZBWiL+E7OWADAX7GnDaEvtSLAHTlaF
fH3MlHnI7WZaJTR3GqPhvRFFntqyq+SNG2EXC1L2hTUDAy1NSpCi5IEaQyUa7Fg4WZIyd1bl6v5w
ajwOHVYhKEPib8VGiayLTlsRYkByboBAw/NzW+Z+dEbx0TWgNoD/ySDNxvfCWanw6AsaXedsVbQT
VIHR8S9pCE69x0JtkcspuQnakWFpD6rmtTLO4Xyb9BZ84N195h/QCSNRtPJp6aYiikgPnKatwxpf
uQFZAeDXEidEHa3jjdwpP8fhrcmH6zqDKdCpA43MqXl13Mj3mj9qPQ9fPCS8l9SaS2vdc1Vb+26I
j/NsGRd2yj66TdvN+yOUpMuqupcTtwQLX//XxSU98rKZ+vVa4QFs/E2xGhjnYGLLp+BOF7U7iQzW
zvV3hYl9G8dHBVgg5+c5OeC6Ps/X3StwJCxbrN7k8p2OKtiRyCNbJ7DfSTVeYMBfLJ1qlzqo1Nog
IBjIuz/PLNqiu8p/CQyE9bBNokHi6iz5Njsz4+kizgOClF8XQp8WRzLoFncjtyVfKahW9D6st/25
XkD8icO/vVjdR6IiR+K2QzkB5HYW+5iawtz3D+veeWdluwjgG7bjlWSCz5jxpL6CSpUS1TAgRLL4
dzK90ESH7Qk2iXRn0t52Wk1iRrurb4gqa1SKuBCbSQxpVTShKdNMKQzf1y8X1cs3wuUpa/hwnho0
YlmRlH3D2blQcNHnQYsaeHU87ISS6RRYFs4pXpNbk35esZZ88KbBQVqPBC5bHSaLYxh+oUWKyeVk
OKai+3GDzPWRBXZUUpVGzNpxP6XmAjoML2xSg0kcnOGjHZUFht/faXJ6t9V/aW+T6mFhrEzJQuBC
DevtOibLJansf54FzXFsa37KDBQ0hv9P8+Ge5wexYknZk9dTqoyKFMqSbg3Ln6mYveTA7ofuoCVA
J0DR6svYww3cvCKmqNR8R9JyHt5NUS3rglDnQOlB9M8M/R8geC2unUUMW7x5VvZwgxbqLnlyBRwq
S57duAYzT/+MqkLncoUKNhKEMGKQl+W4V6C10AstCk+yWPi7+lpFrQDt+qKoSOD8uSapm5GrS/1C
rxS96e5rLkhIazm9BLqf9v22KsDx7bvk6M2IjkTVNvzI6BoWJHPXwLRKVPR8soEZdDRtbG+82cSN
XSB/+y/yVPBafEDQoBmGylsejpwLS9vlcK7QUTmjn2Sctb0ofWcqLGkHCosH+aEXlJU1saAzPFDY
U6ZFcIXjc10jopzTQdt22BpJK0Ei5o1aR3kCXqEsJFcQg82bGvOvjpS020BJ9RODTX2BwAXHj+D9
FUWn/h9j+Kx076xLvtaZYKjv1ZvVHAEgzOV1UY/9r5oqj73E7pIAYM4bWI83C1n2AfclpyyhDYOs
hbYtbL6gy+PvOGFjsjGPfdBphM4mRwk/nRdyNR6pG9P0PiOqA8EYgA2PhHh4MpM8LgukAqokGlIk
Q2XClWNRLQb++FlUm6mSWafK7k0af13krMtR2OQoumIHe6DRu/M5rfuagpTptVXw82+vtWr+WxGi
wILhFRObxD+NSKLazS6z9SY++M8aH15+rDvl3dc+4/KIyWlAWWAu1TTntGs0Nms8Kf6YlZsKAOn0
4oUAWLWf68CAxoC9WfIDWaX4OqbbRTrO0skIN078DX5ZLTg3ONjdHW0qDVVj2ko/03FTKsCVyqst
gce1HGImJJgPaOYzMf0LXTXmc+MQRdS/628ozf2iXG476iJHTuYrQpRNgYlkj0VJjxJvf1q+Ox2C
zwSrwybXcp+zRBRr1C95mozW0hEfnOPOlvkXv4U3xJ6G8JGTDflnGyuJ3Jz6lV/HynyvRojje2Dp
emERRYZ2oQ6cnHFTGrdaA7JDQ7qCVr3nKOV8vF9QgEEJdjfuFk30JLXX2MeAsBjVBff0DeFnjEZH
WeTC4QCWV5f0y+S6+COKwU+taje1f0jebtbdYaNsqqOIGvo1KkxJ+qRGmiWBRxt0aj4XsSaMOPJC
E9iMWYIXkkOVj+xWsfyNqU/WmfP7zIsVUNesh9rfoPhqUUzA9eEj11pWzBbo/iOUeG8WNKitZ0Xd
/fh6Y8n3tdLacwVBxz0WWr446KT36DrfBwVeOuWT6BWhRhwKC4G0Oag+jVDSFZTkJV47vdf+UhaU
DOU1B1owxdLnhxuiMDfhtjIjk3hdcgh6eZYZ5f7YPyl4BFMO6kZ3lx7LMHllOyUItlRa+JFpcvwu
nPoi5gGsN4XRAblMeIm14EScTne5G/rmypgWRCml0rwPV0a7fm2vshxbYbGadr6xSvZRh4abyxkR
cBnvMPkfI/bRXkodvawh3qu6y/4XRVZFLAJB57dr8HHxXyfF4dUwXqek4w/a605XPil6M0JK1gsz
o69R4jJ3rtzwJPvEtgYLgni4iyolQAURXNzNlNK8fLiRziJ5EvRZMjUl8h/zLK75zYgGDwANIsDm
oFXXB+l3H+YAp5+Eh2ypIMdiqKXEHg4ojdQQ2rYOp6/i0/Ct1/+fovHlGXtOrW6JbFz/BHSsYpkZ
p5LeVx8XLaGQNlxSkbbgSvJpe1/3qhA0T/xDbwjrtFypxMdSoztxKLubqxp8qrmHd3mb9gQiPKAv
kkZIjq8km5r8Kncvi+TlJqACvCMkjzgAE7RwuoB0dUMwduFVdgEkfP0um8lUTiTPMyw4/yAgtoQh
68juhjQBnB3gWtVg40LpO6xCLwvR6Y07cwVqp9C/u31WvDpQ4y5+pZU9DhocLPeOK8B38ziNmLlc
CEQvBMcPdU4kr+MZGXEfNcr7G84+lSB5Iv9UugPKMph2F98xJJtiYd1h0QQK2F6ZJJduUiwRO9ak
hyKW2k3x+rgd6VrNRTnO6dHkQYINMkZknFBKhkYnQ5/kKDYxrxaEsqxjGdaJuODpfDuBcy9LeN6M
sNUSOVQy2Fcc6A96GMj9HtiK9CXYnPCTfliqOacO94oVpgBEIYYG74AaCUVcUYcEQV27DhRYWP0B
PeuZSL0EJInP81PIbUFairzh16LHA8oOJbXRGSBct4F9W+/KMPYNUB2EB6Kvs5H2pqIHfLymBf1t
Zp/rn8mxxFGxJlpuLYq9K9SD3rFzAIOoC0jjyEAVtxa1w6o/YDdUq275C4guWBz5VtiVRsDI3uuK
2VzFzCgz2EfsvU1d7JEa9eZIeQsmKW2GL6Alwl+r4RQ9Mx40LtgaqMZXz/1iKbYlcREmz1w9ROkX
p+XZRFmFPy4Rkkb1dF+FCcjdF8OIniMz5Gj9WSrmK0AFqBlRnmilEb2lFnUML7JmGXnWTka7hFQK
DX2PuTCbs094XGhQxI0ueR5O6ISOh+ZRcUZlhQlt/2/NPIKNQc7PGUJ74J9SdQ3Vfgy6cBskyZuA
b+sD4e9dqKyBiK0D8qfeGzoO4f4vIGSdpo4wjzblsZbB5OqEK0zHcjoUVMeS2PeKlRthAe6G3327
QseX39emVT0MCEvxRYTVENHlBLW2EZLYTZgFaQuz9kToXQsbAw7sCQRXv1U51ArnFP+Fw8g6sRiG
K4x8P4M2VBn0QTykLuddTC6+/H7yGvxUn9Oa5asnRxXifK4PWCU69oomyXPVTaPLxr8Yz/a/qcD1
IOBrN9gjcGQYKzb3df2vKx58GsZdbrOqv/AKx0KnGi2AksorvDE2MHigderAMRYOdsvK2BBMN5R6
pprSskfUn3c2DFT+pktE4txSlrm1K/aYdVrxWa2Sgz+MK4+x/eFv80CR5OqtLU6pVzoY6tgvoRbn
cNR8iSUxk+DX4I3USmfZzRZwz71De625eD1cKQ5ozFm/QA6Of1B1qgADSlHKAvS1MRBk/bpw2m3R
Wgll/HFKpo+a+ZBHgQl9RiT9tvaLOxi8WdCrsoxR3hL7s0S3deH0D7oRisdgAEueCoYGo5R0joiD
gCrih4VZT5XVXp2VGM2gYdrFgNd6dXTMfjm5s2Hx2s3Drz5vwQnGA105lnRM2EEP+AW6BvHWXNt4
fOue+zh3883oOC2URq+ROt6HfsRIw5gsdZBQKoZF7BBY8vV1YiiS+qWLISih1g5yEt/AuZv8gBjO
EUBfAeL9MFk3VXb2bI6JyJgdwK4ICJye/M8/GNxVpgwQOT4bkmN7FGKy3zf4E4N5rGldmbLGOvFg
FVCwnwQ142UHX2YCPxn5VtKox3pceOBj9j0vcofoXCUXwudfGK2JAftb1bV6oDZOIJFgsBe2apTy
DUgLxNYo63tMFTdBj5AEb4+mwks86vZ0vWQJohjdna8vp0pYoDXa7SHayH8ftDiYqMwhkNoqq5He
1el4pBduHNdztwP44x3Pl/HcJoyaonpgDDopYWeKq1MJlFlvNgLF7oVJCUf5ucY4k1iKDv6IBvLB
W1PnNIHkoKlThExB1TnQpVGZ6S97O8qoLiZjjcWsrMVplFvxKCzkAFrgKSeOlu+p0bwrfTzm21QY
5cJhy0jDZWR8nm0LNaWJ3d4NqWYGcdC7a0+bPz6kvgTEDPkfYWP82rqgdbwDc1L9tKMiyNER/k2n
lCPxh1k2IhwiofkIQn/dHfwwZwBIApWDdWz6OmacdVm9lmHDSuWZqzTD6OLazO7wobZ+g5iTjAIX
HT5ENhxwgjyj/5ZDgYrZ3EYr4qGx1NcAv8S+BWVKnv61R6/v/byEx5Dp9F4fvxhs5fnG7uIz6p6y
XKVWz0U7vqLgmthgGztMJpjlj03ims6HNIcTCDYcmYt3efMO1wKYKQJQWT6SGB1CpPKrnyfwTINF
4bk0nK9y93k8ot5ApdRZqMhVSIYP88Q9LEcUbTCI9wFE1cCEGls+zU9FbzduM7InIPCOYuW4X9Hp
nyPk4G5dbuqWJcyactQ+hdqz1+unC3UKwopKjj1c1duUvNmnwRJ1NWUZuIItONExkUild/WCcapu
MuoHXvNT2RS6XKE767VP49NgLdXWIgAjZMODFY5FuKyELZyx7zN1AsSUlTjbODFgUR2munStco+p
q6v0jIdTzATNEhP3gcparwNZtvuSNkDjJCskrgqjyt2h1ZuIDqY2hId7jA33jaxLKoF+6fLShrv+
RGPoHtz1oANk8OcHjTpoyVN4E0PuZcyzo4dRxEw4k7hM16qPfmrKRAceHZx2mKUV13SVoHlpnyTE
onVfomDr/h91ZnhO3UPJlEUFvia3azFOSRW4t1sUrQXtkhGmk8ZrDCNMU0hyK82oXW/HE0vBO0tR
uAa3rG+kTkEXbAyv2mJi7Kw3wLQkpebezAImYeV7KYfmqBOmZH2nUNzcj8fJjc0tBDQ0AJp39L/W
IYynhjoFH5oLsved5xScV/tVmsLTC6+Xyr8rLVU/QTcq7yQIAp8cREDafAzcxgtCaU4bztb+3P0q
HpvouDYH8hUNSUynN3KkNjokjKx49O6f/WDCeNnTRWDrjcer7vt5TxkcUedShytpfZT9GQc/0hXu
IHMjmRwGJBcmoHzzD6RwpyMPZesykMUqCmhnK5R23jyYUiW4ZOVUSnQZ23WyGEHPB/0LrIYQReYU
gv/4TuY7P2P9jvgrhh+VTLFkwGRZVDLLGf05cqFgGWpNgT6FgKNoE8LkCiGlm7FiZc8hPrTwyUZv
6fXs4FAxuQeEYNLZp+F8lqEaxGFDdv4jpgOmjw0hebLjLB1jvmBG7TMPZVZu3dpvFDWeiaJ8vxfj
fUOPAUpt1gSB9p+ua7JOKUe0chcIl2FzXdsSmhZozAdYxnFMU/kl+2hmwCyB/S6pbka46yEt4W6R
+XxVssq5XVaswwvkMGdNtRCuSuTyXrH+l6uD5z7XOXeB9hIgKuuk3CE9n0Eg40zSnLN3aTAzCgQL
LWoKWh8ojOJjF5F0OT2gVgbxMdytTSgeOwdxxdVtqTaQ5R7eggMlff1/UkxQw4kk+JY7UnAHzOCt
+g0ayljCB89Ruvu0AN66N33LVamXLBdo33wY9olFjKL6Y0rwM81EJ3l9OmMl8fHkFXuHK4+L5yBq
Sze5vQJdFLPgenBBL4zV9F41gQ8yovH5iIs5oFZeLMVmCw2GlMZEueKcF8MXYJpP6ASxouddx0ua
QnciwqjcP9S4K1ELup7Be2JJ2d0jQ2Uxt/dex3veDrShVKfJo4SDcLOMnuAjB5Bi1ZKY7y1qk0ea
17mC1rkf51Xz2yHB6W0nb8hx15IKmRSz28PBOFCZhFUEz7vEpxihCMMKG2dGOsJhVaOEkOWTBden
WANPi8KfDiuKvEqhcX3N8JzO8Jk9ldbmcDVVO6ogCGg1Iw5Re98E8vyMnuoVIc4dCdfFU69oR/EG
cqN95hH8poWGnhfD7J74QCGUJt6dCDEVdSieFzjLjFMY5Fw30a9/rktISAB16NjW1ROQC44GNHT/
ANQmJJ0c882MMrPab55cCFlOPv2SnJ/K5S/UW3SZnhvMYjxvrwX49MUpTQxTct5CCod/3wgwmJEV
0T1fsA6IHqJJoHdFW7AN+zAInF44N81jOLi2bImI8DDOJHz7O2mxV9vo7q0+BEbn5SLMk4beoZ9W
G8YU/q/v9SyKJ/vd8pqo6WqtmgP9dWOgLu4zlPA4vC36kayCQGZvyQ4AZ8BrGUOk2yMW/87Hb+rP
wV0w2Gqt6fTMSaaaO7SrNl77Gfwxj09bIw1br6FWelzFmD0HcAkRjUugZI97MNjo1FBjHG2cETX6
GPAQSwDBWKTdda1IU1CgUOfDrjFJv/FflxZH3aHQsewITSUYmoXH+3O1Ep78gD0Un8aq5dkTLgna
pN2IyiyrMnuFmizoovn9LBWQuJDsnn2JBoZN6RMAVJ/DaXjPYvm9HNw0lshyRQoSC4011d0B5/BU
Ki7VnzVe4NmLB9FQpuePLgxM2fiT6wN/t1wIUXdX+CzbjiuGAyHg9yYyiLeFV5bfHFEmdKAtycHn
HydXN5ekITcILTxnayA9nifCVSgBfEK3CvqdzdeWgjFoYzewvfkIGE8o4zhliqpCzWk/UiLQBDf6
N4ZBqrR34QFYO/KhGdXju2yRc1tZfArC+z5RPjPTKRhzDO1wWhN6fHOOkHPIAVBITi8aiDF9SF+d
XG5vHpef1GcoLIIT5CMUUjLBq0mWm6amhL26fd9IEeguab/8nwfO5X1ZJL8z6JkENGl66hx3osqz
UAMTfLFE/6WsQSPT17XlF3F/1LTK3HIHZPoSve0uUrsgygjjsaw1eBn9Xo3IofAD1p2LaKrlVvDJ
5v/bmmfXSgKW2qPJTUD5nuGZd2mW6ZzOAylHgPCbQmbuBpZH0cPcN98uXs6TY7VaYfrltdSX1ymo
HC9MfTcB+DPOwCnXHuqrQiBmHnqJiJgUvM9oMj22M61/oijnDeAUY2tK1fZsRyU25NchprLAESKH
DxK0bbKxMkQY3hO3JUq5h9hlSSYCP2qdJmXspXtYnVE/e2gfFg66uOAO+26BlnZ5YusDy5kTv5ZQ
h7EeUWUGTxlBkMfHk8n8LiZ/Q9URy+CUtWDjEth0WVH45wW4bNxVLIOLK/V/tdL+7F7RijxVk0JD
n3htv+i11fTHP31Fiidw2E1xdQbxCYIJ2fqMlNZujw4NuUbCVbjIA9tc5RjJNSoF+DsXl76d4LQZ
/kl7MZN0CQ7AEDtMgGvwrhoAE2Bi1jonVR7akT6KUiqbvNXCfoAM6rKiLNL5838Y37jqxmUKRyTL
/r6MwV37qFyncUHFWyi9k7d5g1S7KLLqhd7PxXN1drDz3a3l02Qk9XU4q7HRj8SbgYeZ+vTzEfre
l5swG4Y5NbNijdXOD8cbzr+Z34UHRm/QpgI4OkqqeNjdmJ+Z0HXLgrXl897weg6Urk+BNFOXAYPO
qUiIYIf5pzDbuqM0v9m52bYGPd0Kyi/UbQHIDDgNoYkSWtlvDZPjLrOk6UtN4/wqn/QevC7l+gcO
Ma/xuJKSYLmoY4D49iPfSeqa4QFh5Thu64XZPkWgXbSiZLVWDAwr7pHYAr+ziYypMupk88wRNouG
QQPGGN26mWfoG/+UlbWBtk5bdlDhx9xEJxmBsgFxZ5qxR6BeLqrdTPPOO9ZZ9LGdPgnqW3sa7uZM
pB1FkCwE8/mPlXWh/f/Js112TvPqFD9dM3cG7fDgmoN/r3wr8KD+6DHspfa3kPfcXVRpfPzmxu8g
8ruHekt+851crHEtsuR5cGMACn6gVfuvHHXn5VJOed2A3v5fA5GSmyos4CD8jiL87uFrbUhe8MFI
qqkWLFLGpygz5uyR69pHaGfFPCW7gR6iZ2d4YEa889GZAxsKm3p7KbvRNxB44aLlK50zJWl9YD00
mmEikXy0fL31DGJSno7cvnmtGzYIdPBKzQ5shYiOfcwidEsHvM2go5t7AQnPXpfxhUt2c+JeadsO
wVyg8JAlb8OF6AyhSMlSRSdJs+Y7tjGQoQWpcDYaJ3n/xpYE/1Wib5J7qIxe5cjE9yG7ChLL9MJ+
s+uDmQfvvu2T2F8UTTSFtB1cZPBy7pj8zYIxJ6m1ouNy2gLv6qp5J65TNLrFj5QSbj6X6e28h4+h
4cN/gFy3R0hrdtv6La2Iwe5ke5/izx68rlc+z8WlP+olijp6fM1ZTdzW49bsn2X3Fgg29q5l/eGg
BhOqpL7yfWaEBFKWedHKE/EQ+rYN+zrAUUIx58FGhm36GYgqMJkP/dxeNnrghgguwprchQto0sEL
vtnSlphdeBoYP53Li3dy7lRESe6Z0i69LHAMEInaSrcc8P01lZjmOPqTcS/zUiiEv0IOtc+xZstV
D+5UaO+3U6dpXNqiq0TG/TLPFr+mDydX36x/FC/K1wmYFdgAeZqkVqW9NNyQEtOqeWzwJTbf/qZT
akI0Jbq9RDUJN3O9jzTlVqTezfYa61ib+q/vi6A4peU3AETrQIJyYMZ5H1ByfJQkzvhQRRmUcSdf
pfFl+IrbyH6ikjBhEmEM6lQ5KWSzmEZoS0IGQed2/rxNZ90hvesc1xLpt3oKAEoIBKyRPfLlvxIe
kZSXWVMD7osZzxWGyPIAL/rTCnd7hVInBJsRUir/6rpcxJ1UAk6MzXclYkCVRHaVr87J6/TajFKO
1EMzeOSbelI+yBWFqS00TlOZGjP/lpODTZvyD6BLiqKbKtHBMYHGxDcj9mTgHTWUXy+iijrzONdt
EKEUwa3Qt1OsZnfTurSme7gQgu5EiJElvYmddi1pkYR7qPWSLvbG+IpDWr9inVy/RGBcNrNOzMiE
/TfU52LQoAcn8bEQcKsJdDOIJZJi0Ah66YYQU8rVhEUicxnnt7GD+TWj8AajgMPqwPbB+AZeqQlR
SJKyX9adsSlYfgivjkFrwFg5HZuJmQfgEIO3VfZynXzG9CtKKR5HMUj73ofep9KH62eytVsYGI42
EmvBPBIgGhcu5sfF5Xk1CPXEisM/rqnr5wZqvD++psmOLAKnn27u3UTdKpWokKvKseDMhsuwwiIZ
a95sXbT0J6uNCp8EFK4LUrSuWXwzXsDatJQ0x9CkYmC9b8q0pW9xwNIz7mqj6w4cf4Z5aevNMdH0
keEOGX8qAYSMvFgMENbEyS8MAZA9HoUfm/Ht+8yMr+q9SAi0ll362lU+HhtX8QHQY5QvqhlUynP+
1WK9TTCG2OinxGSP24JccUgv/NyWrxdbuTM8xfc54g+aPJvhd47iIRS8mStyYcwRxEvFiF/lmIYR
aWCHiZ9BPfyajC0DciBVrt62Ha+rx/tRODoPSHhobGKC2OePSVfXJS23zJNEfbo8ZF6hOb7XXX4H
smqzCN+UrpjhbymreO09qRugRUiGoeHMhq7Kif85G6cR8rGpB8jIng5V3cqjKsBI1FB2Dz6MUQ4p
VYSmjlWDNL1oJd0i/nkbm5ZeyuiBNtcJT4nnNSyh3ycztixzJI0FBLG37HmmwIuJYYyjwRvKdv2O
mYnagjqH/mDyApk1utwvPPlk1oameGZ17MiBqP+8TSy14lstiFn/RYfHHQfKsxO+8/HpAPhAT2GC
OsrCBcmF2o31KNpoVeOs1IPW88Cpa6MQ5mA0/8nP1XrPr/IwEUHJrtAwg8M2Bwx7aAN5Nj2bHN2A
Ie23ipO+SPKMiFhMOvUrhJXrRjCziJdpgkbwSD+dAmhRRi5w2+G+1Sk1t+Eik8FLCFaERnsz60qf
OE/+6jAbNZPPfjf+Mztvv0A53yEcKe4lyMB+wk/EDHezLkfh4O8g8gEGxQrNIwHQGLz/KlBdqBJy
w1bMGRQdubw4gEZikV5ZzacZwt1KvYpP/IxbzJQgJvyPJFRQAs8h9tkS+jq/2EusDafj3za/Zcdy
P6OBQd8nTIfsa7QFozjjLZn2E0SnDEGm1EntHBUSka/OnBEqypvi1Nnfh0geh6tInnPDkVoYSrr/
N2cFWySjbwsJj9jEFIw2Lw7tB9eCDDp3Th03YOk7uGaorwbpi1qQQgIifIt77uPene0zmAOwAkus
uq15/PfKXKkiWcLnPFGnP4PQYgLRms4KUWVA8JRgdaxKpwN0Gxqlw/bCVLUHLRVZ2FZA7uXDuQtZ
K4kzE9NpOTJGrE+gzKvJVc0b58tQ1GsCUbuuAne0S/BPAeVRfc2r8oZi0j/pvFn7mXilBf9qtdzF
C614GQFdOfgwJEVVBZZJ7XxPucUjEowr7nrMQQvM9rfGbGbgUmA1iLyD91XEgmE9qq6TknyUANHU
1bSBlWpTwABqauduNfw5qa/JF65NIEKzKi2CIQiO+sMV5s1qVwjb9hS1tiVJeCSeIhPLa8VU/36W
9oZ5LnPx3689HKqCSUWiKp/5qM0zdTumYmXYiPKCDZMKV7w4+lu7ak7cfhF2XA/rXs5p3nfiD7ie
TOV1pwFVeK9KZ9vg5r7vEQ1g4d7jwb1hffBv9yREH+D+9vHUj7mjsOLnaIbVJEvMf61W/HiFI0yu
sKjCH9AQpq6wXnMn8yejkpBOY2T7yCIB+KejuW6UDBEFO17xtu5KR3+One1rtj7JQuWu8Z+wVTru
CSK/2XSf5w+mR8e5kmp590wZsE6uILV4m5dV50DiDsjGtRHBNJyxPWenyxztxQeOjZYosO3sPurt
m+B433dtC+oJnrqwLu8KaazUvhUuCmgxOMmVfIqkSKkrtCwVLBs2OqR9z4CYpRcxOARC08hrfXLu
2ySjJRYAIuL8CV2wSvJKdcYXfDK8bHiJLXPvw9S36NGs/fHB7Y3IxNDRI9lsr02e2XqJLAEd5NsM
pOiPhEvLTiYOyHZtGwWYMVM8LG783pnGdBJ8rLI0+bziHyA9Qe1WJ7iX2C3NTfP/f2sb7pLP78Dp
UHuQ0ANtoAOQ5Vzl/hTKP9vIWX2RfCwoXEh0rYdHJbqv1eR8ID6SCsRsM+IvUABP3FJyxu9S13by
Kv1o80QHX2RFx8PguvHsRLm/wyGeiaCnX4fEnQ31DXGmo4eprjwZsEWXzz8rb5ZSIqAKiv8HFtfn
GtT3+h6eItKO6ReJbUZii4cprqOBwlEq2FTs+4pU8EZ1G/EfUnuT0Rlq6ljj+hfa8GXJAl5NyHHe
43cyIc1Ll6bP9c5VI//yt92a1pXiczYDOVWQNeslgQHbZxybphdXP6KnRZbVKghEa9R3ASXbHahY
KOWjq8UfNTRcnEBqlaT8SFcqNMZZTYk+IOaBBAoT13ipaVVjKL7GY76K6B0Cr7aw+HX59GRN9aR4
KBB1sZs/UmkykYaX0/L011qltIeBIIAXvsnnBEaOSIWFszwn67jUuSc+VTIjBZDuYuHgCpsk4OAH
5jWKZVRrKvYyABzOURgrh5lY691z5sYsaeddY4VpFq3JyS0SZp8m5ql+LsMm9KhG2HZtqtLX0txG
1wo41vvVluLtcJzBdCuUlkFkDeKiGes69ZVK5t+kGnPHoiSJTop7E56vPyrunVLg8GK0OgMgDh6d
4OGMmCO8OD/nYvizrVDwsoaFVX01E+Yd/XJh2ZYfw+YFGkL/BGGegclB+s5Trl26DnnZMKGoar7t
xRrnC/o0qtfZbVS8Sv46KZzH1cvIV453yl3yi2F7Jzm9eTztGjlsqqdOHirok9Pe4QkKQKzgCbVU
1qgoNfLTB3uDRqu3z7CT5/CcBufv4M5WiXaNIdyKOZVT/FzJ6W7tLolYGdmtzXIIOzDdidUXr5CU
ekE1AlzlH+6/z503BdF5CAffhQqDitBUrF2L+rBe7IC9A4u7T0+Q4LpTClZWNgIqpAC8A2ve8I0Q
xG8fpfRpeCiLTFOVaG4I8RKYLo247qYqpfpf/Dv2nBx9wimfpGUX7IiyNZnF+gBiySkT3c/IS8q6
c1dwcaYJvvn4PlprW+UXSgfOl46WSrxHVAondVtcxfN/E2DdrLre9PJ2GBfWG6uk/a5C2T+3kxUi
8TKBCmp/CGqiDfQr3hASkGyvg6UQyfjPAJqFfKCVnibxr5rEHAoxF6sOTPaY1aWLoRY6pWH5Zoxx
nTeVTZ9yItBhBPA0zopsB0kdi7g/pEciYLSOSKo9V4Hwq9lW0JVUEElK2+n9m0e5BT//XU56ZjCy
p9w704DltxnVmvxLXFIJ8vvrHRWnTP2x+m2Kmm7sMfLD47sQQ0ou5qnXC70gw+RZiFxLLwHnYQek
GTnejzGVvBZLq2ucrbguxmGbzMtWMhhAvo6wWo5LgPiL2lQ18gq7L3IHZyx5WLBt5lS8rUp//G9l
Jyifi/7J8eEH6jzj3wwPlxYiUsqK0KLorP8qZ96vF6ak+FlOiYxlptzSpCOCj1EnsJA5Ve8I2riI
ZQr1NV9L9/mVHRnQhuH2E/1lho/F/9DrMsp/H+Q+KJpL5OyYkE48kiSFzwx7KstP5TiRCU47p1Df
wyMYBtQQwHY26iJ4+vOMD982Kaq+bFmZXXcLjmJchlz0t/FL/+p3flhlAhAjUiFwfbUL2YxkHqko
v3MdPwCRC1a8VIWLNXEnbSr2OQd1fgPyEvlMsjOeA63wmPOSUu/SKxCHa2a8pLffXjh2rLCSPSH+
YiX0mnRDeiYUZEKKkU9msUpSubYxcW1wvH++u2kRQyjIh0FBqBsvV5Rl2YhO4uB4Tk03ohUWC1tS
pCAFDuCNwM9B0Q8h6VLL9jhNoRT8Pr6BX09UNMa6PVBl3juXEBjESJHwu/loeGfX0ug/A+dtyDLe
JRuCUno24wmm5lvZcPC4XvR7C8Y8jvVHee+g1Zh1g4yKDZC6t1slNzMR+dXJaMRHff/NmooyT4zw
TuSH/8NMpdfLVeqiPToohbq5EJFXsBSJMc15fRejaNd9Nqbsa1nCNcmoVfpmljt6P4kBS81ysbfe
eW2ZiEUY7ONKapJQHwmFXz4cxhgp4sI713l1OP6sRrQuwNQlIC+5dM8YeYWAf+Z5QxG5NwiwbsYy
AUQiU15K2TVDfT6qEPe2+/1fcql/qByzXGWzD+bIRu6jDz8ZH3/wBDjM3Fb4lTeINSsRolvIabpp
6yl4JCVoFYqgi23eITJxp7K8qsdUjag7Xw3ldTLkat8ToJYXtrh04nfCC7v3cKcahoVKqVR+JBY4
YTvlMNj074497ywapX3KYlWU6z8IBMAfcfxfiDq5Bk4eKLg9dL925Xe+8A2Mg0X5stGFcGJj0IKy
G/pUhVT+wuACv7nDXeEJXFKSZC4hCl0vU4g1rlNTJtXwwvJu6N7SPTZHudWmrNEJimbgFHqifduI
6L2yN9Pf6hXTgY2PX5tw5moUeJCh1MEpt3gql0BHbvScEnoqN2WFTox5OXmczZbyjPVarKhmHsUk
drcnFNRt6OAz5GubVSDGJu6bzuogyBnLYM65igDPIInosQ482bA/qJJJm9t/VInYS2XtycCHB+t3
Ym5lo+bpjb9DHNUDyjiEg/ofBWJfeSN6cqXgLlvAaK8GF9ArKwP9GRdVifkSzYT2MUo4bhjeRqy9
ov9pFtoLEq2gHss0hYLPsNYspOnBymOrKzgS1kGbZn2ID0s5ZsxRhKSVYPugDJfFw7NAH41cQPSo
jnWqzZVecdEdI4XcAj6013iaFJl4VG8GZn3UDGbSfAQryQzMAN8JVlCoB9MRMoyq760dZIbjupI8
9ycQcfSN3Mxlb2DRJU1URq7wh6nj2SgXKK6znH/fREswSaaafi1iXppgpTxYsg3VahVgo9ggG9kZ
Gc1VtbqZBj6b1G6ViMIFYe+wdSllVJvyvdVOGTLVr16D6PkdyZP8xADcBbu/L750cwgo3QsGA/OF
sSVhuerXY0FcerrcXZFqMWYdNDSfpB93k2dE4tD5DYM0iLaeM6b1qRWNcz4+gwBoF2cb0/Y9uKxh
lyV1L4OZFdZdvyUUDx70IUUyp299jhEf/Wtm5t5kuxWE71eeUWdoOP0ZQJLYeOqZ7kEiDMSfhqg+
8bc1wAvdt79LFw44rUIVKGFPRxZu+97E28ViiqCqzQZ/8O+vrPg0D1TIQJBXZQnvItRXTsQypsxg
GCDZnOJJAfYyz7VBjEywwJtFrHgZzhgrrHgFCZuSLt6pjRQGFal9GpBNGTjesbXOkwkZg48wBFyC
GudofgrcuMO9/YAN/BuDgIkdace0M4Mn27fX5zrOzMqJkvxtyILiLJVaE6b1QvsBQ5U6S82USOIv
2oQGoAoVagJVgovP1jacANIqNinsSqZQDfqauEknSwTvvR6Hf+1IY3F/vDs/bC86y3Mbzh5r5JkO
j1YDQEAOOorB7b1Ia7S1av5VEYJx8dwpUw9r4qRmzbsX53hXBtKiEqNkxljOc7L3JrFSvvzlXBjh
SiWnTR93qvlUTHTHNDaAHaesz7753QakBHUB28DYMHl+G+OJwERmJ5bHAuls4M13BW3gznhsuCZM
0+D3bvj3j3bu935GNJHJI/PySYvPffarKOc5Y8kwjYlqOLH/GMTbtIiBcXcDLSUCSX1KAz1nMMTW
9tAscX70NFtXqMvRgABV2hnTheIZgYTEn4I3AHnswCx4jZYCNQN638Vk5V+yaO39qnDTEypRv2Tu
GQU4NNm9qWqymSkfUwYdCNEV3XBepmq26my4T5eX53I7mbl/bz61XoychF68tV9LwBtPAQPIcgUd
YGw0PS0RTPFdmRxxi2rB5ByF+RPPKOD33bPRxkAYMli9Da1rpPLJh9+VFvEbfSv3nOsvj8jpT2fu
kuXNdsoBKQBp0cIOd4q1aAGbEPV99BzZ4brgkGAUbEvzm1lJOZyg+FqF2NhLubdbI3rMOtYT0Uyd
gkN+r2PbcOjlVdvmUzYVA5wba0F1BQ8wYJG12so2MJxH+1YXEMfjCuItlv6MAnc3/tnmlxTTVTYz
CMTK7avMasAUTYXzinmIXBUJJVn1XNjIGihukCfGqTrhdXM/IqAhaxEmxPJUvJVFF35N/Xa6+qTB
H4VywQq6bMu6n+MDpELINiFKpZg42RtkKK3ectw7w1Hat+9SUubWQVdY3oqhgXPEFRR521LibpVq
87L/sDscCQje+bIJpYwF/CUOHO7NRuhA3aUqeTGc13ccsTK5cu2pAQeIHNB6HBzs6Uz7wBstqh2x
yvSrn0BTlNN1eg34+2h+RCOOZ45ekBEUt0diZOgTaX8Y9B6JP1PlfwelD0xBYr9Rd1xA/89DPW7X
R6iUxp2K3ceTkg/IkxyYuTlTcyAPMFW77wsSwvPu1nax1mk/0sf9i+DxO6EVg64mD40FnUn0nsau
wXNh7ZB+w5TobE8H13AtjkLmZcun+oM+meU/G5eAKEPzcKy42KOEp7Cruu6CxiJ0LHSVZl1dEYy2
IhU3FFttrR1fCDUHfPSoVOqHqrSUPavF+iP4529WiSuDGam+pAorwrhcxS33p2mfhZTUBb1BL1ho
bonlBG0lbqHa4CQoC1MwLpLqj3ylfr1L9hNZEoPjYJeVDIj29/KlNZeNHtQC7DuZAJjRxEtBOlpj
oSEJU7rGwe3CjrzAUJEneJohBJtPcHC7666KIjAJ5cwQIePsl6oyinQiht85i8QHbp6oqUZZx1qc
r5IxRGh9qeQgX8QxJJ2x8f5nzt+Kq4FdLD0t/31W2VEo+AWArp6YonAS1AQZSgqvvhVoJmGT87ws
IUaWU50LxlRYdxVYnzm+O43zcSZmIo2OpJyDX2uSNIVqu4AqW33KeGbQAt7ZE4cadFOYp2qi7p84
YtO3GVQluq1vKBsiOkWF48BMixPN+D5Auhnz8076yIy5+66b5sZkbpw9d+aH7U39S46vPR9Nb9A3
PpCyyF2NG0RwMByKhH+iA9Vn51o4DWLpQL5BF2gjbO0UgtgGp6TGqZOrjVJA2fT6DR0abN6CXnxL
n5EKtXfctzZ83u0g0WgROaljSbZkvbEamYn5nOzeVe02clLcJiN8EaA0PUErGgvY/jQGja4DHdz8
eXHntExsGXdR1VKFb/85pfBsFETaT3Tf+0CfChdRJokXqj0GBuor+mk8A1OUXgavCrZiM31ujiEq
yb7iPbFTd+4SbDLPMvvI9yty/XrVXERsTiUZtfU1lTqYsbCzwq1CsEdDqq+bYsSz7wHp9I6UoGHz
69Eq4v6Sn4rWaadPwUbCVGcFFkaX1wMGxAdVG4buBA8vbWEvxp5nFq7e6wCPsPQLBN6RVPuZ4eY8
Q5BOevBvmUnwxribZHdFAL2OGY2vpgD0Pztd5bmkGIECEgkGmZnnnDoP7PUdnDD2eZNprrElp81A
SS+peTT2IN42q36vIqHwG4SHeBzVf9JQppVSA2qGz1KMcRno8/yQWXqGKCYCwzpFDyofzyzdMxzM
nP714lMU8yQeZc78HiDLq6XJFRojCNW2yQSPwtQLjIxeNOJpGGbWSrOVaQTOuiwTv1j1DwUIWvG4
/iUQfdanastmh7aRWBXW1mdyG8INXSxwtbzb62S1YulWyi6UuM0ab0ISXVkeEfNFR/u0GbTqqlNm
76WmElqvsfc1gAmDiNFy7vw+tq+wy5Yy7pOw+d9CRfcSw7y4IsSpMmVaC9UCLgoSWVgrUl7og9zR
LWTpcAkDR/k0wqtS1MZCYZE2SeOPpMjE8au/kQbuaDH40KXuufo4HMj+343K1MH4IuPfPioBzcx/
pPk1+955krXd5NhckIyVpjPMzvp1cTHkI3Cpf/6PGufwt2/5SCoHlnS8e3xh9Q+pSs4INcjgftOL
oJaBY/17cj5jGE2T2DblhtdJ/AEVWWrFqoHbTG9iIXEvsyXw5ygzApIMjscOtXUfMG3s1spLxJOa
8nCDsHoc75nHoS4oq18bI7qN1E5pbSfbH3DfSH9FBpsNqgOefI/FBQvO5/LaQSz2YrTeI8QC5vRW
TxDeYSslqY0NrFCcQ1z+5X10SmeAK5+9Kf/ZPPIL/4JQF3xRb9DqboUDbl8riZyHEKnZQoJLQ+rV
bijQG9folx4x7umhbmcju7xI3j7lU7kGOIFiwVBHymZMVkJQBqOheQ+c9PrNqvhJjQ9eJIqZRXbi
3Fc+tHX+YZT9wl28l+D/BiINCVe/GrfxaX59eavwTisEVGhCiJaoZauz1UbhqwV9sVZ0KWNXB59O
/zNqu+VrlWXNQewTe6jgoOfX+h6ZG48rIQlYJdHNPQB4+ImFY7ol3Tg18QH8tmEt/swgWs1vv1qq
wdCQUbyJHzT+XEy4aknmxzBXl90waYY0SCVR6xuqVmFKFAbiNJG2OjdO8iNzmvXQ3CpHDjIKmVxz
MTjr0siQJ2AU4GaMkWJURQz80hUGQXHuoQS9ebRR2yJ4R0fZjhj2WAczpichg1kxPcQ1UtTnvGj8
8av6qCZdpWdQZ3oixMw0fTDIVONN0kpwIduMx+EzU+UkTih3vvqdZNugFjVTPNUxc8VO5NxOu49j
cF4PwlncwEn0L97c1oRWeoM4DgW923NoXGYk6d0Qqm5QIG+Oh6jszi31+Crf8jejX0+KWaFiJpaF
DCPWOEXVUfyGjaQOtbM3KvomdmAs9O5Hkq/LVz/vtrGI2UGiTlvJjcek3FP+4qmyp4wUzgPWNwVZ
zEZtnd1T6ie2HD1PL1tLJR4upVxFhn1M5WNRfyCSUyARVaDphBxxwFWq6qXSnT4dedW+C25XpcnB
2mf4zmXwdQjSzO25el/N96CB2bR0ehGOeyRW9Ay4ImgQXlfZjl93OKuDzvWxYOfueV3KNbp98Mb0
t3fj8UdhCnCDqIhPn3xcVfmk46YcGC4Rqlz0xBcswYmOBKa1JFSjQzANzaFrYyehzd9DlvMrURiz
zkpmm2MvKUu1W71Spr4o7PiyhdLJgFQmDCW9pyoTXKUlCDDZAKfVOyfDuUVJxFiWihcAM8vWfVPj
WwyQdbHlk4UZUhBHwjGviMfXrTWa8JXmq55TRR6iyJ2JXzBvx+Mx1R2mAjZBa70Jrv+bzzvUX4Pw
2cAud/livzkr1p6uKBE054p8s5nGXSaujGtav67CQ3EGO+dCcGkPNhgNt+SFxc9hB/iIcHqRtdEo
QwdED0zf67ytJVZdv20pqoyF91oleer1m7E3X/+04VT2ljqY/3sRMsI3vuo+vv9U4emohe45gZCM
hRvgjnFcTFZzQOINYVHXy3otw9OAyGz4xBVsE6M97Zh2Qkoif9kIgZpLOBnOpCwlloW4GFelxd5G
ur6EyaKWy4v4bMzoHoLJxxW8gvH2yKSqoiM0GMEIE59EjCvcpX0lRB74j+fic2CcGQNqDk7Y/GNb
aRuxEdtC4nYJPCbnvnY3St9i/uYPNphFYeK5XtLHGZ2DChxy88lZXdw/Gt1oo00wrxqBrccb//H7
WFP2ZIwxTY3pbu3jhjDrs/LEU1sWHIE1zA9u5c2jRVXQnsEriYZQNA1L+jaVN1nXyXcXSexxXd0C
6UGByijX/NVCc4s0dJRlZPT7VqmlY8sBZr2+p9I2BHjkTOBoGMC4/jkq3Ems32sZ/e6JcJqTRKak
VVwbQGVf1ptVYOHSIU0CJ20GSawGHkhrzdqkQbOKbVIf3xzwt1befVNJ0fxbRuZ2JqY3QnxEXXcY
WVfS+YyLTiqEL7qQfU8uOmQxd5IHFOtwOHdI1Pe6MkuhQv0ujo+E5Q9PDXEHMi1Mh/HKHxhLovot
rcuSa/QDpijmXO/onVEXsDT4llkzZfX/xep8JqaD+G21T63s7PU+8GZ96BO+0ThSx8qKPVM+Cmfy
AzQBfH/GDXmYUWRLT0IZXtcXhloJ6nMKXg5ClcaAHJUFX4x2aTwQIiUdWTKCIRs88lkr3DqFSaL4
DVXNXDcNyvJP/7LNDoqDDWQDKEBqqQl8VwUH9VsJP3WtpL1xem0f/8vyMXx/+O3O/7HHd5dP/cvF
3n7zxfzKc4hMnX6+J5f7750GCgnr49yLS0CZ7Bl3pJXr6QCigA6HilPxJ3rDoRIkqtkol99VdTPL
rxM9mct9Q+mUUALylYdpd2YJKwA0oUV1h1EOFPGw2AziDDYGnQRuSnpIyC87kpR3Xi3swpKTjChj
fs6B3wo7lYcW6lVz8nhcDQdV9RC43ZPPcEog9jBICWSShPB/PlMXbUxQhlvEeJJpO9r9GyMunqBh
Ckc5mf1RWMlyqRu27/frlEqg4grgcRsHASN8hS4z22S9nlfUjWME7Xa9cOVwGgvVBHwpRAa4asPf
C7S/vWd3FWaAWHDC7DAHtnq3I5h0RALMHy+5+TDjPk8jjur80gPajtd0T9jS13tGb0YW42Y4RfKQ
lZfLWjwd3uasIVFNtn2Nc6vf8HDys9vUOTOR/+ChcuyWoYdLAD4jw0SiWZ38LQStOY8ywhSflnp6
QzEA0comb2i5c2z0/4jGyVXrdJVdSfp2HcGHCOzNPaYh5LdkutDWroCNP8TLzMxQqvw0Pu+q+98u
5apL7IcHqc9vtVQ4xe0KlS4wal8bhvrLJtrZEIBevigyA1zDtcevMIfShoTUOuwtuTN9mOJl+5Eh
dEiOgH1M5xqBUXXAhz6Ge9nu25ZUWzHQ+R+0lwbMn5KrGrerXCRJuJZ1ETi7wnePTDHyMqxncGU7
E0pHSc3PjV3XND8LDZ1oRRcwmvSN/JMx7BEyRYkywJ9Zz/+NSc7pBIveugo3moIaVlt1A3B3IXxV
8tpOB6TOwGlxiut4KKiXupnN6WD58nCTnuiIO8WiaL13mGwGK0rGL09aQl/0YHWf+6585hwtfTzo
HDUS4dITYaosubHjTjmG5Qj6duXlMqAXblDEIsYrvARVpLFq+MBCPHCdwGHcRZ1MoWo7mwwWK2xr
DBjdj89njxtWErlP/5pogvECj9xcCqtMsZxT13ITF4v+HwSjdoKV1qhfie+kT9EqJBG2yUHVCZF3
ieKPQlmyAkJFeL+2+m5eh54FVmGtruKeQQKn55O8F5QwcloUVXk3zDGp/SnjRAvwLxHLhNMgTMD+
d+Zn8nOC4eBWc13NBk4FCvffaWG465tiZn3xGmsIgJdlarHnCxQcOirOqWw3xMq3OgQSQA9Op93a
zCQ9w4D3RAdoDwE0uGYt1HCxcz3tnfWUrqFqOnVqLTVjsIrlRQ3Uotm/YsRAZOF1RBTCsUcDuBtB
83iiFzcfjf6wAh0PSovH3dAlBUl5xV+uN4ddf2I7VbR2ZrLjxGVApz/UfQdQ/+3+MXnQQXqK4D3d
RP/JdMlsSJ2gUpOa80GnxkbRggXhVw6iNC7ZGkhqVIG2ySBX5GV55qEfiJ+Z+faZ2/E+byTWSyIk
d7lZF63psDq+qUgiQtBJDPqiP97sVn3C/HcmwzKRayj8YH98MzUpp4p6jqF0khwqALmOIssD3NYn
BrYjTjwOvPm04kZRRTJ0/1VhK3wgPzZPDgNb/EbkIRMi9cL1v463RhSLWYgpLEam5Ww/FG4sWorM
7dx2kCasR3Amz8QqMHqkMkcUEgEQgVImuJzFc8eWovzlj3xG4KcxoDLt6SebD7WbwrqBq/TcaJ66
mWiSOx5xgUE/srrL8q+HNXlimp9vzcDPgmIrL2xPBFLYKA084neCiQYVVRmdmgW4As8mm0Nx0CN6
oBS/vtjgJH1ffChWJs4HhIuk/1ciIWMDQ5jHgmexASSCIpYjHY5K7Hl1OrOVMTgVYpDtmu89tu1L
OuTZuan/yQQsadRZ0aiTtCW8hvZedUd7jLRWqq1c8bUYXKFQ+x3AZU4gVXsu0XNpk56vD8FrUyrT
izk9ShHH4kjevwkjRiqLvXrgOKl5I7XO537Q/CZgRWUORyQJ3dWQ7DjfoxXkjbgQNW++9NIFp/ah
3wa+D4Ayoyu/ihHdqkhSaJsAIFUmY6fLg3bpqy9OxI2b8hHKPIqYVq4nvGPU7zmuNWUwcLA9StPY
FnPEqoYGmpAis8zonc8Q1K6dEiSvhPDO3PhGa/OoiVzX0UalQXythkgUcOvetKZfjsXYhlbyDBh3
Sk9J4H7G4CALaWIBdova4itcpeiaXPNct94YAasV9Xb3K+9h2Yw4rPrdalE5NhOc14xM3fMZrok7
DnWLcCKD35kws5PMHXGscA2gXylV4PQOrs0jnDEO3KsPoWvJNzGrmG7RcB2TrMIX14ldgMcJ2iLL
bRaIyq77d+tPZNXpmYNQ5n4HprqBjplpW0FoF35CQUCe0bkPnfBzTPXHl6rl68zY4Tdhon/UMbB/
ey5CzKlgQDlH4tjSvoKAVXADglig1ci3308bkvLBu/eGWNkesY+bmUhlWEZTsQM7K7S3W4yuj95U
mwbXJ3CA/x8PvlsZa73/dR/XdS8NNtyE31ZY++HMM4YDFOkslirZ4QsOhCyzPShuSqXXM+0wdTew
9kBiT/sZaIMuAi85lO+pgqVzp9GW3Q0PsZKfRpnzGmVbSzOkGfLx8WK/aou6xa81UZ4R/CaKNWVb
RlerqY9a6V2/Vw+9S+wBocXtLeYj6dQM4sdzanITESTXygLHTQh5wyrvthkpnm+s3mHLIuvyw2gt
IEsUMMSCoAPe0lfZU4d5yXcL44J3EAR4JeXwAcblKvsyADwGRoFiBMlUbSzlkewHT+apkb649yI8
BRqnZZAFrpRKBoCjteI96fvIw72iLN/GLewO/k7agqkfa3xcDcNBB8s4qwgsSnRz0r1g9Kcng6Ac
kesXRvAcACJ+TdXHcTO8plDM+30rtd8CiAAFlrImOy813ahI7fThJDofIJBdJEdsm/0O9AXUHWxW
+zCfqTf/xM0H5DKAvhjWf6m1t0UkFzpsWbgF/HhkijXCgAGqTLf7svOq6HheJRcXtkPCpCHnQlun
KIRI7pdGRyBW6AC9wXChcSWCziltHVpBTJtpVJAtfBISxx7sjRtX8IlhW9vRR2aMRyrUZA2aPhEu
/9Ga+eVzzc92EBo6ObTTZXVTcDH10Tf7fZV8y87YVys/dRtqFFBRIeJorADaQh+D1vUiqRD6kTXw
0mKqfhTAJcgCaue04J9xjmgiYZL+efxScSh/X/gysqDznGc7dh1J9MJ9OiA5t0sjwsQYytZopcN3
ECE1mClzemBePC/WiwlpJKMHQoyZ5dA0FZ8C1iTZK1dFVl89EX2fjIUVTss6jDesrp09Abi2vPvi
dOFzHDnyrDJWH5bZzE1RU0Wj/xTaBfXv2HMKNt72pOnRlhPbD3m2nNqMPYv/GGETOcnEmCIbtDSJ
iCciEEzfF5MtaEbQIgV3Yad6nPMpFaR/A+Ik8Bw+RZopWj0RhCu0o/348cqY23ekJYcre+0xflk5
URYsdtdNYL7EBulBg3hXt/jrYDzHMCIZGHHdK0JkVxWfmlofNWSUttlkvJYhYbbbDzlF63oV+bTv
7AnpdlXI3XMQsXGpyWMiYyDGVEH3n9a/Wy4jrFuAt3jCM9CzB9W4Ht2sCUI1phSbGPMrODwXtV3u
y1vXvBsgJT+OFffZTnyrfRNmVI/w9JYaU/Bs8AmxwwBTJN/uVwiDTYt3DxWlLa6NyBa1ZT1Dqb2N
oD66LlJuwQ/YbRlFnBgsybuyn1xpv95DQb3USHtuwEIMuWSMXRnWYnK8MPTtAO3kHBl1Tdi5LcwR
ThbGtC2QcQGSutD5mxxHnkOpYLH+ZnrIKGzW+e0r20kTWzNADsgm1WN7Q7zA+x2Bs9VRVg1Ev/Vq
RsO/pcvjHFqDYjw9EK2fDdQG++clFBUBWzxwrWl9JREsVnr6Mps+MxDx/IV2mqKyQaqM66S++QOE
lgm/9FdiSCf9EcdEKAA7UACRQgX6UUn2T0+eZidI9HA0GYbvsuQiOwgddxYv/mCbdcAKzGtT2BWC
6/GLTdK6dbSZPO7LXu4zgP3/AZmgHTwyTM55bnsnCyICR5J9SWYrM1ayBnzUUW0PdXHSBV6GY1iC
zYuGjXv5a8WRaU5fALAwMWIhYCzChmK1Ts+DYzHyRyOlU1Dar8iJIKBK8TEXuDRifetg89wLFjZq
auax4Z7Opn1WYdYXV46QbRdPJInXy1BTZ56r7XZDyskbhTbWgt7qUgidl9OU9zWWt6A8M4F5tn2B
Oyla/qPuUSQg0wTbRb29hbiSkAMj1kxBtXc+CvmLw/alH4J++rIne7kzRltZ5FcsITJd0pjazhzi
VTksLEi6ybjYd1mV2j4oPENDJM0/Z74pTSiYzcBTrBCcQruoT96Sev3LTmQT6BTNjMXk3ApwdhRz
eWTczGD5L+g7PCu6y0arln9OZaVwHSIdr5Z8l1+MbhLySbbhHTw71+rmq7ThhbHTXqyVUimeBoMg
vhLHusT0yoFS68CdRlf/RaJ1rIOxxB5hZPz2ex2bBAPnRmX79DU5PdeuSedURmk9Q7dosNQKUPkw
zpRpIcS+gjeMWC+7WNjyk3KEbXvbtnDXGEZY+KZ1SSqn6FHHxIIBQ4tq+YIZWSSlr/g6lDcztV1N
XIyDrs3aI87K79vVS7q0lLMauI2MJD1w9P9uGYTSOKqZO7XvTvow6nk7jS2k50FlTEW+oYVJqVB1
qz1kSxTXAFxCZJMOl8yfEfwhqFPAmhzyj3bwbIobB3eZRjVkNso9PO90d8NM65ODV/kkqyeWwLS+
2K+aiAr692dyT6QRXY2+klkw9ZreaA17dieyep/Mt4x6JLuhQNDGK9TAUrEDH5aRR1FuvHh2TFcg
+msdWBhVHPLjNY5iAUpR4rdYKlOwXhxbqCsg0E5XkMKvHfV02VLFEHqIqICewFav3xiZ4ibltArx
0LsLKeBNWjco1opX79ODz6UV14W6JQkqhyVMYttJ+Lp62ZpdDV6BWSudNrRBRK5ZKvcWZpMBrGXq
rswg+7puILEDC+jsIT5ASmhQPKK2tTWFB6K7jVjtbc861KgVjNhsLVhRBuUdLT1GbC3gMmUTMkke
5jFhBraEfXdQ7KuNDkFG38sOorOxb/qlRxhwsZVOfr00VGyVypObp//fTs4ROhUfFwKlBl4dMrlY
iojO/dIoeTQNGf2FntX9tHMZ5+22Bbqxz60YuMvxmTV2qCPAkZj67PDvGvYgOtdOsH1mpEahivPW
ICnoBMCqMgEKUWtvubwgz8kSzay6F08Emmu1qLI0I7iTL6WnxaRsu0cbJIK5zmnCxZYjX6e/LGfo
KClj7G5lSHSeGUmtQB0dqqeAHEbopVzlq2Qces+pykS+mxOtqFXnm2XKPAtDgPts4RyhCAJ9LEUM
vQh5vBDa5rZqNyaASrUoYrvuaHCFJFUMLEU28El+jQloSyuFPEfKZnvFAmfBOfMfck6WFZbzeO+H
7Mm8GY+fQ/3ZlFZS9TldIADVne9nTMh681KNpDAnf9iBCitEMWg18H9DHjCQWykkhy6PmvYQyb8d
IBBA1CNtN/7bKv6KPUESYgcYArdpFnSXNxQMi+aEwWQL1wEIizw4P3b5rci4NijaJH4Epmhgkfd+
4qaMDWvs6B2s2skXNdlZhdWhpZVfEIvd420aKTHNnGRu8CsUojP5WAh2sURp4Ws3bcBzHmQuSuBE
Z0PC0xCrg6hbuSd7D+jogLYBjGBtYbhNyQTjBVZhtlFs3/5E0QMTjOjIpNW04dsoaiJju+y+BO+O
+7SclkHSIy9WRp/m+Tt0OOnOdB7Bvn7Hh3RqarW0h4hCBQcxT2B0hk9KczlD73WwM6l+fJEpgxUa
/k7dYaiIokwBHA0BRD3PSCM61zKRb6gj+ZgAhLXBTKzRDwE5s7l/+9Fi/9fzIOREdi5C7zR/mOJs
e1WDlHjDg+tBSVmGU9i0AhQUowryJp47yqy0c2PkEEKm0rBmUr5SW5p/kO8CbnhlM1xTJDgHWnVQ
RIcfUZT+iYEoK1HFI+PeGduxX7X5azNgc3ziwRoHpRD8+W5kDnFnapg/3ARH3+GYBgsiov64jeO9
jhws1i+sZRFOuSo/w+PLGSnrBZ7Yd7jCSc8bQjlpIkdHDpgwxjcTUJzarD451Qp4ubtNXsdZc2EB
GGlXRaMzNXqOHt5BX8KbQEOAMnrW0td1BBjfCF15FxacOAV63vWTnjaSOJKFoQmfcrJSyXjfj6ye
N+IPKymBd9KGjyWPfBVpkBJ2B5t5G2KYjZk3i1Yt1f0hHKhcoCWvzNl/qj0UrFhbsUhinyIXhXf+
+QcPcoTIHeZEn3Fk21QD6+Ghe0LOT8JBvlqU/aBBK9J7FqReAKRwoOeaPormAfizCYIacdjK4SBo
oEvWk79F6xw93oTN9SdcD0LuHLPoqM24quL/+7iZjo4ftDoKKAhhElOzQUzxX1x4ZvMgJldVeRVX
fTOS2Ny+eBlU/6PgdPQ7s0uQlw4fX1Q4NPmfsBViiggtFyQo9GdTi+SgR6jchiWdokhLo1+TRb4B
Ucijjq/aTPf9hiFgAtMGRQh4cR/sMf3/mqmRS4+ypmioDNlDB1eadjuNDGEO4JY87F2HYdkmHW3T
A4iF2+5KiBQVhVp/8Nrp4JLy8ILBlGBCD3Z/P+mUpDSihNZfh1wqcNxasNhtZmTPRbe/PCsuGKOp
G82wmBmzLtfgEPK1GwaCt6OEOB0N9mE7Y3BfdSJ9rqUaTaHILyDBY28OIdk/ONovAODqEPXTVLFm
ZMM2doNMeWkiLru0NZDwraknKA4p3mFmjLYWAIWC19B2E+2QiRbKnQ9u6oECBpQaL+RXw9lIhcDQ
tGPvNnIoLekvL6uvO00bj0n3A0PV2TDfPS29h1pKwdpCNYgs/uTGe/xL9+7u2AnZ8/tgIwfsCMzk
TaCO5DDx6Gzh9sSJ78UMLJcwLJmCkPPzfOsrarzN6mJLoswQ/IKweLmrdE4waFwzy6UDVWefZE43
r3upNO42quoCrTI5i/Xal9d8Ym60Jz9P/ll31P9i0YnpzcxwpXRiMPqAQNwazhi482GRRxn65DQj
XbAvdQnQUG+fvlUJcs/JHuQBbEtlyr/ohdVQ1nr3hNrCLS+tZNEDUt25+fYUQd/P2NjdKogpvKrZ
4d0a7LFpyJx+iRiHB+jhUnSSGiyNPkCUzDaAVdYms2vX5ITwd7KNjdB5hMnSL5TIIwZV8tfBW+xp
HhmuPi31oTPPQ848+Va+inlYfktPOIkPnjJnjpKhYQixEko5PqYpb09/Z7IuBML3/SA61WR9l40q
kD6I+7Yz/kg++8eNi23UAAftz2RvoOMv49qmXcA2skgdGFDhwgfhfnHAnTBr407m9n4BhDiU9ARr
9zHrQNGqsY1Xzhsw8akyERPsTIItvDo5hMyYMcpEAeqcC6Oj6ZQ1BKQqzv8PFHKrZkVTNOtdd5ai
oyfcVicm6hJ6EEBvMvUAxlaNGeCKaXB4/q7o/yf6OlPlCJiIaSajswjOLMHFtT6u4DKnfikninF6
pJx9hR6LxJcZcisghvBxZIKlGFWhgFwFI7eK7ph5jbKDSksLVZdEZsShWXNDUhJJ6gHX1UFrYsDz
vgq4u/7QHeWKP47FYkLDEYvqQcuh9PxueSNDkUVSdoPM7G+slTuJdr1FHlqH4mG6m1xhyCksRECE
ZzkHs7nw359FnAPWTjeusNbWZhci80pgKGWMXFibGmYsEq7r6ByHukXw1tMUgVYzkrRNowyfa5bL
R3HaRL1jtritl9TAkQqO4j1tIAxKNmZmw8Cx2dbh5ROe7Mq8hfuNcrMC9gYefw3dJLzdZEY7bd7d
RtsTRmFLdTUERe7BWOUF6jn+Z7nfN5rE/44Y3lT+wQpDeExg9hRs5EJpCUjxcX25eYZWjGKDzFoz
ebT83JZFC/8zk8Z6iwUWGBRMTeHehv0lzcE3e91aCT19CRQOxrUx52LdbZ5WP+KTcCMelJXM4pc4
/NMblGjRCyhlaNE/BsMMqW/32Tef7vGG3VEu53CbrANDVUejM422K7sjZLNxbKWU25JksboAXOoo
v7xo5P8aKtR6od9DAMAoqemOvLyCtrI1NWLAds3Dt5VeiOYUVkDj1QKVwdnhPOufUL6QJdpoL9Xf
sPuaFxwQHqctPm33a5a7KQ3zNPZ8PbZyrCZWbNpaem/IMaSVSOqWVTy1ulNCwebIw/Ru8pyvTlJB
z8mT5Thpc9a4T+cehM03NJQXOLisceBzjL9f2JyExOY8Ba4/b3oZY7MlkDgnbmJZY1ajcf6nPUj/
ffKhq6vIrv8kQRiJMCcFh4zjUd2bC8vtjFcaFCag+AY6JUngdWTzj3wk6MBxIcgYqjCM7tUvAaVd
cH1v3vQ+aYL4w9x+mphLLF4K4/AGH+hrFudBkHnaJpPYWPd4JJnXhcMaAMGe5GqU6jbAAigwniQ7
Xd833cc6nA6JVMi77DT99LmZ8Wrwp7URMAjK11YLRtSjZs4ZcvxwHlOTT68inXhx8bjT6a224EDa
Wf9AXBnL6p/I2HL5jzfDYfEBiifr9XOEce/VGyIOC36JYp2WPgj1VX89Fj/kblww3XTjSzRw5WQ0
wrRP7FQaLf1z3NLWHcEPmbipxBEvcgpsBChpNoQpZ/QoZ9ROvwDG+0e21o0z/XcJHf6sZ9VWJEYK
wjeDymwdxwdTWGcmMz15hvcg7YaRkw79uwufBSQ/kVLrhcAvScW3KprAfpj4GvTZ+UccP3qj9L+U
Tg7Huai9qUftYM0ovaklI+0uGZLG5HyrgexdzDXwNMXFyCM2lEMxE4zAFvDWAlppmY9dMoVwrVGz
LxvUbLUMBJ9UdycPqUrE2WPsoxGRRuvRAIi4ShBLt5u8JVUIYNtAZa3iaR0Ikl5BPfF8Vhs6rS4j
gv55bf51y8YvsMTSMQfEspxnqHHOWwSy0NtLtPX6PQYL5z1nQYKmXKaCCGQBomuYWKwmTwLlxcm2
YFoe1rLCUNS4zzLEepSmiaVCZ6KrfRqfGdHkFmz248kDeCqHbZCL7ImscX5JQECZ2+dblW+gkSTx
ITx+bQSEh0bitt/KC8ew8sysRn5U2uinkg8vp8zMrSHjo0vwkoSMIlp1mJbjFIJWL2T//XouP4u+
pulNGu/iX4wZ1rICX5o57jyTvPcf/xZ/7CEbYCsTBUdc6AAbdiRAoIS+GrQ8CxNW5FQT8nFV+9v0
1hcpz2ZaAQjdDyBgBbJ0X2UjynB98zqcl7IZDKO/N2JNl9iHT5p0tjBimRDi7o/UAl/5OJQMhkJa
nQhFQEx/JpPxBr1jpiIdIl0griG/kGbERA7ZkYI0JVXVpMtVLCXeT8BthoI24I45IvgKMuKKXMJo
q3WQxmdv1ag5qNEsjXul4dOFuucseIXO1uOY5Xwgxdc/CXNC2uPK3G+JrMvZvVh77mcjMnJRM0HH
FOupi23g6JeF5yPQ97Da5GoO5bk0WK+ataSzRGJ3ABmW/2Wvg0DpsKaYTfZ53IJqXy8X9Toj/a6O
UgaCgksCkivVCs9CIUPQabcYTnKEdLsEpgIezHBoDnlaBuIlgNlGtFH2E98h/rihyrj8gJ3SfFdX
y+tBn4wZjio5ZSll1ftcEt7V4Aer+yIyCixptFLjI+60b8OvdiN5+pwDexdFNy1TJdxkvUpRJPbB
KpLMWhe4zDLqOC7azbUNsoSq42SgNbTl4KpJdXJedfBtMPiNrIpglUMJYaFPVZheehCP4ezFLtzQ
USGUjo4irThHrl4FA1Xi+Ib29RE4JodPdIZVvH/68tzCInNKkshRYmqXPATKfcP/AKY43Wm/bvKX
vjCI8TnrF1kRGaIhmUaVA74JsdxxmVY7Rio4Cbv99A0sXh/BpG7sClqgOve2EC81A0JFO8nLUECF
obUxXhj25D7qxwCxy1XaSYlI7kJaFPWwFcZeG3PfDYAHQUyA1qqQImKtsi/QTwwZPEkHkSrTMDUQ
1fiGcuozZnOBG/iiWOcfavvmwX1sXbfnv25oYp3yDsBjI1YjXkaf1g+PdjcKhBEZqyszRq+G268c
Z8SkibY9bSO3Ir8XrdPcvHpIlqtOg2NGIiPmfC8Ak/tVAarwg5uWO5ZpwsFgfQ5/BYTpMMYbXuF8
CjkFyWCEFzbi3XIwpmPFovTNx2SsY6SmqFcL4QR3RMb/nbV9I3b7PbB9Zx31chujJhBaL+z/fyO0
gfHSC+3DnRDerLzouG5IGbgtchjOGdDB8Igo26hm2jGjIpmXQanYy9ObY3TPmNtkkr+W12wTQCb9
trBSnzyBIQxD91dy05M8/4XVq+GLIoYyLL/CoJEcKUnfiI4Y1bxQlZq+MfV+xyc04ZI9MMAcczEb
hjOkBn8FYLhEjQiUbKnFMbvxy9R4dK/75BUM6VVaTB99iWmpJZe5jhink6Y/9RA3cYf47kR1hGan
ieeViMHkPYkaKoPpJzFIp7F/nvRMryhMA1slZDsPM81rOHUeShgLEcZpRk4r5e73tbSlx4pOFgYx
G4unrXDsyOBL4+FcS7wd3rzl08OBoB2jdlbrlmuhSjaNebzN3meDVFEX12Ze3GrSNdK3BE1ezyes
gnmuxyNZMU1Q2agcr+r2N3h2vtZTlU+d4yiKm6ZOwS3quKMpSRNNLo5ospYQG2YjI4g+1ss8M+Oi
Sdo/ivh7NNtzdqbnr/Cl3NSvKALUUvNkPvHCHyMo/Ph307HnntYQDZfzU1Ep2e62jOS6FkkHbPjp
+FBRJtOW5shwp4xg0eIhzIVUD6nQmPjwd6620EI/vAaTO/NZkEAsXjUyF+xaDNam0nmQgocVokRc
f+LMYcvBMaqhaN+AUL7a/Ko6LfR3sKEeFhvGWLk0WDXoyasOxbTcqVvagF+Opn6hVfeq9DLu1hHk
2a1LwaWeeuP67loksKgeTEDbmG8agfDx2/ieWj80gTZiDMOyXeVr9bN9b+iNFhr2L8yCaQkJxNNy
Ijq+Ou0G56WupeM8uRGRDJCZO5zf7wTf6l//UWmLWbAuuXTVrPCSWDmlO2l33l5u8cBHZR5B8rzE
V4GuPmva0VhEYx+x3YOwGonGgB4EUItH83WkFxmOo/XRlTmdwlpY/ozgVRpXj/Kwb7u47Y6q0pvh
4H72iKZVEXz+KW3uRyZfJaWbEAqGu+fnzhuwpcihx3ki2IuYXQJybZflHwIPistEC3g47KxbHoez
KJIc7RdkB7Abp4gyL+/jmaiub9dSofWdzO6UJwH2C/UWXmBJznHYs5OsdCPwHLho0zUjzt1L4qXR
ybiL8X6ddTFkOgTCKwAdbcBAOvneldz7bhH3IzeHkcjetZt8W2VeDjIfccgz6+qQMmmvOi5+IAU6
mBurLb1mZdPEF9s6AYyYQ8z7JAmUcvCDNLN8WTLwBRJYt4VBdVMxu2G7bFfh0EG+eTGzpuzhWVsD
GEcEfNWMrdMa/fn7njNwW1XWLE6QaTdtPDrq8brtJ1c11N265FqK6fTUQorNbx7ka57O7pGFSWJI
IQ3kCqEzcqO7lgwhSq3LVJ5s27ldhM6gHnAd9WgLovL3jMmgpArqS1oB5I+/EviNLX8SBqifqvuU
g/fd/5Trrj1/gkXp75JwTq2/21B29kB0GMa14xY9+Ylbq51DYPH+zVWlyUM76B/dF5vZS4Gu+cIh
A9wiey0DwXiJoZIhjgYi8Kmp4H+Df5xBZs/DKFhodvMsnDpi64M1NB1oNgxWgzIqHVipS+uhIHOy
3tsn6WwOwom4JkI0DGRfdOyiEZvVE5zpdANq5NfZDQATKpD90vBgMxAxEB8TvRwAb6/5nyTYyGHU
ERCfHQpZwH/t3fWwuaIe+afezyMM2nPreeIG7TCGo7ehWJ64s8BQadfEGlH+eBPZWiPlxpbSxg25
lczFMYpTt2iq7YwotvDRfebJY0nipp+kFaZVdAI91UiHlGQEV7yDzo0hKm+64leMJApIOAzQgp6w
24eTwCjjdfJpyvDnAuvKKZM3AIEVtLa4s1ZtwHQYm611L4xAP+HNZovT/KkYF73tr6FxM9TtIGZm
VED2ihe0npfLvYmXRCtIs/0FJd35YASaN2IRrTdgu0IplNbwvKUhNluXUmPLRN7+509NR5CJWhS0
aEsrqfA2g77b1kB0HtNXxL4a8mfsF9NWHKmd94eUAFUueHHS6AgQ/cLvgMZ3KJk/h6ZRQUJBfZ4P
UJInAZSD06CoPBW0WdFYMiqzAGsh9uxYDjAM91IVcQRdRNL7bKFjsVgnAIfQJyLeTO/3l6EiQo9g
XP/OZ4EtruaZui0OKl8Wnv2H2adrV8Wlmy37nKBJIT7xW/uTyhxfEeWd+trJw4lVRZg20sNSqCdj
OWStYcjS6gTQ+bmX33y1atWrhH/NSUMLjo+7vizvmGZgRsJBOuIht8RpdCsZiuz94iDKOqLzG3Oe
UG6De9OmHF6QV9uW/TeEbosJSHMvWFJic+1eJNUpyiArf5LY6xmMM3Mkcrwd74cfXK+/589ALhtB
U/qx2af80Ux8pWV1TqZW+LcvudZ8Cj72aNDSuGEmdnF+4aT3l07+OaykfX3bEXuwtsRcCDlBkgoi
aXhQOYl1osV1rFjjocW6ZGjGcn8nwOt9KPCA59ifBYwg9rA7735iCreCJRjwAtw9XHbHZq74mHZy
EDBtY719ch1jVfYiSxqwnw9lih6DUnGiR0Ft2P0Pj73gD/KNeM1/zgfKWAuz0xAUl28KIY6UUMXu
zZRyY1UyAvYcnf0m5ui3oQ1GXfAlVpRmPWF+XMvr6RH3iQMKA3IYyukuz8gpwRkaPqp91zXvFPkw
eOFszlKWBejgThPTyEC51NAiAv27QI7Jzm47N0bkOJ5rElS7aaJGVEmZyk9gxPg76x1/6oEdaOWv
b96MYP+hQIbWc/cTEVo9k8CWgrR9pBftuVpahZAeNu/fzVEcHASQLFA9wGu4XN7nALX1XJm7EpVp
isQD+gc+Oi47HnmPYDWLmzbiv1um9ySa2zw19C8kW9X+YKtsuQ8gvTDbJXanmpvVXl+yBb1fJKCa
+Mcg/3O/ZGgNha31R/Y0MDSLAJyOogIylrtNZGUDhr0EPgO45KMXX5HejZyo6ujyOdb8uoLzsWlQ
sVUi/kmr6MGXKfBlTowKFUGM+W0g99G2Y7VBQM1YONfz5TUb1d8c73zvuyqGlDtxyKaNtQbezwxR
2obbs9JKqkXCRN86lzpiHobeWxvRBYgirGz+ex3fpDbrv+FrQh0A7pOjulNkHcxaRBAbBWnbBG/o
WbxSP5h+cVSFipdTcF+Pmb39BGhTnnvvAz+kA1aKvc53DUwiBCZUnXzHhvT3+bkGUSOkQnQALvFf
FqYqv+MU73t3xtS6tFf8nkqghu+UE0shAnhoSNL6QGOcfzcGo13wnw6tJNZfcoJ7hKIoICVlloUb
ERKLLAwIgyXyOJONcQepnDfenVBjTFwTATL6DxnegNkReJO7oOp5cyFKFI1LCzvIBBa4dHn4buLc
asz5Hg9h8CEpkpo/9keeLTVsC/yVCRAhDHY0KWxSNsAjeW9MJ05081bVW3bNnr0hNbK1bMJntLaV
VePhRSS22BsuCOGG3GYUTX/ZDxnB0GGcSzhrg/5eBQ2x8QdjWv9lZLd+8wqSO8+wpWlS3kbIpTZN
+1BjJz3dwYSgnEUR0LRWStceWpyMOl+ThvYafUZP5pi5EXUFbEiCL48i4dLq7Zg7k5NMylPYIAi7
JLnhkMFx2fdvEHKQA0bLw2XgnufrSbZ5yzr5kWFE9AAmGA2SEYiUINj6knpX3TgrcCpPXHrzc0R0
icehNe8FUYByw6LD9CYdKH18Qdc2I5yn2MsfS20dskdA39qQW2E8QWTbyADjsi561KndCLL02HQJ
EwBhM+PBJI1AfDZGvVPTsel3Eob3KlKVeFYKkeeC5kpDYloDNN3yrGPaiILtCJ2OOB1DrMAcLsyr
qd1qRCsBXEGBFsLIDs1Q9tOLxiQhj3IIPy1GEuw7G1GyJzmNhAtjgtZMFENh3bLuPZv6ZHRV6fCN
h+9EoR/qRYlGWHc6FZW47OSQLxMSigJ4Ht92inS/eM1A2UNCSpGHGobpM392hQuYO7D/+GCGcxE4
RNhL636UGQDoVSVn6+cW0AeB44sDP/Aj0pKdTzLHZYE+0E02xTXv2n994p5sfFOsZ+NMZcmtfTY/
+r3FihGr/N4zUlxLAtE/xrQW8I2Vf0rjxqXznmiN7lC3j4cgo3Jb6PjComk/X1ebUB6H0EiAw+q2
EyVcPXLTiVqqcjYiQ2hVx0MvKhaIn2sfmLXiBO5CLZuL7Iz/1TdHiq/ITgYDEIg9Vurrj5xiAofZ
oo9aTP85x5h4znLUJL04tMYbhaXLpK9NCo/AXR/VzaJvQj8fu5+V2cPuLFsQ/gMJeJBD2IVupKrz
Pj+G4mXLYl5ydeqIV/3zrrdypYAdKVfTmvGrtGzto7wFkSO1VYDZavm7zZvUY2x87t8QiNtEqdY8
Ellu+hs1Hx8fWDF1DeV/t1XcV0wGlP+dxQLRzC5OS1b0VSAikpdyXIUhQzh26ogi6inv6JqzACHp
fcgM5lMn925bl7gZWyMWVUadaPIQvYVek35/x9kPNBX1SACpNRQeIe6libTOoc69fUK9lcNky4Eq
tUrhAOy5+d1rQnD4Rj9k8rX36polx0VU/VmRoQdthJ/KPwZWoMpcZBllwW2rzd6j3+MKyqbv5BGB
HfCJsXozmt2HnLNW/9yPCURbqBDsul7IWKiwOh4cZlld8HkeJ6o/+IAYhfL0m/qLMW12RSxR8fMg
nlrviJMC9Ypej3daTUkd1vgbB7A7g9cg1mt0wns/LN41YUkaYzuFLIKFcaiptgyif1Ia7S3n84Ej
lx6UIxOVMc0OUWG2lJzAqNSB9e5PVv3F7obpbVglPT6HSF+QIlqcsgs/YX9vIFHEpDvfALocd5nE
1p/e4/wnflvG5nrW1vF0XZJrfttB+VpUg5k5JuqkAx2k29IoJjxMZmY9vW3vDEoBNSopKXs060bf
rpA5TUEprC7BemZl5nSdVKiSEGQh17AnVTbUZpdtfbp58MqIxr+02rGjGFrz09b20veoAk4bPhJ5
pOJjFtdUYOt05zmnxgz9TfJWU8NN1MvWMp+koAiSWXUrcGG/QUgQ1kHEfYbmT7WN5k9nJ9gZJPjc
2u2xgcD5wUDHXzvkc6iGsf/twuDZSnK1c7o8CIsoF4ORbL8364GgUvh97RykielbI6QoR2cLDY+H
NPJRZBJeLem6A64x95KgaefMu+Oi6ScLewppEKHnXAEyK04JVk1P3TKn5/+7hE40+v/3Ig8EYUku
XV2iHhVw4DWMfr4+FUQnjRtit0otc7WHZsLid1r3b+ZzKwH73UuCPD8SGv37X7YDgWCLjZfb+Wm2
ydSAV/gM2QyQAGd3Rt0vdR7/tFu4tPxAlHk0BOm0a25UL9sLH4LZabDKPCf3Rys08anGA79ot/hY
uvj87oDHEVtCiEho72Xr/k8J09uue/j/hzbwuSJv9tn9GJxe22t1LnzYTzL7MSgF0CtDzLMtcByy
O73lOjcBcY2C4IByGq1jEPRWNMdpgnCLLr3gVB7SW68pWOZ3PeUF5Dp6dVEAGUATnNORaJmkk6Gr
nGS8RLD/sOGdrO5XLSTtejplJxibsMeSwB/Jqypzt8ihJXeICtVK9TOydRLMTlAHGVKUGreYYJKJ
tG/s35eI5JWChULHAvCiryPbeXdfYHDztJBrDZ1AfZz/+tH4CxyIGQTFSkFx7dTRZKiwLduClZtV
iqw2cdYltpzUWFwPNfx+XgSzPsPvwvc8+KdgIjgEy9gLwpNUiaqezbiroqtBhJPCpzXjqGf4Gqeg
Gu0aP3yV5557dlKbxkQqVHcPmDZEAc8z+BwPOPmpAkva14OBxV8Jd6/40pP5olV1FEcwsjkZ49vw
K2hoTuFpEYN2MRXoo5PxPghk4xsOgwZZDK+gR6hLFMq6Bd42b05ZBHC00uhzZuSGrYqp9M2PwLcs
VLW5nkWsekfpn9rF1tHpALS47FcspJ2q1KyxZIOrKYUot7WUna824krEPjZ9EuGTbyxE7FvxQ4YC
IuTqBdX/3bl7RyA8BZf2Mf/2uVVRm9N6hdP8B/QcD6vjQo1LKCB1gsokcjeYL1gGmqW171Z6Q0u2
2OjV/VrIk90wec4vCWrZu1elvAcBiXKWS5yS54qrg9uxDWnhnrN73kiScPtrTZrZyJTWdZ22wgRA
qY94NXb3Llh4Nf83VmPD2EaEFIPklCKaU2g//UldC2vB1cT4WBEZ7I/mQY/gydwdFBWLy/rxXt5Z
AWx3YgmbKqEcJu7YryipJYwjj+xM6bsVKLUo1sef8T1Znz/KVeJmQI5ABKdrdTV4/ujUGMRgUIqw
RPa4c1VCNr5M9JeLIO/gas/4Q/M57Wi4L+k+GdFjRgji+sHdW6/Wt16QT0YFQ+6u03asYlKydadw
BDrljJ7IDckRHA7g0u9HRvsaeXty8WB/UT/J5DzKiich000TlSRTbfthZPsquobxD/AjPR/HkxNh
j4JfkHZY/0bFeIbDfhzIkThRg0UprXYse0TJgrvLQGCZztSgO+HACsQZ7iI7bVtZ/FrXelnu+2WC
NyNLwLvHrIvUPdJ2FO7NdhzJW15n/DZsZMZahRwgQDMo9UQ8wej0Lr4isYzooHJMYk2B2VwhZpel
YFNikt+cDSkOFX8wRLYuMgATR8GP7inbu92OBf6mVlIdS7SqQxfXp36BR+RVRzRjYCh/lu9d1rJL
bcelEEdQN6vB9mS1uDp8h1fH/p1rGSKvw+QrsmNvCY3UHRK2wzUXHZlQSQ1tbrf38aivUhe2Q1dZ
PdPD4WzggWGwvmaOWp9ZCgUz4oZ4sz0KAgDQAN6U/71m8aeMzKhQO8mFW8ZSyrgbc1lInwCMXyTY
YDAzVQl7FhkneIJyKw3WmnecOJ4ttPZ0qLuXyK6yi2wAAYMVZkPiUIvFsizW+E90JErWqSWLPNSn
AEV10S/NHznqxScA7VwoOdw69SY+SWXjSkdGiJDze8VJ44Yo1mhHHAWaPHM7fly6D6k8qxaf+A58
+Sw4+6IsOwkLivUqE9cpwTdncrXUg1lUbwoKkgjYagKfCp62uPdqB+75Dlp13IY8fXlnRN1L7XHM
yv05+QEsk2YkmO95ZNal4F3EuK5rBDv/pPAt/LVRluYbzh2X3084LebNQMwtI8+W/Ped88YLzOqA
CkwLqSKWn5jprCjH5zdGgTfne/nigwyqtN3lVA06B5U2vg/rORAB5GqhAPq2sy+Zjko/VL36ZnnB
AIbWZwajxhdjA75qopUfFxabYy9gJsqnL6MSUWvyGxT7J64S5KtSOVTI9UpZdFjuJKjx7dHmMmW5
isjPNUFADgtTOtdcjpO7Y72nRuJ5t0a78akF0LVO4R9bE68X7yCsBJiq0eaQhFHlKMtMVpJKL/0S
F1mP9cl/PMBkZETCp/dt+LdsjsUuC5f+/OpiS1kwHAwpcYta1UPe6Ck4ynKkcJ9NPtD9V5enDV/q
IPIJrW6bQfhpLhGqiaL16nXYDTztZw9ZjN/tDhSSczYURtFYoMSzspfojz4fZDjhIwLOy3/taGce
ng8NN/rXWN/RtlMdpuUFDOiy77qXUUWS2Aoy5apB0FgE9N/LbPM2rWExejrxFZ60Xs3mvzOpup4t
mu+8W2RtD5hnAAf9syOlL77yWP3bmAPfm0OoZ3PtHiQ/3RZCzaPaPk6FXHecKR7dk7nm7mJL8iaA
BlUO7czDb2TZLK3rIkyaM59TKIxeL6I80GOJsm2atMuxCEqCF2LK+wo2Zxw3r3tNKO07uvwriwZ8
riYbcxlYziJD9ElNWFgymHNO7srhYSIwJ/bJQZl0fSfppU/NsPC2o/owsYh81LAe34vACueZBaxV
hsAaOgIPcdO00eVd2zypcktc+slxnWdmqHvAgV28ofZnJuyr9T5axzfRMz24C2Zdn9+RCVtjSDZo
dHpoWMaNizwAGdRD4VgDTRFyQV2y5VllEmH+HZHtu59g1M2HR7PydpLWPizr7ohEx57bEhIsK7jW
283oDCmjsKqhODnWGBN1s0HRNf8MHoOyzcCeLp6x+58CmzHEy4e5WL9/rPqRtrKt/24YI2Q4trBs
Ee1DJ8MS61OHS6VJRbTLGvn98SRmHudpud60jR9pxatuvj4uFHJGlJODrp8eNRujnBBkzoIE6BV9
4SBHHriatI46EomWPmJYOljjX7/UTg1dw2bUn0VBi3FuHf67S/79yHb4KGjl6R5gh5/fzPmmzlvD
Raxsthp32Jp8gQjSXJwtVPipltraoaAQEGLXwQpnHI1EMZ0V+Ma8CEFTREBlEQvlOmEylKyM5ij4
vQHhe3ntcN9AUcWhHDWGQ5hpwXC78B58lvAkODQWyO8tXYLV9wWQvSiJkx9XnNj/XkNz9Wp6AJ87
PcUDXWeg2P6coOK50ZYhIuIXyAaQ4c6zOKroDm+MG6ZcK7JdCMYppyLaFbaO3RIiKK5yqJ8A3yXR
a6cpYumA8teL2FY53JUK1Q26tJ2mflcYBOPGNHf5ZUbtgeRPG7gx7qPIvqTjVNLYIC4X8TFMcoQx
XFiwHnzMEmLKGZcp696TrQZ8dQVFSzRkfj4DQEYSd32Vqs6mIBpKmcVU/oduu8X4/z0Mnh2gFB7Q
4oCDaUQQtWU6prtUnYceCg4UBDTUIVrwKR30Gw7Z2UihdC9uOLkhbeGXGocVgA0FvmkrLBTWqg/G
+rEAwVcn8jvuG/Qva9xemjEgI5/B3M1n6gEBpIW/ZUMzu1lRNqD41zd1B3nuZ+HO82dnRugsFQJK
KTXWR90ZbNyRqrlutt2jBmLws8fp1t4j44L7oPw5LomRRSD9p+PZ/RLo/AlP8FgFOxLKlLfTdvVo
LEqaGREgeQiyTMm0vhk8l0YGDggm/OaHWRolnulYcy47+TyZL6KcoXmSxzR0rrY/MAi3rjSDk15e
nAdHZORjNJuCC+kQac7qR8yK7tY7cw2upQUQl3UwrMQ89JztE/vYdsbDgVEPUPl0IjMsbJy55Xlx
o3SAVZjsH/s4QOAuA02YHk7e37b5hJBhx7V0fucDzH9VxhNsUFF/OdVG+WKyzQZfZoBKejRqWNPY
FJisDWPzIVxxVMbPuIRu2QKeX5S3DhYQTYqKDpsuVsjbnC5+7hMx8zZun6g1wJEU5MtsahsvknP0
/42KzTUs4TxMps7fzzlALdfcQ3QZgnCIGBG1RwIfbi/IzdTjudH0J1Md8R1xixg3Sqy8M7YMOgUJ
2oLG6aiEkz5LuDOhrnMJAVuWZtOfNLSlU/3dQpH8MSjVlFi2b0JrcQvwZtm+aig4ATJA+XDKsfuj
HPxSI4nvbl/F6EeIptlcXTjrautnoNs0d5edDeAmwZKHhjI0gGotgckxfh2GbWeJIBWSfYb8ax5X
xIl9fGNECMNcKdELpF50np46odpuvKOQ1Nc5k2LVueTDaj2bNQ/swrcmNOjMNl0WM/dIMKnkyxOz
7g2/3JFRrmaU2ZwGgHgTRQfY1ep8DtpfQCNhHvHMwz/cnoU8rItqTiPkQLzAh2gtN1sorsiGsL3d
e8I8zN0NvvuqyCarnQZmr66g5YbHIldyTMRB/qYLLWAsA82h3tmnlX+6r7CzR2uG66Xtwaf9lRqN
SoEGmf2icHdxDbG4ek/6QyMq1mswBL6vgtVjRU7zqQWFNMTChyQGfkV4ArboAUYmTQGO23VN/RMO
zp2CMi9gu+MewLJawAl6CDmWa1zbnl776RSNbRYXMb4FMUx1CbwFGFkaEJ5RsnCD/e1reVb8/qzK
h7Pp/zzm7HRWF6BpDRDXBy2JE6nQZgCBsYjrk1tSySRT9mcoySWktDcsF3A7u08fdi88ubkwY3mD
Mvc8GLxam9Sh9HP5WWwvu5yrhT4D3W8Qh9PMa+6fIqJNXWUjBVJot9kDOUN0XxSLZRCm5/LQ3nxG
z4aMqyhDArwj3qB/08fC2kWNBqC7WAdTkOepcHOCWHqewTijgm+q5xOtXUuQhKUDFNSfGVV6UKFA
w1/GXwNohJCmtsRQqj6kqCB7W/vRIyvxPw+dBkmlPismPhMRlBSymQpteQz8B2xQPKfIgD3645KX
O6rkIyACUJMpth/xDENkZq0bg3+WgGgTGbFIA4U8VJeq5oobqmifExkdsa4LbySJFMMtZd8q6Mo5
l86Z8Z9wKp/vtFJ5cmEiVAJ+KfR4zHrBbZrFoXitDpKeIuOH55ahQfHgO8ZL2ij6LnK5OST3Q+gq
gRWwYpMbS1eHSRF5Dwn0Pj9FsBUNSqV6FtkzUL1uSOMisOq1HtGxHl833/ZnHOC7YFOsPRTsP4Lu
tZ854hYq6m9tz2scp8ffabD11gRVWkhTHa9ywKchow4rCqKbCLeWLZXvbJWO42cnAKm7YwFu+Jme
W5bbM4WhMNbRCYXiXNNGcYUA/EGVQeSUndv1gGwOGFbbYDIzQCDoPmmnicmT992PNtlU4NP787tp
kbXuaJnki90o7onTc3plpizZyNMnIY0KBhKh2Vubgv3ZVX0l97qynsBRh8MIJskok0t3GR2CJsOY
KowYeDQ1t4biroKQSHVvSJEJseGIX2NKLO4zNzCNOwhAmoe5ZbEJJaxHezx86k3NNL2T7wD+Fylf
Vdihcc2hu9vEr8KWD8GS3p4HGIjhTKFxAk/A1RS0Alkpb+9Z7IZmRNiFtqPMTytk+bV6vHWwzUUx
TJjHwX9YRDzS13dgsIiMyw4j7uIXuUwg20pRXvJIyCzMayZIqV3yEi4uAMyx94OFlC79i1ar6ilV
tk7nodrDYcDcv9Ai9yTEaCHLgh1N34bx0XgNocEH7qX/uJ3N2rR9pJnTqq+DIuxEVxDJ79tcUHtc
raBi9gStv3gBAbseaR6As0SuWwCSX7fthAAC/6fkXybf3XoJeixs1MQMw3zja+hxEl9TFxzwt26W
T0406js6R3M90Kl0hrwhFCu0KteSJDM+vLIRX8VJ9uw3+K8H3GAlXsph1bTyJD/F1tFOqqNGDrSa
8SwzPAAl1jBpoARzPFmy7DJb32/iK0OwS42AKSgFkRX//nnZ7uFtCbJ8X0SlIRHScgCII70OM1gd
cbqs8qb8ykUNmXOH3PzGhX0FWkJ/WsmNcI8DOvcHiZm/z+rq4nRFfRizRWzBj9OKFLSdGtyI0mho
we+NrDOa+3qNH7UnPXQIRpVjE7ptGGUXN6X6C4KY6hrg1xVnGb2XLzbz8lPFNpx66zHYmZU1KIjp
zDk9K2e8QhJAk9kupstwrbE8xTLTd4ENvSg8sd7z9bHSgiAWSYLq50XGF12yETvwZ16Oa4ZTQcJg
od/DFYvvi0TYMQXWLNuBcdQOIi80WYpJG8LIV8cgp5xaDMP4S2rhXwmfAvzQkvG+n6b21LCWhfDD
bfJEyUiRPmZj83kz59TM5hFpY/cXJlod+KQwhDSlaOaNUw30hl4XqqcZuHWzYwkDvYyrbSBinkTC
llIGl5kDtPiY8mV34fS/4p8OEUXYhyIbVPqhayqHYWBNtfDcTmQo1ZADWuspnVk2B8bcY/XVPBzJ
uvcvORxMPJr/SQgO1kk8VbAI+i2OF2uHxD+0cNhONPq4pMFSpNpiMWKi6+sjGWaIGwuqNiReZkAy
qKsTiTUL8obWSmldRojAPcQdeqqs1p9aVL9AHIu27Tz2FsiEvyG05c5AK6e7LCWCodmP6rzr4Iuy
wMOLyWY9dPs7ENYFiwoXxGP4VqK3q3USHKFgyaJ4M/LN+mpj0QZxfgrAyEexJ/QN2Un/ShgaJ2T+
KfScOuGbHJy12luTCYOYBU3NvOZWSvPpRhipAkWqvSPzrBNDp7sv932mRyDEt4GpBuZQSzuTd0R/
VA0Kb7wUdxa4NtZ4ZGXAcGf17RsStUgBLdVpSO8zLX8BfjClnXy2GvNMqZLygAGZmZ8fkkwaoaWP
PLVH22YD8lvxu73Fwe17hHVKoalIDB8mw1UbKztx1bSMgTeU1oP+W/57nnw+ohQMciFB1cXMa2Dj
JKrIWbcNMpC+aAKrkxkDGMU0WZBzLySiiQB1nntweLsk/oqizHUm2YUVqCB0PNN/jPQSFAQJw+J0
U16hspH4iNfSi0XWbD2Enh4r3SEd+uUg9gVWFwBGOpM0HELNt7dS07zLTbNeH2JeyOLQ4+pvX+ZS
YOHxMy/1EmHZf3D5exAxDf6nk7tVP6BSSamg5j/XQU4R7AjDD//dnBi2Pi60B34JkRUWMKE1rz0X
Tuc2F6lAt8XiJCzw98J45hp3EYXZcOUVOMfnl4vyDzt+vfLOdtQyxTzGZDLT+sbajb8y2ZUlqxNn
WrYiIGOdlYTrQdXsc/Xt7xJ+akO21cBeVUHyN2OzRTXIZ/CmlEwvBd8GgE9AtjowCPC/H7k6blpn
OQh+CtiuBLalK/5MuKH7WGZ7Anv9Kbw4RyP18b0ExehIKVKBaPkLEZPdapL0NM3K4amRbTqKwb1I
rsspu+0ZtGbdmo0ziX8dW5tsBu38cuP94J37aoUrv/Bfi0XFFVJp16cKPSlepLKLj3nmqgqor3jd
eRaBAVBOxU4o1LsHIXetDzNuwt8XZc4J71FRLq4TKKkab4ue5QA66FnNJ6oCOlAhMIomtNyM+U+l
Xw4ao168xYCdkQrvUb3g2cdEAeNmmt4yy5C+0p0njvh4yVJng40Hxmd5dCOEK1LqL3Aj5tsgpf9C
ypN+/DkjixZhZwG1Qk1Zddw9ta0/WoJtGs8zM8cxZqgi3bdR0N4BdVn/HUYedSXeocaZifihBWXt
+O1kL1lmkPCEFLyKxNso4lPXKHxxxsZg6woFvgIBLseKpTYNZHqYRWwaYaSVF8xqMjvsJB1WMhBG
d6DUBX9Q8v6oIXBA4XU/qLmdKzeiTEQ4nPiymWuC/McovLW/iBKMyMdql5YQ9xqiTD6qilocdbe8
HwNDjinmyvyv+aQwkeERma2/o7PzMa9HVizgyAZHi7TaRe7OFoowSYDzw6I6qtCpmgVWXmjKJUlq
nLALkzkzRC3ajB76mScs/Hhi3Y0eRIoOtoeb5iJFDuMD2+ZUZbJ2/ZHUVQLHNBpI1GotuOnH9oMV
BCg+oAjejW3j8vh8nf/EsKOaDQKNcOHFwrLk6nsz+OxkchdExcTpeTlgI84nZMSaftEK201V/ia4
OTIhG6sHKPu7HC1B9iWWYXVnGdG0v8nAEpJhHtrRMnCCy47if+gxANWZsU2LkCsW8+JVC7P90f6v
vOHH3SBSDRiGAKS14d6BmErakI13VlS29899LNiBX4R8MKaYOZSqN2u0wBmFS7TxOiEuPjvG12Sl
rqZTe42XNmKg+h4+Sgg3wbOsXK4176J3pMyabO4o1lPp+tdr89EFJvT9UhEUwnKq53LklDhVt4w3
/1q1znosv+qPZjcqnz580GaHFFNHnRMjlHmLeBbqAD+YlaGjp5iL5kAw2BvPcjRaRp8Xjc9xRDa+
8SVTf6fn6nhmPQp3Ns7vInX3Ktl2hxvPUe0LxXojFDJeehbnUS25Gtr/vNcBcqBecTStGEP9bNTp
FBiXpPqmPiRj2dblgBB2q1XkDzqPbn9O+Kqrt6p02CLLS3zDTdXiRmeJH3z8TaFbj633DKgBh8Ct
f1d3y30w3jUtLBOlzS9e3Ehg+zNojYBUAlmYhxqxI9xmW4KlJISYhVClMbSZv71dA5+smlkNeZUV
cRRcDZdVKRvKTJy7Ia4dz382l6GiGg/ohYKPpzcTcm93VlJ6wraAy6/pkRC56BODZVWosZ4D+ApG
n4sb8iowRBCeiFameEDIbM9qUGrZbNuMFxOKrdpG1Olg4DMJr1LtRwkVkz6s4JTrPDWZ8Gt7hpPm
jxNMw2uB0YESAovhuXoaSBTuMLF9pFZhdFRS3Rc94djdA9H/k14syxm1ZTigSVsiYDtPMD2doZR/
bEZ10ClCg0D0oyTuQaZYHyJLzhBgWXyrOsKRJJoXc8jPLMK/t8pbfn6eQeXT3v10pYaT2we2ZeY2
bx2FKg4gimFtMFkQNQtjIlKCamgTjLgdba2pikMElJFyEKe7zXp2ncew2CuzuChBDfZubjYDtDCp
tpORy9GOk5pEyzhrOGDzZmq1RSPZR4uNwZRLPVRa04aoVxfh2UKa6n7yeLU/LqutOD8tC7f+yC0f
rykIzuzFEqBSKDZsEYcNYxuUb3KQONh+PncBXh94qwho4of8IgVIBASLYaXTe7punXBaM2EL59+T
audCGktgGHwMvduYjH435u0bo0dkWVad3KHnl66zcF6gDu/9M+5bteTsLceSdIP9+gOoFA2CmL9h
3qvAmsh93OygZOP/4udeVdd0KBwd/30m2MJX4GXHF3OxzuecfSRX4nhJihY+3krHHxMW9wb/1KYI
MkVqdUS6THOrXhvTMLB9UXU5DlDc345WnUOuzlA7f+F4lydromUxlZ3HI0c90iRq96WIOudv1JWa
y/FazLq9ZQHw2/xprlL/vTljJIYdRKiF5Am4jTeW3tL1L5v6b8XE3z8bq3FAPJF60lsctAfuJdrz
kbRCQHuCiUXgCo3hHb8rsPrcGAjy3lPm/Hq4JizhhzvhDx9LGSvc77x69IcpO+Qlpa6OuC8H2wSx
C25gXNDCVsE1a7tqKxlyVLLdYfWiMuQQ0L2e5fxwVin5poULyTI0V69D5dY9s0Ly6ALvxhCp6anu
bM2f5SiC1j7uNrGLn/3cHQuRxgN6JCH0FDROp3IWjO9BafwMBkewcxKnNJle5xjeztk9JnehwPVd
eJddumLixIMfd+6Xj2fxYUxq16gm2VIB1NXv6Wgh6g9ZbTP/UAzNlVdaadbQaD/a0ybxQh4luJ+M
NF7vcplTdt+r7l5ChLqPY9zDD97/t9bZmR8kE0BsC9YExw/zPoS06HmjewN43/gQPer50Uv4CKED
OaP5/u1D4C9UbxsMnhQFS12kXOAXEAsDeLGZOvuqu9a6PIcAPOiwzQaERiHsgktBOxTP0jT3bvcB
DO2C4mRXuTdlhXUjIJrnhvY5682DSogNT6yg1NXSho17W3I3OdPu/VyP51rvm0WygOoTUITow3Kx
/4ZpNS8t0BPusbY/2uzxyoiRnkMBofje3OB3gt+Nx2CMbY7b2kvloZwb8Kk3ZGyR+wq51lIR8tKg
TISc30cm4+i4Um5kbgVklp0zPubEdRLFdWVopO6d9V86aWzc91d+idhqgA2F/ExtIQxjJP7gLnbK
zbG8xwx5vsSgBOsDzkz1KWvYrmiuR20ILGB0K59k1pCMR/4FsHFhG4ijAROdCfVh3SikIH/ova5L
KmW8g+P4G8w29BZuQR1Kfajv2NSYgdnrpwi24P/BcUX++/7191LEBRrux9kh9OgWX9gFEr50XiII
qlcJI+TU7WwW616ln0tdPtWh3z8tpaGajHVOMsju1GrbU9dqdC0oLhuJAyF1YkP71SrBhiO1/ASs
3zT6+7MbrYSBqncTJQWOWLTy7pz5EdqBr8pZ5bhWo9P7IATcBXYKHnXBdzOX+7Ouo8k3Sb+lE2/J
UKWmw5iYYao/8HXoXBIqaa8P86e5Q8cIZa/j93hgE7cPLtxKN0CpHBcR5mfFWUHONUB3kAKFBY08
W+Dv1IBev4XRX02OIxRonh7J+163Gd8xrDt/V+Ky8BCFRv+/18Pa5piXS/nZA5pMWj+fmvF2VSuV
y51S8BLWDhzUNQhYVOc8+s9tcGcNsY8rmVPLNQhGHiw0UnPrBs9uKVCfU4lN43TU6UiykIOgkKl8
D8or6AnyYc7mHcyjGQPeU+KN+d3XPDwkmilkK9qFXHbkjlR7wXYTawHN9ECeCR/ByEe2yAizr0XU
kSxTi3JA3Lh/oVTkOKq0aqiNQ00DicyH6mYUE1K0cdM/WZDYM7fwm6x+kKYPP94yARN8/DZKLuJR
7j5dFThD6E/+dQc6Kzq6clbRL3ItOElvFvE7kr42939cphhniJLSaQha7yHI7JLYs1jGcPhCOjpf
NzaliboUNGOuGpCpnv6oK+xMzqb7vxa95cyQJEzN3D/+8iIxmODVYLTJMtvQ/sx+Wmjt5Ul66j9F
X1VeIGtoT5vRnRltwlSc6xAr1CjdWLFR/PooCUwOp/z2p4k0zKlLCho+UDUFOcQ6W44wlhCYWRWC
cLbLVp4NDvA/HbSb2x7xZ3phicEkLAhCOkERhiA9E5KXvuqQTFv1/2RqcgyI5146dDCM8fXKvyWJ
4knqBfA/nHYQPHKYZKW21qOOteT+m8TiBSgiGlrZN57Uzdd8ZNE3Hn9JLTzAp5wnihYiecLvavgs
UqdA/goMn1t1O3hDQfVpdFoMC6hI3vl2HuKc0XZJ6V+aPtm/V5C/5UXZpGMJtwHNLI7Cd9Ri6hdY
s85hUugRSxXlqmBMjjIgQQdvrlUH/cUg8yZYCFZKr3swccZ2Mjq6x95uM7XF3Egdcm5GKtx6Hpml
fvxHY2zDXuZVpHUUJqKHQkEFFp7I+Zs6XwHtYD3NrHJKFhfF9Tp0deDjTehu0zX4tjtnXrZhNDcH
V5XSepo3ToFG/oWGTkj9/Bf4piUH0PBSBs206R7HPVgg94YCWOf1d0MtllNdnw6x6IMFifulvyfd
ds08K1NTpedmTRhNrQ0SDbKcZhAXRHRq+kGVkdrv/e0m9Uxo2VU6n9VRYrwmenSOa2nFTKOYwSoZ
o9bvM9VnZEE2hwFrr6/b4OAwQOnvq/CmIfzzQIUCwHXbft5v/TTvGPBd0baeOaLcr/SRtMhBoEgR
8Gg0A3NVE93VqvLNnA1+qEPMOdWqFYp7PjW6hxGotcg57SISDZGmx4o7EtHKfgUxi8Q39sBkjL3h
XHnT84nQ6VmhdeMLyfMaamFuFROg8GNbuTzzmrWYdACvWDJa5eA8xBWuT6b/WpDN1WeWfaaEEpSt
D0Lqr8WxsONtn3oRjWHud9kHEg1PtgfRSkSPhz4JDFoj+pgz62bxdEaeyEQZqKXGRzAm0yqslB+N
bJda9RjzD1k2zZRMFehx9piXc50Jg5mwY6W2LkG7+9p26OwhZj01ZMtpHcQjPnb9Bf7MriByYxkb
YRH1Y7jiXcZiUrBno2ZHXETFlulpp7I3M5DIVcyHQeqqUh/TLqFZhOTOw45no9FXW7upGXj9HW5Y
QSNQ9TcGRkAQTTg0/AOI9d6cFrnCB/CpbRsl76fpVNfen2YmUf/FJEmKctznofqNm2K3Dbekd4/E
QTZItH8BWk//pEr1KtbQvyPeV44YqKgeNg5WkRkpCn9UmC7avcYGm6L9qxHZprNmwS0eW2PvRUV8
is5iPNhnwTn4H4TeTH7xjWW67YUXP3dBIHMWfl6N5yi70meJNXP0ymXY3gasXEljU8fr5tvGrXao
WL+DyuwOdD5Uxb7wW7KmkQPNw/eKmSeyNf1oapBPlEOraIZrtCNmYIZNnrp8tRBe01b+AB92F09R
apEWvh334yfzeG9OUg+jD+ja+SF5OMscwu1mHAwl6WeAasR2sO9rNi4e0SVY2loz5tPraDHRMTqf
ayeajZQXIDyMF4zt2WEquxpZXw30rRpFT827g7JoT8pqQOuT5C0aWNDhGQuj7MnSTjA9zLFVhfrf
RlcBS6VjFORxuO4XGFIn+UBv7P+wb5kJyUX866y4FWK/iHooS6PCej6VGjS6v02G95dFUJs2cyk9
kI6hZ8ulagxL0HSsZBZtJVtDR5AH5emG/qfXw8G2p/iLhvR4Us6bakTABXbFttEtzlNm33o+DAMb
D6mB0T3pCHdPNMi1XWnfZgVtROnrrGDbN8ieFATXc4ypValdNcfxlvA8VPtNqFAxAJnx9Y/W6aqO
lCQZBaTfIN7VKxg6ek/1zcAU3DuXPkUkDcrx7HoeD1k8lcM0hXweDOF3GyN6BcqunjvCk8vMS1BD
rR5OJQNAV9Aw5UgIz6VLHqpM41yzgO0fmR/Zu6ZT1uMVvbfpphc8+LaA4RAkqVfZF/KPHClP9SRy
IntHr7hTdRMp3lLQ5avO5kcwnu5NDA9zPy7nZtKwBuaE5ipn2s6Z2aAcAuWZDZTB59bq9ymBEWnw
ZVirWOr9vDP8vIAWPiYJLdTPJCcIYR6NEhHQnO1NCxsSLj4vHj0X4B5PFiaGX0nTk523itdgJyYl
Xhu2nXKnTyo6U1VNXNIa5naQiBsaMNWVmUgvToCIdCgHW3DLJIbx+5q+m1C6K/l9rEiSTalVC3Mf
vWWxZMNwTJoVHg5mok/ehvQG27xmT1nl2LPOjn6UBeqnmu/75inmkDaUaK4i8QCbzBeElEBxwAM9
R7RpwQjbc+iYA0XuCl6mkpRYUtd54RCzhEirDUnMRu6nXWzrdhTT7Jy1dlhjv0u3R4POY/SMwQ/8
Yq1p96/zZ/Ah3YN4Qo6nz3SHM8KGETctxqMieSNMBMAtgS6YszIhFRRl2UPID3VoDxQu8fzQmXei
B9m8NmjvaBNT2SR5J9WfTadktbQ4ipU/7MDtYRdyaW0H8qLWzJNo60Sd2ETz/Lq4jiLYyf3DHiKh
pDn1bU/x8d6WCW+w3RF3TDQA/9/RWYL8Ecll0/H2H4xsl2sV/WYIepvV0tVBYOEoy2byEiXkpCi6
z10V7iGvG2M4cfRGpLWOn1m9v3C9x54qOfp3Yng5uhEkfgEMV4Xo43CFNbrj0aSid356YiZjfp9/
JUfbR+E5w/Y7hK28erT9LwxWs1q94HWXtwT8cBLpLIrJgR9BVrFQ17UNuCo147LYJhvUHRV8Gk/q
dY5cn046nXP0wO/p8zQf80LeQXi/Xo2ulOHoXrHnIIiVlQhs66drDaitpUiK8O/fZ5MTeiRsL6Vg
4ve6MuHZJYhkUklmgwT3bgKmMsCW1aWzW+jMvgkumA6C5E/AtodcJk6wYXnYh5cIrcuwHkkCyRRw
dcnuqpA+j1sH47nK1oSwQDZFxxpqLapEy70NQGn2/tSAa5z9Tsp9lr55icSsO6mvnZkv/n9OWGjQ
SXVa2cT/D+5vTMbDUeywJ9QdQfAuyky0jM9v+FvKN/F4BIDsXz5BzHCJPn8a/feCrqqTgZoJLEGc
n/zgiJjJ5B3wNH2JGZV/1skZ4Uc++O6Is7m4Oo2DML0jdZ1JZ7tHsR5ky9yES7OqcxXV3fdukMDv
nFLmUDDB/Ut+uxkvi6y0dae4d2epyiEUlU2ZaOR5ykZcWync+/BwKfaXhc2EoRIyw+harAepHYqr
CwmzhCfAIRtE1XY1akOw2m+LnhS9MN5b/Wrx8pf6WE4fTVuSc3MrWC0BcE0y/en/cP0blKxb6+ej
vHDfAIXyxQ0wICKzUHUymVDQXIgsu5RO3k8gwtZAuWy7Dr9YV19QWPG1xh9A8z4kRVUyjLDqDY42
/VwwxJNIszjPdNwuNG4Ry6f9XQiyr80Vq3Kn0wk3RS6P2hsZ+oP/cfbEkh/4xcaJRw2N4jv05jbL
ERv1UqoKS3uRBYYEyO3EPE2iXNh/N+lVs/hniaX22iglfZ0STANvViU10HrjRoZGGQIwpkva8whn
00SnH9DJkwMzyvWjuNygLcG32Y0Hy7IYGj/SO5DHCJIg7Ad6cX+qiSgsPBGR8/+RSg0zvqzC80NN
Jy2l1iTq+y/J0jCFhabRH93cjKVL8PO1Gh6ba3GIlvUAFy4xmYsYwKapuynihYe+E7nNQRz26Ezj
/2kHxv/6e8NoO0Xm9+1Pdp3Ra9KXDTNEUG72dmPu6eNsN5cwAXqnRIgB207/vkMK1dXGRyVY7g79
HP6jm9q+/nQ87lY2hdUHaoE2ZLlawZO5TvvQX6PzGdABpPckglTbnYI0DNJWT09+kg2ynEc7CBVl
5ZHNEQHoJUaBmn4BTF5+SHMqchA6S6CjYZw8GAGH5zQVUN+/xUtVWL1F/qlAmhz4Znkh6kEHxthX
sQiSHoCdgsDnhXRKvCyathvvu1E9rg1WI73RcDe1x5ObNlplNqiEE41NY4c8R3eZ6PgpUfK/h3DS
2qUTWgp6xW2B5YU/cx7r8w7SWEVuByHXRt5o5NC4nM1RvD7LMlwtuKegZ9ccVLlMfAMWETPLh0XM
pmJAJWYX4q7eFHACsfOoJ1y/+9TpNDazFf5sDQkDnn9dFaW7B0TfyTF6q6h6f9XOv8Fw+gARULRS
5pqgaUMR8zztZ2qGbQnVu4EELZo2wimD7+ESQRS9L1LUgxUBd4PUyK9Z06QpSkLYYm6Jl2OD8vLp
bZ9cTEjd0aMNN1pgUJ/xxQimE6QuP6k4v0uaigzwR8uavZlWaybSl1ymXPfJU+3PU0YswjwC+0Mi
nhClH1WZUqxv3yW0kssE4p33JjL4vozTA/b3JFrMtUjMKEgGrkunxf+zLDE8Q2KMCb2zXJcXoWa1
b+JtVLuxwHQHVhlLeKMAi7eNeqaA+z6zsFOeaTKTCyv07xPcOgbABoKJa+eD/zoMvMQJt413maSY
NyKfHQqiyKQVlv4M1kk7ch6iuFf9S5BFye/0Fb0PsGzCnQfeqv+w3bNUKOORn+pNP3Ob6nZRX2YB
+d51oHmvCdtqZ4UpIZQVIB2lEBgJWg7ShuJ4PeEDeTzmv7Sk0EfbJdRbEd0MfBssRHoN4ovx/Vy7
Wa/ZQfT8YCYtuIU83XLOnW9z0eb1MRT8ro6BN/rPPWgdX+mjqouM+aFLxl+pGMZCNXJL36JFhARQ
pN47+1F9tqF5bCWO3RzWBuJbm5iDXs2mGc3VBWaVBvlT7HCeKRyXFWdgt6ZmQlVWMC1xfR36FhRl
ALM9wP7FZtqcx/yUC3eQZ3G/Gb5ieLCeYD1vKS+1lce147VqpO2KMIDcwLptfbxV/dbykgAy/F/r
wKOmuKgJQoun6CtAyPQgLypj58CurKj1cd8GGprBPrBLSb9wJhWWE3Js2QVCnZFI7yy8kMgfobIq
QRf2+Jimyrxwl160RlDqIBeAt7om0WgMbdo3a4+zer9Ii5m5o/h4/Kk9eW7fuIQSgbZqxZWpukgb
tpSHxEJrqqDmlB9JzyC8QNJhKF9Rl89xpBlyK2pl/nLFR99hnSRvQkU89A6LZOLv2KcxtsINkRGK
O2qXxbKvaKI1PX0zYIWI/VMz+ipEUpoNNl1W+ucLEL7FNx2O8gzkomysAwRasqUFLHGpzbhYz8s/
rXMeNHI/QWUB3ZmmONJviOulysEYHuNHXV2GWFlt1JuMACq7gC0iPH2208ECDQing9wIm6kLDlnz
jPRmeXZD3Nhf5gVbnPMSI0pBPblmv4TkzwvFRdgQrMejRI9uyvwnsVk3YuuKeONX8r5XwtaS2AbV
ICj1JwS79Q1YWiYfQwwR7W1M1F3zDhmH69KPdIrQFtwK9HRXyLEX2LxMVJr1kQwvt9Accv2ZgZ/T
SUaj6MxFgmyrxVcYCpvzmqvtThE+kPLpTfc8/evyOwKr4msfNz+EDihXKPbElUBuC+x9W9aIJMx3
S+30LgRrOjsRcfCm1y7IeGJy5Cyj4VN+O8924ThQviHEk6HNo6qptTp+K6JtUjpKoyu88J++V8sQ
VhMzeThwNya1CnDp74zt+M988XsYgOKNe+o6DMwO/GdodzQKPRDJfe6D5qBv3mXM0MP4eRAR2sRq
XRpegsozhneT+kSGXvydVv/WkkY+rOzjBHxwOHxxOctdm36QBrP3WPJtma2jjF+DIxgMYskO2hgo
bGq0/TjzzS3pKousWZJPBlnC7vrxy0J9L/588ybOFMxz+oE068kics1ktc8721JXS2SzW1XwU6VM
pvOLzKB+q+EyFueBNaQrfFBX2ouOurZvWgI/ysW2/YtxfSCYvXN99fG9Ge1IBe0KNclB9TTXB1MG
ezqjQlnYTD/OLpUlTY64TDtVFxvFDQCO6xg1LsGn/utSVmn7KaACg90jE3FM8fKuRyfQVeP6/YDH
8ZWwXsTUr3WpdJeQ50vHy9SagSOo+jhbX1q5H5u+6jOiDM5LFfvJ53oXb9CkcHSAt+Doz4ZU66Ut
WoRO1DSSSeD1tkVE3TEg0hZ+xmLv3W0S8M4dKnpwvHvrDpfnm+rSk5KCRt/0WxN6HzlPNOsudkpD
pNKumqPiKVzucYBNSmK8xaYzLYsWu3ZM07ZdsQ7hqXoCJYimzRoG5ebjibCotx1SXzmyDt+1FSLA
pAFqFeeaeP5592G1dCzCO+g+YQ8szlOwXt+96ahkY273s33UMoY4pDEVSxSTsQxNo2use/AwdeMk
aOy4rNAQzvjdPfQMh12HlHed5FO3RWeEdP47Oa/2RogUW4zstsyUnZhgOVtvywp6jcjjgeanh8uA
Zjao9HAdbm5MbDi/p2HwZyIyPxdeHT8jHmc4U8me2SP1J2T3VIPPsivzIKODfFumhcJCMRLTEIWa
EyfxymKVvanbn56RpyvUvAKq94H+1Z37CYHNAaT1v3JD/YmlaKd/9YE0v+MPneFJfGUSsn8t90pP
586mx4m7gyprkJ6GNqdKWIYMgqfPf2rqV60Ga+jLWTRwx79P0imJfzrjOYFIB7LTaKrCpljyG6Ws
ofITbirA0qB/7hczQ0TFiCwCR9KmD4w4k4wo9ONWz6HOeJEzm4jtgrs57FWzWWmW6oYqehaSa2AE
oBx2ZvL8PoI0e/bdvU+oLv1PR2EmZmkL9st/sIdquGGr31tmcYOr3pp+MKYGY0t8YoofdyDYXabC
FX9/FToo3uzjSTG57FE7OYQfMp1sA6s/+oSibv1nVYZzi/TZkKOjq0HqZ1h5QDdIE5Y7uMvuOmoo
+anCBsR9EUgna4MszneEV3we82UvsCZorjpj+eSCA3r4AC315XVAWm/cgfPwPK3B0g39nTeR4G+J
TRHJjPX8wGtdwOBnePZ9FlWgmBj667dAqy2Cqa7BZfQe/xtq0UR2pXXro8tbUwoZdUZA/EGQKBhS
HyMHo/Tf/erD1jHFYw4T92/feCOmsqIccCmBDIvuGtuTNaDqXxPswhlTC5cRUNerCrCCA6QsWLfb
At9DVm+9KG9FfTLHJKFvonl4hiqdYCy7uDtjcNMxhFqfiOxYjnmkHoCHO8pClj/7Nz605Lz/Vo8M
+t9fH4KOAnb1bC6yPsh/cFJorEfUsjui1TkOFC2Orni7zBmPJZo9wNAxpJ7d0x1LmPfTZ7SK8NiS
A/A/+e7mCvr4U75LdEaRCwOZOJQ+mG8MgHg9K9K1xcmHsB2mZ0Yu5QmMnNdKnBpcpoHOssYmdi1o
v4xalbEFblOTXO0zfWn0kifDOBhd11gWWuddukllJxiSuuXzV9umQSIxviomvJw3603TFr2Yypc1
6owvfX+h88rhWQlkLZ8eqJ+o6Y2iAHFiPtfm21VhRaOv1uhXrBtJ64Zw0oTCDQjYWIrP2AGwC/P2
FGt7HlHMFGtUoTF0d1reUYJf7hGx5BHHdYsuuqY80/REnNDPlK/gjxGFBR9ZToelEBdgi3qKMmt2
pT0eOMoe9dpS6rTRg09J5S9xgPNK+KM4WYS5UBhQ0VabPngbRay2LZuBxYUmAlxg3TqWKhcoKEAZ
+dVoy3D8gbhu4xjfRuVVYCYNo8D3zZ6G68+CC2B9aCfRXSonokV8KYDcJESzdRnOW2VJ0xj7q74Q
kCrlfsE1mY+mzBXpnbFosPRlcqeyauPHvnLgi3JKSOv/33FcyJ1YPJ1fmjOqSEg5XDXA1j0idxi5
7KUhD/MqDI4QiyrxC6A8EdlbHnmI+7rZ5JP2jq4p0cMbKEbFlR6/3MTEOKg67LgBhOPdQKgdslG4
WPV2L7E45BrAyOE1SVv0BfQy/bT0DXvMH8ljiH8Lsa2y+OtNnu7Xmk3DDwoKahucwdH5rJfKHaRu
XrG/GGOn5BRKKhXT/alFKe3HzjAtRJbiOtKAd+50iKnEAxUsI6zAO6Lyy3Zlcj+/LYsoowBxVNXi
UYDnOdixEX+E4cGto5AO7W0OTt9vm0Ci8e/EbCEZjqK3bxBqvIiDmk11zaVdvWCEFjExR4oaqsrK
nInnMuTeD/VLYXze8JS/AYKQy6P631iSorZv7EBYx47cUHkYZZvjQ7AtGI7nLaEws7D628IYQw+r
gIyQRKr5gIFRzzydOtaGFyIgj2tNgkmWkeZxyle7N9qG8vRIa5E9hfSST+0GQWitmB6SulXWk00N
DMG+4ihy8soU6AqOZrBLArJeMh0ytcFmFq57A/zegUwAHrNWX1h6dTThZNYBOjSmx9hOX6k8/gqm
Mb6jZofFzl5mr95oFdQWuOV+RMyQ6PPgxhaOQKvgbXzALuEqVeYgEeXCHH6qQ+KGMopiigd4ev2M
VlygvYi9As6jIu4WbGamWOVpkzUt9YAqtH9YVZq5p2CxSKGdZlEwvGeYKA3ay75BJGZjaJRaGjeL
i4m5qOkr14gx5hCzyRbhV/LGFpqcgUUBa9m/lVBI5HWhbTprI3RdnOkWpiqUK+vagUdUpRZxnCdI
erhshBHLY4Q9RMYhOgQ20EA60AjON2jnaaSqPDw2RDXwF+ZLiNk+PyaYDAB792Q5qAcpuO59q7QG
mJ5ZdIoBc0ElzuSXUNHCbOXmZRiPCBZnJJWpTC4f0ESb2N3hltw8zYxtpiB+fhD82S9wkBebTWlD
J7UxGwvY4OQKdgAEt9Mpv6WXHoyrLokWlh2CRrqRa6nMlzyLSBOKUuzIgtbsauteaauJ3ZETZkRo
0RUrIBIqiL7+eUnaFJ3cGvA4wIWhJqZCCWLhMrSres28exgu+xz4kcssT53nimiqfDY74ox7MpgE
Ulo9RAEGDC8nDkDytxjsZu4+B08DaDk2JZHqcoj8fRw5+7Prqg7KOPsHE80gld0AakAgh4Vg9IGb
+vFpdFC0kymPacLTrI0NX/uHCl85XTytYQUTnDE7Tml8o918eoc/8MCwGBL6Ii+Ukyv8Y/rcRcBo
pJU4PKWsGt/umP6yNIPEZTWtpBnvq96CEa5a1xocLQW8R3TeT+D4MwdFsZ/DSm/Tk7cEw/DMR1mG
iS4gGvJH1x3UwdruymLtTm9XjflAvx2XKLyZ5RCpug85MCyk0405vONKqfcduVD28f2CaR6NnN3b
B8kIUUMvhsZAazKS1joMuyzGWHz9aXX1pazpDA8Gb++vrn+SiJRyRrIH/Y4L3+3wUQBIWJGE1n4B
MAneXYkMdoztDy/FfFO4I74hzVqeymVQl5kacVqHpSo03PR1ge+P1ofSO2DM9dukxJurMT8xMkCr
OvoxoZog6XK9Iq5trIt0xF4xaTpeCVoeyuCEChS5h8gBLHpc1csgVuYSd4ApqUZaAMdf4bmiquEp
c3iz1aCgzpzcMBsrQXSqrkNUr263UutegS3h59rAdMf9OzvWDi40969I2NWFZmgHJA1Airk9X9rv
1iveiT/4ofQ3hY4XSUPiBXmtfaX1l7ztRMmOxaPmLKyROp3ai8C8nfu87v3iIAc5Xbvy22CLaJLd
EjvGxdT42SMCM6LIOlDadhnQbNpg4oZgVDPGvFy16sxnunNCpI0F4DpsR+ASVHkW1MpKiHnA+OFJ
DTDF/10n5KqEHT5vpVgtVV3It6P+P6lL2VXEViD/7eGnKBk5WiGGpijr4pJBQRtCPNtcwQv4mVXs
WM1b8GLG5/FgHaeD0gCxjLZDxb6j1Gtiv9HQW+5Owdow7/KpdLNLf2ndoTn+kedlqV0izn8Fdcng
kp2PvCLG6QEcFINV9Rd1rideaeZV8m+jwC6/d/U0C5O6VJJgAA6vNC4ohAwbPklSmp0dIc4S9xqT
coq3Hx7yl8lgit694utT8Z5vCZlkKIsO/JD0xVdz617CN3AWgndhXgX4zeiGMIG3NpnI+mRbBOrm
19CkcwDEx3afa1C/CdnmlK9S6n5xnNUsdkaTYfRxClpmFZzwbK17FQP0inVJU8ucB0I4IG7w/SUr
A1GI+VUjya9R2zUy5uhPzf327zcMbjMxrRzVRA6vT8yFAR+qdZl3CAHlLpvN7p1zE9ETpwj9vQEM
Lo43n74z+zD6aRo5hgsTDJyoBDD27mxrN9fbMMZoAr/crHMcXinnnvKEX1XI3a//kDRNobLf11Go
vammETXWIGtyTpp0qCEkNvrO8vGUywArOU1etRHiCnMEB+XXKJcEP5yi9yuoIYAjJxEW9y556HE9
q7eBrpDfUcVt7wSmEui7Js9N58LWR5uRK1YjSsxOJhqE+wKMN0vh7j4+gCoAV402JoeLtpYaC6Wl
FQV89IOOgbLezOlS0KePzMPj1e6gmY3uyvYZyCqiGYsBs/O41gTAHWF7a9g9iBZV7dTsQyZTjr/x
v4yLxZVW+itdtCDY6gKaXoh3v5PLSv/xE8v2VGVMRc9NePravzd93IoGWjY7pY1MyAeJ/1ZmUzHC
nJnJwrtgL0GFfwzfV9DjgkCK0oy1SW2m4goXiUIxb7IAQmjlJJ9IM4eHEnPUWp+XkmmNzV9JESVj
wbVFFJtef9xZECn2NRDthbWXd7CzFUf2T6M5O2vguhrhxusqkg+WJK0MDcYfcrxM8tKKRk3BOwbN
OSyfEClXQWhtAomzm8ARVJ7GMYR9cuRUwut4k5alpsf1X/gY3BDHEJUa7w6BZfAgXuQNweM7Adpx
rlWICy2oGZGPd5JuSIKPb/4xmaWoCOniEnh0DIt5cks2R3FVhdvGmcwgFuzuEDaoBgAAzuywuxbr
FAXRuciSaVFCwFhATkF7joLOLpWMZeTFqsJJz+OLoNFYWwhkeaNM+MtLYomgx81ytQYHSJLbKG8w
nxYNSl/xJ4ogs6sFkUnhl0YzByob34NGHDPlZdqYZgh24CsKxGlsLp76u6GPwxeN8Fr7W5JtYAG6
xneKrntnuqh7jOeefJsAPYTUdo8PZcJayKGJVr2pSZJV0YrLI2LlLwyQZcgIdjRSsCCxL6FETdd/
rfQg0ikCykpHlBiRPNyZq52beC6PVFfVJZUuUHDeRXwJ8B5QQDwAesC8gItOnXz0t1uJCMkCaIKN
V12ty57cX6qmlFAjxFQR0yIbD12sjg4nnFmu0NRqwESDYh6c6Orw0bzlkm6A7iIL8AKjhHJmLx+C
xcuT7iwHQQP/JFtg2w4fId7Du/UAA9di4aQnsjxFL0dslbGPqW00dnegGoi9hSAD5iP71JgHdv2L
Cr3LnmR3NK6QWGeY4Mi1MAXTnoizu7/6C+R8QGX0fZsjrLSNSeujAlxj3gbVRQ6QIcv3FvH7e1gF
jR+vlnWmWBCv/2L/LIob120ew1utm4nTrA2Qq4TfD88J78gciGBG6d5gNNvxuibScXjGL2/u5tt/
5NVs6CZAkfj7mp/of0ZKP6d0dSyOHsR1rndMsKYlDOSfMREW9ky4bWUmFz6xJFcXFtDdKO8+Ajvr
NF0MwiPNljdM/LPhnyNsDLZgi9oqCXNCRAzShMADdBj/hXKuEGXP/YkisLuhId/fK2dqf8Obx3KK
Xe6NenDjgKotY/+m3cZPjjio1+dJo0cly0ME3JaHz7JR0COlOGPDS66WRhlcm3Ssf9w6HJFrS/6T
N8OkFBLHglVboZCynYe3klQ2gHjJji1jAJ6R+nVwZCRT7p6vvbCJsF9GJHsoQEVtRe6PRzgA4GUh
PKL2C9Kg4Mt/H51V3Z6BMUWVHEygD79ir2yA75MygnEQYbi2UslWAC36d5O39pJPXwAguz34+NxL
mL5AH6MjZc2NynLsaPPK7r/ZYlOmNX9DP4edRXMFxgjxbW3IsdpnWWMhO99ml+K5GRa5c5Toa0E3
zvAHhw4rRvqjpV+Xz5w3eqVTAaoFt0u7YNlGcYxL+XHRgeeJH/4RYnz48NUdy2UdFV4S4sGLy9Pf
6LJugZH+g2dygCcLXJ9f8K3wwo0HUaFnk8RwY6QF8Fue+Aj+IhZWO5U/Xy/36lL1LTo7Kkn46Kru
y0cH2z1FSKs9Uxj9cIFMlfo8RvwR1u4Aw4d66jAKlQwPG7MKqPCkNeRAP0zOb3hf2WG6OhdB7u8P
Jx++0/uT2W24AamZl78pnuuPbmoExXdEgM5WgmoHgWvoEGysDDo6EpQvGuu28KRnskOjXMkpyPqJ
pFal1tveifJ4flyl450pm9GrSam03IT+qk4f2DHtRoy/UAVSeMQAaeeRw0yVaVPCsjUWVispdPlt
/5W8EQvH3394nJXZDZNDS2JXRgT7v+OPLg9wULZycWP/avGIee9HBq3G9fc7ByNbSAfDc0gDjCgb
lUupATgN6AbYfRJk+7nxRAAS3g23UBIvKgjGuTPZvckwJG1D74sVKIqCK6LkWn1hpUxvB+D7wF24
RaI5SQb23DB44LpCa0SEypTC9Nxwd6KlNx7LfVYA1NvwyNKx6tMD2/iAaNJ9u1HaaDzzkRodyc6o
cRrgXR6MzT5JNTFqw2D5dwVc/AWeL8TEfVuPfVJw/SLFj2jWP6iahMk6pb5eVumkW3zagsMNnd45
QDwjLkLOhMdh/vlzSGG+uuZpYQQ8b5nL4ZlRp7BZj+fvRkBOtZTlo6V+NU88xf4bl0W5XvDqgK/u
cwe5EpKVH1zs4VbvOAO4I1BqoUmVkGp3QD1TPJr4OjmMYPc2PkEzFPuuFmSvEvjsiJV8beaWgO9I
Dh2iDuBhjTO7PhZFgAi5hcaxE3bMuKlYz29jKP76grXfua13ahRHeS/kIpZz4U+n9i7NkqhwXiSN
MgYb2s6hGUY8c+VV+yP6sVYZil/w6Wwnrju7lAs55AXJVW1PDfZThi5cY/M+zUYsx2jJnStMe63q
z/LrpvuLaMXYF6lE8+C9yseZz2AdhX5S3Wxchd+cv30IEFgbI3ViJ++3siyvfna4ruwzT/zssZNQ
JTQpOD7qqTn46jyr25t2xEhhyIcxQhoCuhJcwoCOfUDmriaLJ6Vyr6U05o82W+Aptt3weVdO6Rgb
bm7vnWURhHDWgS4iwwal2gelp0DOOF3nlYcPszPKY4ihAzA8REEmOqxKeFJ9itmMu3xvHThEHzvN
VJY8dbegm41ElViVxsIgx2bZP07CSrD3OCDMCm7JpsWDWGHMH12fKTe2M0jgBLhZOVBBDT5BVUxc
pCsDA/7PNBNxv887Qz4nx5PeSuxPOk6yU9UPjxTV8ez4xM1ZSaoSYjtzzYsot9MMgJEO5kttZUlh
P1NDGJSYX/5te9MpnCQ7uz8pGTrMZ+IWPaEmAOh1FprPnhJwXfH7HXBOoBBmc70nnRQxtR6ADO4/
3Drm+rEy2j9X9Iwe1kfOP4P5WwIsz04SV1zM3YXRLq+q2ks/31Yz5RWsiNRDd1/bDoJ+vyJq1vQJ
yVCHfERX/ldytFeT6ufs3OOpn4UG/5SlG7Bomi3M4zYAL9awRoj+mrqBMYC1fyd0ngoDA7wDN8G9
7Yfa6KHet3Xt0IbwJNzAu77eVXa0FopAZDRAAKx0SDbUdgzwNP8X2CaUyIoxHqqPGmx8SluOrkig
pgA7qDawcAH70BonQEHhYv2tW1I81xZltLa1H/DWwko0oUyqTTqsJy4lirwdsDsFDxFwIwMkz9MW
miVwteRFsff77AWAgJfn6V9LsGHr0W4UWgvrf4vW8hJGyIBjnx9h+tZxyUaQZG4Fwetio0WaztLQ
vBRA9CmWHiSV5x34tSI7t6Mt96d77lznp6jUgEsGkZmHdvYw/a5HG/LxcuRxfGU7L3SQWd9Jhzj+
zYFFQPij4/AkMSB8wBLG+UBriVMZVxk/wdpy6KJ82ekymgWQnj4R8l/Zt1xElRWJyv5N1IdB6QBe
5PQuMmbIra+45apJjYMZ3sperwWiZp1pUf3+L6cqeoSmNeelnCu8FnRlzHpZ3fUS+RfrmGiocp5+
e+5ilAYswZA8dHBokNc96NxId0aQseNCF53ofAxSBWPhAR83II5RMC5qeaT0kgoe8NGXej74tE/D
e7ZqrkWkkDofy6A9O2q+PBINjwKox3Ahbjsa/Uj1qZxLr6OHNwqzm8FxIa/9+LZarrL1ApNpPI4i
2d4GALdzN4cCsophFSRVrvn4789PYE3VdfQwu9q2SqP4+dVDm1g9pTHqvtuh18oKnCOxyiYt+syd
wJ0QywwDDsiYnjQU6n0ePKnSrMElvv7QmX6cT0v9DPphD4zCs2OEeqU/mEXhr4bfqA48/JnlVZtC
AusgfTFIbHJEbmwsQTJehERtbLcAd+gSwTvhLxTQARPUVFq2twe2mc9HC/gWEBpWacUdeTCZQXVz
W5KdXJqh5V8QZT7P26JeU1vcP4AKyLfPBOXe/EP9yL64ysgfRarSlT3t6aQLhOrjodtyd2euhnQh
4dXtpT8Iv3fuVb/0DMkWULX+ns4+t9+OdCNjsimCFf5flzExQH2nZ+JKzE/RxPZ3D+zg6YwWwpvh
eEHc+BIg409JQaHwAn6/VRTFNZtFzt3lKWZzb006hVB2mMjieTUweM1h4K/X/qelUaWf2piIxP2E
I9de9EzkQLNLmcaunBZljCgqwLuktk+K6lB7oTszh6dCzKVpFiFBqGD3F9v0+HnY2HuriHVZrius
/Y03Q66bTsOCQaAxKiIrnnYpraBItbSGrcOKD45ZwSy1Sy2ovUvJvSpGizXhbAy49JL6hiarJjp5
GjG9T5z+sWINBN7zHbehA0b+pRG6aP7Jo+pS9ZM/YmyZtRzXF8vdCXNPEGwwzBRihPjfU8CIVa4V
S9A+cqoPyHDNtfoHtPNN1t89Y0lVNeMglvm2wUTgAY8Da9nldQjkXipq+5ovWGc5aP/SzWIy4mip
/8NH1ENaqnFB6zxGssT+XCvR+SLJq3hf247OXnZ2aqdmXtrxHsg7eY/y2t4Zlsmigt9TlX/ui4Je
1LsjPNyPQvmfULTgIsNliiq8zp8CDBnPzsB08V+1QTDVgF+FW2Hypmj8aTEoKNyfeScqQsWsZstK
ALAzOpEJ6cl4CRL5w2zwG84CFkvDN5JXQ6Dup0Kacw0Y4MTyw9STtB6E+OfN5nvwN2JYS9EnqJI2
z/0H41HMU2M3+ygEIQnU+Be3wK40zUE+2mE1l/D4IHtW4X4WCeQoB0AAqJFp9EB0BWZoR3Sn7CYs
1fIDbWZ7ysKmdrOw2WA6fRrxN0QrdYjwAnFf/035CPXBmigGEfjfKIylKg17YQ9vJj8N+nPrgbDy
XPmPTGRqnlltqiq8DibN7wDaOD3u2sOuAL9rda26F8FtSe5B6Y2czX669G7ekSXW7rGdV+qZdSjl
nXXbP9hmj3Xtkn57UmbpqPT37Bi+TwxnGyDYLyWOScFR7vdDMsQxJq8QXPpVl6Iaz54ZTmA+Hzu7
rcB4P4/76GFUEeMV8nQ9AxVSXv+LghAgLQZ2MkVa0DpmNfJYTeIQOOTbDT0jDDDj5uqmIcQKF+j2
wSg5W7KlXFx5wPqMmK5qJdDzwJwXA7fzf7MvOCjdMg0UXWyY0uUZbE/LwsU3jNev2VQi/+aFIfIw
3fpJ/GEJyBaYpgQjAjH4I0w0aqMpVrgOe3xO1d993nBnyUbybmhDf0mRkNI/RKsHtSEz/jwhla+H
cVuY2NN6SYxkuHr0wMtFa8QTrw6wXcco3mg3dj0qRzNnMptGi3871s+J8D9swrmo0YwjNvy9zRne
69MMWX+KMZlDSfK7PZNKlmdTnG+P4tbJxbbmC0l3ip/FYT46JIl+enFKpKsXdFBcxKWVo86pXSzx
KjOPSSOSyy5XG9O9TwB6ltecIDB6N4QJFtEr58fArFYZg7mdDiK/ZjB0hX7CJ4JFc8VkE8uzyQZE
qNuFPayZZ4ubya+q7+G5P8fjNqMjtPPwa3GrolANd/vaSWLiNjipxYbXfUB2ZWoRZBbBoJXURQ6W
BQMoxJlhJnQEHfaiN2f5iyMaYaLCQSxDXDt0i/PzLmX7WI8/3Urq52WqCp+jwpsJb9ZPiI8EGT8p
aTpMPdpJqFb8kqaavJN0ywFJwOpeJZtKpEVo/L9MP1+QwJVIozdw5EdmR0Gsux4/HosiT4Eh3iKC
OuHXsei6zwKYXBkmmhrFXsf5e9jWQypjoI77dIOxtbdsguhB2zU11dw/RePZRjtjeB8B4GAkJbAQ
BuGjST0wUDnnnb+t0lDhqW+EKzw6rgfwzqlCeBUNX2Z7gOwxe6CFie2pox/6EjXc15TXsjcuD54O
BKXWxEWOPrKOAJ2zCSnqMnYsvhiJwtL9uYliIQzuwiIAG05bWKdSDTohm2EWp3hI43jUfPGAVdr/
zAuxXrX10wnMTwonLbF5uPpPScdJ7JWWLeEMSxh3uJiUxfXMmoQuYm6ZhIJ0qvIE4BSYyEM41XHZ
lP1mLdhlHJlg/oHvfGRltogEDz8ftJJbDt4Hj8NGsu3MsFvUwxp1TiBGmsBjHiTtMaxww1qB+Nm+
pP1TNas7jSz51UR5ndDo2WckcThQ8nrluNNaGQ/36UhJBxityWN/Jxdv9CyaeUIEAyv5XDcKXHn3
c1k/+3dZD8jTnfnAEW16PcDTDY0qZzXiEAUEmVJsXvo8pgNikpLsh9GfpXyzp9Uc/502IcglgyT3
lSBVaE+uqYpaujhjAWlf/JcRIE2oGtJZjFN36krpQn5qWpuDPa1XupBguezNqCgtEtEokxnNIgAc
WDHBdsJlFsC1D7qWt1KXJFK1ILUObHrCyx8a56Qzn6yKUxktcGVQ6UhvArafuxtiPZA1I/N5ilWu
SVPIw5qXaCYOXEvFH0IOGQhzTzC/jslwQSTolQ+Cu4PTICOvXrCQOtkaw7NeVlkKnV+naRGFoJ13
qf3XoBUdk+D7FBDiXlX4kfmbhxhhEBSMi/I2AguIeA8X6/UHi/bq4mQTYCLUHRO2SgjKRqJ6VL4v
a96vs3A69zpB4zKcRCa+v5W3zoYzeJYZh3lCIW7JSa51useSQ3TNuWzvRmO3YJQ0yZlBQRY0VhER
q3j4fxL8pqGr8FxyLgnwbGwi+Z73XoLABGBc5qo4+6VQtzdfMn0zOe1sgEcg3W1f3bFVX03lwimZ
CAAX5SWNEa4FlmdbyqhxHxY6JJlbRAvH0zZsc2KeG7jF0OfXNaIU/bpP35syvyGGKBjIDR8iyQe2
Nvqa42Mgy6WdoiQI1GjBU4rWMrVeleC8UOAdw06Ju9tINcQJoWPEbU4nFbcYsL4983YQDacsM1Hh
r+4M3o1WrgyIfjk3RHWhjGJt+iuGwHo84HWp6vf+VWmr3GAvBoXCv4Syg42Hqbu5Xy2UXZas9Ln8
V9pLp9av1GnkQBmM2E6BWoFL1Ry8SLWpz70uAedfPXkkWXPJe2Kn+wSMuUImLnYCijCtgT3gfInz
cc2Ss5mysan86t7lpmR3+uGiryUQLCWaTLBdL95vjsbOM8xqivol8o80eglSlYHu7fbzOh5bLU0i
Zn0hCdCTA/gc/9yMt2LBZjUM+ThDxv0Ul1lV75Kzh8u11NOgWtWgU0/ddB+ZGMAyYLFKwlYSTqfr
is/T1zxZpWxW9oZtU03yTfLk9yr2e5vaxHr+JDibgCLylEcxG7sds/ZEi1bNlP/2Ih3F1hCKTWSm
FMy2yDeK5qKyqHqmmeZQ2dDSGcnudv19IfM7/fZsAOKEiSkJhbDZjdgRoGwDhzjS8CO02vSt3A5T
p0UaCRp5AmbvlM65S+GQ2KLCj1ce1w3qyHfYq6U5tDoiAdAMCnvNTaVix59vuPKNQ7p+Xgtpd5gZ
8f1hUvg42ibOFB9fnmpLBuItqPKpoddKOwTdBEap9dLAVnlAgglbZ+d15J23IF5f0TieC02LrPm6
ovNNX9M1BkCij3pQFgMGy+f3Cj3XYRH/1jjV3UN4O4wZ5PzycfJ7EcIiJvyX8zB0q0O9Cw2+E2wF
ETOWYo8fL9tSIgEg8HqAsIBEVVEGhg1bUQWHMY3d2DYn6czJ6oSm/CrFLOl9eHIhI7j8VI3zN+ZG
AHEQOooxHVz8coeXU78x2+LiS6kHagWoAqFzBqp4MH1YNER518mbTzJ1wiD8EpUd0IeINtvZlvsS
XOoihX5dPlQ2byZYq01P6c/QYu+pym2Xvgd4Wt99ylGwB9P+u124ji4LQZoUk9Enitg5WB61L/5t
P9EI4UOSRO4v/8NWqmXOzWMVf6vYl3V5/zGnAmeOsqfe73MGipNgvParRB5kLRlz4HCGUgLXUPMZ
euCNIHrKNmX8woxzNMjwNY/MNqsuz5kDaH+UxQfT3Yu34sKDZZuk1V9uLAUBnw/w7erqjloejJI0
ZkN9ZVqGsM9wR1q1KdLZThFdXnTubhsmiP7QA04FzjRqOrIkAocfsXFrH0D9we8fCF2emd9c+veH
FN4YPdqZ0eD0kKfpzLcCZBv9oVmbIX4LB5S+hJUT54U1TUdjYQ6F0osvdJPO4luiqnVImoZqlGRv
6Y0jKFyzkCqBxM5ZfIOVd94FqqeudQ/iUGZ0jUJ5qUWvHM98982AtbYews7kTD68B7KCvFJhXZnv
MyOQVAGQHPz8RcNAytyJCueXuA1sv2Xh5xSZB9P2m2iJp2ruunZISJqUbhY/VWfVdCc3YkNkSAHk
ll2avYPZ9iVhieYzyipxzYokodPAPjWwCb8qEK+J6T9dVt3jC9b85j9nHCADT4Nl0M3AoIJQap7v
HWMCXez/6lfbllpDOZQChTdznJjQWRjNPmMyaZGwWqf1Oo0kzxqg9iZfiWZRyt7KzQmUxsghdchP
RRz6QTGXDRrAnjPBmigMPdmY4izqyBWqF0GPYfDC/plvnyHDCPgrDFnyhee+HcpT/feRkPKWpSgq
pQCaoWvHvdUv1Ssj0Ojcs4FiwM6zCiNeEI5AA4Pdygihvn90J5v0yCFkts9EsI7zCK62zvqLhUs3
QkXfmR4isH8HCVnnmFR80FPkUSkpwMEv9NfkOBgv8XLpTuHNGyWbjQg4n4s/0LMcLleBbobGsPNq
RCw8F+fVaD8zq+U/mPnJckMT/t/TyIc0/UqM36s9QDwvOxS+lmwDVKlO0J6aQxSy9BIDcESb0oU/
2ClOcT9OJryi9NZ1RcQfJol9mL6eBm8UqCjRdCPvcj04+Rbym/u/311lAZYeLUHP5l7r69mnDuFQ
6Tph696jdiYkRBwH3gVX+yMiIErUW4366o5W/qR8hFbao/9gE76TEMyB80CseMcBdjDVsYuXm1Ws
p9NnaAFE+Dx839VwLYL1IkDhTyYAiLf0ChXr2Tsem6VrmvmRJedc19g4nND+bLugZKLZMA+7mrHc
F2ARk2sCHKcbvZTuRgKpa+uezk2uvRDaPtRTfh1cMyk0nrWX7caYqP4UHxyFvwkDjxbPp9FIMhTZ
GkJNX1vqe8jKHneAK7NHX7Oh/yrQE98FpBT+RWIdCxSKLcfILVZ1nIXgs7g3aEVLGEWAswutwCJK
au/YmxLJ4j1ZDqfCeSR9VFS3ZELRhSIR02qxMp0CN+qGP1hCDO5Q4GMBrwMKA4hU4j/sse21BtdD
3qoWjlQgUO6xfCLHADAV3S8TMHjeu7P1iJO7IThtFzvjEL0lEWkHxOgOEYpV6buEvTohgGYuH0pQ
/Ml9ryr9cm48o4T99RRJbPaU1bJwJtIZBnN0fyLDHvEuGB1cyDiB41oR2bf9BijKsaKAbcLhziL2
Chgk3fGLQkX9CYISeA1225JnZ0Jv3TShZ91SQdIWXPvz3th42HrfRcWyV60khgdusGzi9q+sVjuc
yKHPCm+ldxDhfJJySpoC0B2E/xp4/ixrJcK2dtByWKWueVi8B428cpVeBN4kfhBpz/dchrFoGnD/
yyY3vr/OhzrBUGt+TpXsAXxP2eXAwOLjgURtT3HXM1RQFEvQSMU3Gl0k+tnjgWO00eJ3LHTOAEw6
c0yMu/Co1lLw/kBzm+wiS8VViYBoU/Nd+fbRjkNmnM7Av+Sk6ZW/tsmvokcediyFBiaf1QjDKKSh
fIsvnBlW9XaXVIumKbkGTUFev9tMJ7TtjmcJRxKjWcu17iOt7QoZNGXBATNBAJkK+H5GGl/lMauc
L0Otywt104DrTL1hhAuPbZKmj/mejQYsHVYeL7Yed4TZRMHroi6l23cTnFzSoWMrsTg/XiqHYDNX
tJ1F77oTG43FFuaP4+D7nVzWQw+IBCGsnz7NS9dsQxhKpf0hTncl+XfPjFfePiQ+bBvI8QetXTs3
5NFyNoQ2V1lKbr6WaQxmbqSRad5UMYxTPuNsuc2lk2k3TvBguCAscbGq/sG16L1ThoK3ajHLJiky
8lcZm0sZOcMgdAxfmY4CJv5DtwPpJmE9GZSy699md3Wq9VIx4oBGRGbnAM0HfAs7dCnkYtc2YDZY
t6R+71JVSDEP1DPsxvb1iCqsPcBAp399xQH15PZbpirkN5h+jLA2iNCZ/3WUl28hBWTRXKOzgRrp
29afUe1WBmkhA5xvTnVkNuT5ArhwQYDjhUj9+AbgiUpzuTh2bJ3zdnHOeLOqGNqKI6Eq134SimEn
yJo5y3OEdw3Gl91ywbvMGakXuCp2kI+6TU/PkjlCR8wUKG7WjoGCgGzyllrBizU5dD1jAVqVD7Xq
Qfavgyn49VB99vBLzts35tjg2vNHs4HzqWC6kzeQy1wqp9H+TLEXzSCmyfqFHhnMedMIb9i1fPL9
qoGo7vkBHvtXFubEiNpIpIhsap4DHW06jbqjsbLDH7HvrSp5aRxRozeWOZFMzuCC71FST/IcbiKd
/YSeINtms7XFu21cW+Adll6L8lgv94Qe2v+dnl3+nGkF1+d0cKnVOMO7X3VyDGr+3sW7g6Whcx+C
Kp2ejntUqJAhbedd2jRkelEFvg2ZmRn7NJ55e3/4EERnTCzfcJQe9BTERPJOSjCL7c6/7qVJDE9R
BvF9Um/7Jgk9Fr5jKtuJdrf4uq8XU+RhLDl7FpbqcbQ1O5MyXvGnF4nXM4/L2La+nt9BJlaGaf1H
5RAQJJDURFFk9sihRp+ydqJg+THzrVnF9fzsQHyYjSFgT1gYNfJ8yZv9r+eWILPDFqDCYCGjZ9uT
lhA6k+7YnTLmt2yX6jgjTrupRwRhaKpTcUc56AY9jp8Vf1CmOzwOx/vTfvlvwB6dxVhhXNUP95ka
7mDiBJY6VKVl9/0hCAJd8LTddTnA7gwDGNtqJIKYv4Eq9yPemaaU4abApWeyKJCozi6mSJEvJ7BQ
ulIjORHGydMRCrGRMywwraSiiTvP4mNqwTkN4at0Iprq0l2WUg9FQy16KknwmUdhzJfKVJxMi/vg
OzDoo0PKu0ggZCwEVjpWTc5FpV0Z9Rx5mrTQeYXxUm1PmZwN7wwSZ8qsTK9D4rIHTbzIq490/2HP
lBkN1lRk8fAp5zFXZ8yFdhTr698n2sHGSj/2uBMTaPyDgiXEdiAhhmvRGoZdaCc5zLeXALQxRjWH
2t9mnfzJPv+zT2x3yfkA8cSpgTJA3ueZGdsg3WkCMjheybed2SrG3OpqJYPHHaR47fFxhas01rQ1
sjbS/5pPi10PKP3kEhGpXw675PqRcUwC2mSmqD4GeSA23Mc6cOUTSdIHGdDWgEFx7ojYFdG5IZ20
eCIOlVm3v2fVgIdDJbWsJ9Okj9qCs+IShJmDFF7kQBk5ddoSk8XGm6YwtetYJLNXDgZTtqIKanNX
ooliZp75tNzs+JjFYtQgWV8/AvFMOkJoN0n8+RAnRvm8kRkASIofWTIrEK0ayaP2soJlvXQO06uO
rfnG405+oZj7lwSjffD7oQiyLsc+couwjRz+M6kMvTnpVnlVePazjgS6KX2PmQc6QxLGEL67UVbD
9cEEt02a+Ub3/WsivP1mMAq3WmTmvLa+MsF22ZtDYJuTzdSo8E2X96hXlH2nf4AaQoV9OiDpHsD3
o0XYw5nx5rhq8aqCwwkDwQvf2aEHPuTeQcfqH0GsaQGBJ9cM8Gn1Ke7Wal03DiTPhDIVaQHsK3nP
a/yIYQ/+Xk36bdVxA3vWfLSQT0ily9SMxf8g5YmcF0fzxxQugAbXd0jHw7j64TwAoISN4N4evFzT
jJ5A/xizQimAzPdVMHo2KdH6wEgQbExxxVDNM5gtyt+rV+vz8gghfhCYoYV5icveFJ1AtvzZydET
rjgXwLA3wvLu+p0kXOJ/1nre2dDCFhtdDUEvXlI/mj9x1ZDuVEChJGFfEb8Ab2ZKNSB2aJhaw192
kwuwnJMZL6umzckFdyJDXSNuqeFY2OGCKJGFmq44sojogY6LwPgxnrqfAlyHuuSVk9g1JM42WijS
7DUeGIs2bkjeDZi6G8tAsCoZVMe6fc4MdtOA7f/J9OW3m1NZwAnTzykbZcQhsm1w6y90A9dkz3Mf
9JU6WG/cZWfVN3jxPZ9EzK4M4ByFcqK6gKDlLsfEaIkd+pjeIrvKtdjKCdqETj5SGFx7RI96fXce
kV7+wVsM7eU2QniHInOqLCy6Bxokdod6OB4QTXVDdkJCQ1zNuaEALdfKohzacEJnYyBZskkSAfDn
nVtoOzpz3c88Nqm2Er4Ia42X9d2/6WzfUp9HvLmBbLc66T4rXU+oqCZbNVIMzHTVdS4gsMKhyOix
3i7pFepJuKGzBOpJzO0n9zP4TRcmVXn0+NsZisi6091ylgdKIgrCUjzOWuAoCY9Jc0Hova8f41+/
BcSMbBa+tLqNrZW2GFN6b9vmA4/QQHgKtVMxOiBpTs1TW0vaB4wKznkglhqR84F/6KEDycI7Mrkz
yPWAL+xfvI5jd37+/NpyWL27RAZxts6X1duqOZGu3GEepmL4wFu1U83lv2oqR8USImVfdIt9rgYm
QZqnayyFXXe0P2lSi24d3iK/uMVn/65shNbJPHuELKno5ZHdM3ZZSRU5x/l3TSursfxqUMSBBVNI
ZMLCQzh4fklt64+JdPaSkvl5nF4zDnf963WKJaBMZGdxOkBouUN40rM5Nbg9gyWtEO+79XF/3mbX
8CdbVOQTj6UX41jtjCgsj54c7PFbdbia/lke1HyVGqgVFwoGMdRcjSgbIIDBbhoR6JXcH/wmYuZR
ZtfHMsWA6MFuDEosEBAm7AeKIRKWl+irtqb3hYm68GIax01Rsn+lPAbd+LUSK09tjWpDFmLueFMD
jlZBndk1BEXmZ7WT6X0c8fxvVHtgAbaH+ZZE3idgVMihwiyM1oJ77gFM6HEn5RE1UIH0X5kKZR9n
BZHXIoFZ1jiNf5mHWa9Po7TN1Ij4Wflgmugud+iUClurTTNDtxirVi6eCGOeVZdhIbOvgAtDRuri
lE+0tpecWwRbY7LKujp85979sI7esN/HyQMv1gx60NIJ8y3N8VXlOGFuO7kd6UHu+rTx5SHL4HVf
qcWkC7JX/ZxxoeN+whXHi6C2x6jX5QmTA4Qur5zgDGzYk2cu2aVlYXIMTeyFDb611yYOm+snbubh
98P0kx4nh9YI8YQIi5qSfthLzwPttpzGRq/KpoRuP7zylHc/eZzf8m3WEiJ4zF4kNblDT4h7eo6v
wRUezvTL3PNDHn4Bz3LJf2jjtQbI1NC5JcxwnTYOWf9HWlBxbGUdw33Prc9fds4I8J80dZIe1q6H
sH1BaKEb8bDa/F3XI46DX1ynmEwS2aAl98w6Sx/OaWTXqRzITw3fs/qzTuf/Gw+fubVjhXZ2mk5p
8ARsbfKV3jd87t1sxvaE8D9L8LfjYToomSdB/kp73PVOZz0Xi84AUOePpexxKzpml9FOTIjrTdMp
Qdq15kAKU3Dab8CrHSwUUFiYrl1Pu/oefFG5KHR8VWkJse11b9qeoEo4RXcl1jFwR4ttbWYIVuGG
q/qmoiZtfgr/UZdDLw6XqAJKX/+XljAAqKd8QQ6K6lmlyBioMQio6qDXYNCeI3x7eejbfrLpM05I
kfK3hzSHvOeMq3EQ6LdwTZL5Hz1eBI/l6m5GtZM8gUaQ+MKtFHIipVzOur5R2CPdk4QmS+VxNwsj
KCTEKjgKLWUskM6vPspM+h/639hZdfo9e/rgt2BsnAPlMP1QrHb0U1HqOcA3AkzEEZjex3ICkwOL
hHCBKsSgWmIMi9AQYp8cfQM3eBLRt4+oxTEmGKFHC4DOIUx6cIyOcWRjx/eAFNxIw49FF8LITv4d
ayCT4OWbPXtygbcUrG0yoXMKzRAlJd71l7Glr4ns9F9VDWEYi7tQOwmCBxUj/7Vj8L+/pOd5hQX2
ON3/bQEYZOpzJDt+PdsD70AQmiiLEG1P/b5U656Il4PnOJleDN/LWsrPLRccYjt5UveaR93l9jIT
dSMfq5yZf3QS2ww7EO+Bhcd/wTGTsMu9m9gvLVykIVmUuqabukuFlrglrLvYm5OxinBbXgaQgqPD
NhH/hDdv0uywAqWo1a2ZjPFlXoU3ezr7dZvFEWY54hNwQ7Z0yyaNJGfp51ZiKrQlVoaxc/cFnnL6
xNb3/G6IAOzf5VOQ5gBx3oZW1nf9upTDpVeUjKOUWV20fOHisNr6SqoTkcP1SYkPjzROwKTle0jp
ie0JJNBxkoEek1LcL/CcdhqD7dopAsx0KZdtwpeaH5udFBCPIaPCnp4ob2jGrEdVpadRPy7je9DZ
9gDVW1k0izaETjdmL/k7iAzIiT1Vd1fuq/oOHnykIQ0uBBEfD5+K6r60ElW8wFf8fxyfKaDzucou
eY8uevevVvF1MgsPY0RW0YIAeg1XvsV75H54+8395tyJ54xNLubdmiOWBiBuMSy4oYZHqW4cLu5x
OrZtzp2tHQsqr9dYEX9TexoWGU42G1sB7PanKkiSDDnQq0C06o5ywDN8jEgMAQbgmytqsBr7jFvM
F5T0ToWGTfASbJZF4LhWdR34gD5MxBJAqE30olE5rdAN0wA9qSTUUbTbh0k6TT3dYRJ7hXU9UeUC
1jNCxxWELGUZdAavco6+XUHN4+scD87OYVB+iQBCG2k5XHlznnpZRVqca88mPairgDlZAiSZ2NAM
RAozowR+aZelSfvMCApq5ltvd1Lro6YkCOlLQ9jwZmJF8cqmnmFZlyqSpOQgvUQoVLglcV6PqAK4
WoOIOEnEST8AI2XbfghAdRggCXeq3LuzwqrLOjFnhTteirAJzDEu3KUWdKs4Vf/Mhdj3Sg8KSx6q
q/qzfo3QR9yPHV4yqDvK9DicBRhZTaXiFy9vqKT/lf/mtCrhgwgwutpmazCCYMzfPu5l5eTka0Fe
r3BCVZXTmZLfMm99JeIDva8jd/a2lE0LkSQ4hYMQdh9MhdRDQI2fNLzc18zXVX4p22/pQoo6WDhc
xTOGRGCF5utRhXJagZqDnjagC6Q1NIW3TUKRS525C2zorGzPlOhSyC5gCMklUtU2N2Dz4747VnFR
rJCT1ospVSe3bOgEkOAJSY9srVC/YewSQbF4YFAbh79d5U5vPxrpnE1X3zERKlhp1SxhJa0Hhpmi
iIGjEfUYhXxCYrjk7RMLhG0Sbz3K3uCUQorlwAYUnUMvCJ6Vp2AawLDwBeXIkv4mOi1lD6Iqn2n7
pkNrzHLNIiNytNqYRM5faUGp+ecCvKw4ULkniZWuYXGeDQA2R8gccxJVVoeuqdJyVhnqWTHscuKy
HcGyBRSEYaGXVhjyO+4JeQJJLIbRLJ6ESVy53+eD1bcDe4q1csqcr22bJMepnm96YhGnMeTcdz7D
z3ETpD1OiOY22udABFUbqDvbrWt/CUP9ibmsChUo/dFPC+vUQT0b+ZE/La2yvs0pXdehw8JFDmPi
PeW69ggftjVLl2lNkRTH2Xs8DT362GbX5HDUycXQ7OX4/RRWtNFtwrq52Ea4X5HCXQSNpGEL0N3b
UYpPPkcP8KyDq8f94aOp2G8AbxVHuuaEEwo8+IdxQj1wf3037xdaJs3wAA6er/L3xG5muNiIV0/c
M9HZwiHkoruE0FAxDPvqB852cPd6N8KXO3eOgLheZej2BEyZVhqz8+J9P+lgU4e/thWteuEebhmU
UZZBTg9HtLjFcDQ6lCn0anJTB4Yif63SHXPYclyu2vOZMXkjghiz7wMOFRVOLjBfgFkkqDvaItzH
cPk8OdDJ4KoXyrcVc0nNV7U51XPhmS2cx31tRyS0ErwAlGTOiLGzd25HZnQCLsQm+xmokSllSyyy
PpJTT37rJtuyI3J4UpR2OW+74NmhZ/c5Jg0omev4M6cx77Fs3vSczpZEBcRr4IX7YNnDOIEmDNoR
GaU0O+IfrJkJj9OBJ2lgXdIf1+ZIRhiWmN1upTMnk8dWkK6uiRuWIc799gy1ep6NZXGspAafed6Z
p7PHUTNNHZbyyXyEtZHubw8KvZmRiE+QsvcptGqqM+Sm3bArJfJY7Hq4Pqpu5m5GlLpNz3C2AIKT
gtyY0YbHgvjGzqDKX8HkPxT2WXTaMy2jE3gNrtOn4fKQKb5FlapVNBpdO1CP6E9DEzYrRjpgvS6T
A/a4Sf439uXQDpVQ2efyu6YJCO+gDJo8Ssbc++Ahmufz0A9Tn9qhH99/qQiXk+Y2P/yhEc5BbuZ4
/P3A8bYi8OfHoyVG8I17CDZ6ZDNKcTYLJtnKOtVNi8HdK1H7xSZjlVk0fr7EBDAByQUUE1boIz/t
AxflAe8W9gaZ2IeqKVhXt0qDyMuTGv3Dm7Xz5bqKYNIXjspwRIdo0EmyrpTd4lx4UUhDm1Ofz0/O
j/ZOD5rBhnRg0Ga0egiRurvMorWr55G7znCYnzyMj9/jtZHM/B/zlHttiP5IxX+zpbYb5eICpNY8
33mKdgLYMpLo6icOXi+0239Ob38Bjv6hfPoUxyH79vjPHsSlCAlbmOZOPWEhhfk6ehUhk8a5oqu0
i1GaAPjW5iJhXgZXmMHZGI0F/wor8KuVXHBknZm/Xu9wf0FDl1022ayieaTEkZ6UvL/5yw/JMo2r
V5+faNzSIodAMDMg5YLQSnYl+JpIo7M75OYi8xkMc7KzW5Md2hqokshDSNpY84z/EBtZXZmZwvH3
JBAIwlo303TusJxOhW27xCHZF1PryD1DqYKpgXZN7zOKBP40EHhPoDOZ/MquxHg8cHZIK0yeC81u
eOOW48g4dKBUQceaSD9SYy0OzqAHcXyK7Zx1Awfr2w0NGxFjEnkf9NRmkn+wiWp98/zD6RnSXXUg
z1JvcoCNLWHwSc+kAF/ocf7kjPaaUQShzPccBoB1Ed11cyTKTascUoKgttJ+P2y/BB8xgolAX5/g
8oiJ6NUUKZ8b//ZxDyBK4M7GPB3PVdFU28olWUdp7jUXo+rD4ziLFzTnbI7eGPZI7Q/zCxKufaoK
8m3tJ+9qwD9Lj6GWt3eTF0SlANEI52x4AiAjWrBzOn2IazcmRBa9Qz6BoJg8vYIXhj/MPJG6jzkm
SN4JuVgMZuLJIi8gvYCO4DTBXymc3I6LvZ9bwoP/z0mLGqRqHY/wnynpr9nk6De4NYtij/bztKQb
NK7xByTp3Icp9ixZw1Ho7X+HgJY2CA6pFgiMN6hZ8yL/fRS6QHZ+qZMPc7Ye4r/Y1IuN1j/uOVjR
yIx/6AuzDbUO//TG7GJysR6X6kc6UwTaX6B7vKzyLO0FXXMNH606KmOh8tsVKGwEKB9OPfFFl0OD
JgTdefigMh8OkGsOv+FQWD8VnbaNLudOf2E6wFADutkVRknBQzNDr3H/C3CXujHSp74D98MOgWC9
qn1I9H21JLfLMXGg6QHR2etuC3WaAtF01zszN9SaR7gHlbaF2owBkqKfh424KWwGBCVE5irBtiXB
1behfOUfU8eHRLtandRyeNkgd/6Wc9dygFlrKQi7kAwjNyeZNdgraBNZ+oddrlA2wS0zHV1yJ5Hd
LimeOoy5MsTDFMbprHYguzVjJHYWgQH6TFeukLWH5FQFtGiSZCMfZg7KsIYy5quMJi4dixyxbs3a
1RhdURMpXOJhxK7sn6BNeTH9vaR2rKcPJuVKNECSK1RDu4X4xZv9jzuXcHNg6T2w+gk14UnTIk3N
XaEHNml1E0N3oNAgIN+ySq+vW4QOgUwe+Gm++GqFY/3s+eMo/K94SRv881QS2kzCauHA+tIAOZsS
hODbz/nOKslkVHpWEFsGwugkA8FrZTYnzY7ibyJFOwAJSEJPrsfnXxKNsunPiJ22XUSFGnbXx+6Z
4g6k3l1UtAltdNCOgxzwjDKKBqcv74L0Fd4Nqm6px54YGdd4mVQ4vS9Vv5poFCc06uiv2p79mFdg
KdEz1D6SKBjPmAbaFP2est23oqNPDcx2qfeuIau+jD5HIjLOFidWrOhXC+5P0JEx3p7whB9Kl0ZI
hhHK4EmxHLh1roQGQ61pnUcbu2R/DFyN8GCsVFZ/72al31m7dLJFCGf2BWbJjkUOkHEYqhbyVGJK
+qs6TEw75GqZpAK2/AwBLTBtYwp057E9XDLy8H+efwzsEkuhZiOF5AFq2kXVRpIgvUqqHhdoAPvj
h+JzavWGzwEdLsEavK6DjXs26bGIanzasTwJxZ6IQTbCsUP65KVXaot6oommMRJSL/hXRGm29p62
+OFK9CkJ2L/z4obu7qlYjCRjwG4r6PLxiR1GX13Jiw1KprofKGElVQRyU7+y70LyP4iIztpXwme4
uUyztKZ5yhhc1Ol26RWXeKA0/b971GZZKbnCG5+4bomzEThr3IqYsgM2/lbEfFOK46Y88AgVm4AW
J8OKkh3aXf5TJdn1t0MpSAZXLkbzFrN9hVBuPws7YchuU4c+utwN5LTrgv/UqPtJ1D1dzF3Cjhbm
4qJTXRhR3PJskuInqsUhzudVQwdS6RdgMMEyWImiEVpQoDkcAkwNiWfO+AIOeG/WO5uzN/1sWea3
9FGUnpIaI/2VJtjyEM9xJ/xV7+yVjCH2oqk8JycCgJBP4p/blj1Le/Ol8Aap6KcipPwEYzIv/RS6
+/g8rZOWrvec/uffY8IDlgPwSXqvbtOLePcwE3nykd2lullCTWZdEqZMoh7q+tod7VcFmqP9ezOy
ESKgskGXu73SC8HNEuyCT8/YhXKQ2F+z3BDFfadMZUlW0xOODfW+xcqStuJHVZ0mZT/3d4t2kgqt
xJm4NGNYGkcSY4b/AVOFc1wDqe10UhUFhIkWXKIAYTJ83XCQjvlVSzDHLjreuokgm/C/IC72YNRR
QEboxFG3KkcXABjdUxZzwax6+7fCyesR2rTPLWcGSSk/tkXuVMj2A0uj3oVqXwb+S1A4SyL2FrAM
PFbDnlVw2BCkAUU/pq2ifvlIywZzIEUpBEz+9hzoL55IK3EqBLZnQdookxIdumQpk3ThKWxyoGsR
AyrQBu3JOuQdEFjc9BXr3IokN271p78XeDgegWvusCpmlUIYmNb6Y53/jwktqLqnQ4L+IBz9GHSc
zFvwSBofElj+379NnY7jySsMNuUIx7GCCSiQEBpCaYo0W5RdKgobaxoVUxCRcTelC9Mxd1DPs6cv
6+B2LnFkIHM0nGCXKXY3rh7iLrVpVVpwcH7VNDKKOzR1ZcFcllFViNcfAnDfrlG/B0w2pUBG77JY
vvWNdIBGdwdpLD6Gagg1E998AZOtbmD6a9aKD82xoimHczGDvHF0Nnfh6VW2OWgb+/4xPmyWlZwq
9yIdwtfQKOp66StHDJ6uUGqTL7uFLWLrOy8e5pa9NxxsbG2A7FChJYLFbRUitOlBgoclNOyYgigp
nFCVCCUaDdNs0OV+vzjWuIfD1CUnldggZDMcvqR0mxgS5aFCjePvFUwywW7nzGfEUXLhbTSFjCd7
BhRwTBl0nDK37OdJBZtv0GxKmoNW+vKVUWDYFAQpCYPhXn3X0XxA6wwE+W7GTPQY/KWHXQz46iHg
DJsoTtLH80Xu6QcGJT/OSqxrag0jrfOaB7Vhm7dzTlMnunUtuZmsW5U29X45rgsWU01h54o9KSPe
PZBp20xIl38Nt5Brn8eZHanJTRqLTpXEVNNX5T/982LMkgow31ckkAoQylv4jkSbUxfKgOgok17b
lxFIQRAOAMYXqoLodNgXBQOtrDmrSy9+Zb0UjcifjRZwVXU2h6Hgx1rBpdPXrhjHMA9/xMGcbkHr
Yd1cTSfxr4dHo61y46/WoUmLvmDSCaYiJFIWBk9eb8Tw0KPWjpd2KGa7sdhisF1TWEN4SwSeuRJd
svrrt++RBroQFwRm0nRK57XKWGmrkMlVapMEiTDDgrN2Xkx8VO5hpb6Q2TchhZCgmqxfR0Ycjc15
gU6yM5VmX9Keg8CLMWNyKUhh76T4w9wQo/UJjqeHJdYQw6KlfmoiFeMIoswKvLD0k+ZgGRhKpy+s
+AyZsVnn8PY3MkZKHfFC+jjjrl8YojD5hUpQxFnWIJT5TczE2WTAaerlxL/7V7eeLYxZZdQr0BJ4
IEvB5IuxchlBXDJzwlisWbFvoT2uVC3xH2MPaPfzCxNf3rqrzCP4n2iehWochwMaMYT5MnyzXO2s
kWFp0y9YIIJNlOgR586TIK+NzPUGv5UlcrDNhRzVt197p7WXN4FkD4JEobkBkdovp57H+RLBpGEU
7FgCASALa9PjSgGjZBK14Q7WCMV9cJKW/fR/UQG50jqU4Rol3f5iRXXtTAt7SYJxAVbkaSR8pNFJ
Kl1G7k4FqDKA5YZMWOr+cbDRIO48HRR7Fe7CnE9yfh5ijj5FzW1VBdvSwbZdBekBg+hl17PZpYHj
3JfsTku+VLUCpt5FXjPW8dpPYmdAzmhU0u2V5jDQta/lR6s39EP5e5t0Be0x+ZVcQLCrtyTk5jVz
fbAlr985f8W2gAOfIludjCd38Sp9JoOgVHe5Upejru2apkseaJAT0EiLZXW4RVPMQEAAVPmA5yIY
+wHBiNrf9CzmfdIF8RWE6X0Uoc3cyJIWa36sSvrhl8niKxZuyG53DgzJWiSqqOzQvcTAnzY3Wl+X
9Pw+11gffbXSMXBRlV0PF0PnP+tX+ySmmDNvEq/ljSoLL+rpbSamykVOoYbsxJftuUSOjSMqb4CO
ntpmnl/Qzc5z9lyYpmszzW/69G/lallNbF/wz6oOpY/CyQWNmnEW9vtWNiAqhdyL1NmyrM38sGVG
/kZHlwk2qpPq9shezCT7TyVGAzbGt9TBE3mWJr4mqMsTqjZ00m33C67zsLmXcVYXMah+178lBq/4
m+JYxPnhynk6k2ad7OgKQK1HV1YuIHE/8IG7b0j5gpjCsCLzALWJSdNNJEnfyIe+xbYJVdi0xn3v
eSDJcuLnRUQ7vPil/qqLoFJdEuRwzszwkFTXLUb93zmpiRyxuwQ0VZAW+HeY21ni2wh2SNLDADot
1co6yBRpJUY38N8deKAA1IJjzbV/TM1CTQJylyyxv+UYJEnzKcIuzqrlKRT9n8PshN84CDmUMPaW
R0OWAeQxao68OQaTwAtuXF1dIMgXJR/zawL0pVn+URaHE2CYgYL9XdGwUKzq224rHfHSOxreTMIY
ifiP4OaF0IITpSvNQrcEQ/gLyeul/82OnF4KKMaVVNryG5KEyzVi9+mqHDG/es/Py9YCsfyCK9HI
lnlzdfyQJNPVv/+hnjU6SJnnyTN6FGf+N6sFj+Ng2FBh30Ms7/JLf4QkyT0xQBsIXCka4C9JaA0p
heh/o3HEBueKpPNudlfBCJwl7ekWq+Am/mFgwRDSiFT8o2OY55EUeH03YMJQHHeilKvVJDWugTde
+jf8eNJMUYINSgqMgi7D3f4i4ztcAjbNc6t9qfH+dKiubjsMdsate+eH4KgBwNcw7l29gJgodwfp
A1NKO11Zmw5lBdbCit23JvYAy6l/UgpdDFJr5ahr8FgRKTnegaAtAt2NlbHYLaeM9S9jinrXHWG8
3GOoDSA7JG2OOxGW2YWIBd6QuVuBh7YytAUBoP4+LaIZGEZkl8YUJKJLRvZWkgKGeE4guRskeXQs
Y05+HY88XoPTD21QKk9/fgle/+TkGenDAD+hbq7Lgze7hWHEx7flzO4FLrmIIPACpnLBalhvHsYV
pHPGA72InrMt9E0h7tMEERE5m0FrAUndqbxxyhVcgWkNl60ltKmHsaJ8kJj3JG6/3eY+4yxgo+ox
LxLPNPQQpjOX4h+YpWfNNtpJHN3ojBpJ9umxI2Q+593C5ZCx7NtrRyph7oNMq/G1aE6KwUIa7Qev
liXhzLZF0HdHVdPT6w1WUWmlsma2+snkXdPvehw7wLCxK3cH4gDp8M/npd8oizUB8lcXyRgj/BGZ
CA2anbB8SL6uFGxLtZLHVnvRqdwrLKs6wr4uFVO25U6fUwwVXuZ6jfLaZ0W+7m8Ek2Ct3LH9OQ3a
VpXIZZdBA7Z4PBpc+IE0T5FwYaOvk8o0VktslwRwLGEJrEr/lZN9RYYHDSaLEcAgV/uC1Uq5jMjr
VqvZWq38kH7tENtvjiw2RnxNplnTnmo5kbufgB3Nq/OVdJM6qgofEX9IOiCeKrwhg+IwJfWKVZgV
Yea9L0e4FCpOFEcwp+P/x1KUmBU2rQAeK9Fl9+qAyJCh+heC9VjrLdKKXB+R2ATxhM2IJxzD50dU
tJjn6jn6Oq9xsrwf3XKGnb/ShnJ411HGfrlwjSE1ewsLF+DdO9axQ/2bUMIqtu8I3HhIp6ARJ330
z6lg9O169zHIt8CCI/Gi3RNB40RUi6u0PYMNiCSgT7evh+FCEhq5wmun3UXfFRXtKfJoEBjM3W5Z
nw6J8hYpMTkxuCLplrJ0daVt5GyS2BfMQ9KRcyEo1i4QlAG7vn71NPHSDk9kqxep33OgQdDfvFoL
+jxjGockqjy0csfrDsltWKHYRTuAeGeT0PSewiMVoTifNa5m8Xzlbbok7Mt0vmFdWkzhr/AJiJqa
Qg7zYRavOa+xW+E9ZHh6szeXaqtqQ3WiWSKpaq+rhq5YObXasUcs0buJB2ilVvDh7p3SkRvXh78z
z83LHKO/Nr41+Vgb4KDi3TYA7mizA5FpbB/b2KitVC3Csf2CqIYWDTlhqhjnW+fPC7mIsRY7xDIM
khK73BVrer0hGV1xVR7/7c4Vibn4bdkGDNhM9xeEcyZftCV8vZk1c/P6wSR854iEVlILtNSCVJ6H
04iJMvx/dgP9Hb/jBv3DchwEk/Qh42VOQaOB4yuZjSJKDV4ImgAq2odRGcCeR5Ky6rnHvlAsAkmE
IXFY/MEAhKITX+zt3dkkmKT/ln5h4mPiEIXLY+UHCdZjiNNQIy1sToa8ReRLmnClMlf9ez1f/u4Y
74mgfnEcsLv+1npQdsQ9ZENKYngK7hULajZn13PBQKs8IChmKz+6beuA7oP7whxIplXKQdMzzCSn
bz6LG6QAM81CjqxaVxhOP1GmLnHk3VJ2fxQQPogxSmWTQ/j9JqjUtuq9fLXl2sKiWDlI6fzC3+zY
E0Z5VesspST4JAWWSiHoSBZjFXkZXqnF7QePCUZ0SPLuCjnBnbM9xtMc9FuUowcvxW44dDcozfp/
wNPIKVnGf0xVaBzrdK1oJUqhfAgFTPFR0zKx9fgyv/wBP9M/cB4sVp5xeopw2Qxr3XpAx06VzBYp
bzB5X4pWVgiIPbbZiceUmaYOuCf/5nfUpBhBxThWqoKEOq5FKfa3XXFmXe6L5aOmwIk5kTGXjPn/
ngcnk2VVS3L0UF0+rfaH5e3T5HS5SWOHniLaO0ZPtov9Fmiz8wgJkHxMQsgKfLniZ/mNaEtG5Dbw
YfkVB8NH8hkpXDAEXHbi9wHbw0Qk6TQYzRuKKdDn90OxxFlfQEA/eq88PksRz42rqVs+w7mXAmaH
0RuddOwqdcTr2W3jCwPp9fVYLw38P45rlRvoUpzEqh0BdamMFRmTDEqTQfcWqypNpQgED7rrTvTQ
lUPsj0Y83RW35LLbJuFufsnLxjS+hMsTmDj8D7wh3nuJbwB49iUNSw/L2CD2xgPYlmCzTwvlgeu+
b7CoSHXkiPk9JKH0u+Qj+S+7j+Rz6vVboku7ebQTlry5JaBNoQ+ZDH5+GfT7lJqGBO4gjV333/fA
jpm3IyPGLPa1JEoiUV3yZCYriKK/kH+cxhbp/khHLOCqYqXcVZfZHGTqsz6wFWC++x/Wq6HHEv6d
4xYEwTaHyDEqgzoQ6ElAX6vFNq93kCQnlwsSlaipAXvG2ntD7YYg78ng5PZC10JtFhw4ZQq0vHFI
221FuAgm2E43vV2CvFajbWDc8UpcDQHY0CVx1da/SjlIYZly1yMH7mtjUshOQdzUKiNBE3FSbpop
DdzqNHTSVHtf5NP+iyQnHYXfc/qhhRzSzVp9ze9rh2zsx1YQME3lDBt6U0gNOSPfRpqnvKLFil/k
PGsxg/dPg5J5U6NJNqaLKHnqDlF/3+S+9Vyp96+wFFLoR39UI8NOTg1BB6yHqZIR+41J6UIDBIPS
mFI+D6XsQJd2kTJQZPRA1j2mfxEDzus2PdGpPUTrcqPZzOxxAgdES4FMhFfkEldmMX9jdl1ait0d
CllxlQ9BPKHSMQzVMfvPEnk+v8LcWPUCbuHpY6rZVVZtGmdCXYwBF8y/DXfSh2ZPDP5G+20nBD1V
uggPXVeTaxEvyNFKm2Pu9yZ4nLj1Dhm6qlFRO7rm6cIj4BDv5Z17RF2o8ZtHl85DMQ/65mVlSgGm
LLxqDOw+ZlGjgXXlM3xt3uGreJ+UJRhDxS3IDdOufoZDOzagL3J0PB6pYAry+tm/w1WyIQf8LKD7
qciliZWpffQodts7I0mnwfBxKvBSGtmk+K2Tbsae8hGiVnxWgBqSdONq4kB+nl2bOa/Xlq1p3aht
egpaIMeMtU6muRtC38OhFmXiu9lwrYv7woTD9D8Faplmu06QVIWqRwB2vgnP+htl5+a1zQPO4NDE
2g0cKLkm5bFOA5vX07nuKTYM/y3nlgDkZl7nc6kU/B14aEa0HFyeRil/wjteB24DTwBw4t0MdX0X
5GhLGzwUwyTjbVZFdrFbnARymwH+T49v5j5PbuUGsVxuIorWSu/KhvfiezCJa4xlDKDP7nPap/WE
tXzLTOOxpkKxt3sM7jjU2Zl3gO3mRmdAIP8Y65vwQGm5WRJU+1Zg9U8aZzJoc8phFX/j2A5bmiDP
aNerquu8XmYAkAyxV3owU4CCQHv1e2VMBOMvSpMxvEh9O+6rTrrHMerwRYIafhwKDBtyVs5QSdtp
UxelPQUboplcRqBv0CvtWSsrsXRXw8rDGZyPQoXJWiRfPzTtVveEXRrIu+y8kKDjfUsqHbaWXxUw
CLVGn9ejKH0ZaD/d1IM39h3vSUFh9GW1BiG3LiVSfpCq2dRadz0iICMes87UMMy92Z/bD0givyvV
ypembPXPjIVAZweQT5sTVao5vb6P/wlsNvLYZ5/khEQdvkSEakO/At8AdDxVDtnoz23dqwqlro8z
sP9YYYMglThsHx/DM7wLoqhCaBFKMUXAy6ArvSZX2rrxlCGhLyf1yveT6Umbx2LGVX2/sqWSgCSw
HwFHt73ISK6ze4rekJ2oKKqj+mIi9kMY+fEs/SwMobityfsrCEWN/SR3jENK939GyT23RgvUJe5I
P5zKPmf33v5W6YZPUu2iLOWqNTrjQYVwX/uumYf8cR0IErggdDoIlDQ5ovsXycdTogFnF0yFod6O
ENLaAVrXG0zZot7gRmbV+emWGrcPzeG9kYo794G2N47yHEdVIPg2bUPHYgfQMk3lqcCyh2TOjNX9
TC59owtf5LiA2UiQ1a+MB0bpekflOJ1FrKlMTTRHIgRR7RDFXFMNfFbE8J9bddmOm8VhS6Wgq4LL
VZfvhIHmW6qaziEKvQWMgxnNFDvtNtSC8hw9LwzW5WqpJrT8440UZz7FQn3x4BrIomPanIYktc1K
Mmeg4DrrVSR2TJT1O7sWWCYow0VD3QG1nqj/TY/AmmzQmERJAoM9n/2E3hJlApPq/az48nyLoxnK
5pOS2legr+tHlNxepr6NFuBdhkY2i7iPz0sVXZFugA2M0AO3Fo1rqRuwuOplbPVPTDMS0iZV8ldk
2t9tQNF5Eud6aNuHNBZqhn5CnBJrFkfwGxEfLXt56zwGQsLyapdf6xAEKAeJOIBu8gBLwbnAY3C0
LkoXFuYWp3xV1E69AnAFloqBFhRKlguzGMgVGRre0BLG2aCFQL/5+JkMOf7zeUAGjgsSigDOMDo+
FzWsNCmXdKZCePQW4PO1SkQCMC77W9WjNKsPr3SExeBhdD11o0UUu5F+r9CEJraKFaakC9bXTaEO
b4xzHg0JCW8Hcfy+IGJkSEuyBFAdOD0xcXQGc/Bcc8S8Iec4Y/J46dnP+uCXdoC7Jf8SwbJNxPRs
G1QuQyjYhzWycYAGdQTE/+mhIZuCs63qKM7ElrMWUSqDah28xyAJ7DYJ6jk1NR+FT3JYZ2ujSA7/
c+4xIHV3uSqnPuUs4zUXcbdX6Hgqk1WY0x02EsJw0QTwcYUADBTjkz+LQHthiilRnWzStviLXNKD
G875WD5ZI0+qlomyOQR5XLt7XYCg1HOcKMe7CMp/2DKFQS0x51mfN8J8TiVYGgZ26EBaKesx3/rk
Tk/zPtf7Fiv/m0K9gmcNZ/jxQYeXv3YY/Np/e2PuMMBiEot0WW/zOcgkPc0Y3KKvGLkim0Hr6vMz
LsICnPIWIsnBsVp/4W9BZliNDFH6uJbaahWqydWZZYTqqJFSbmRpJYLzOTCIXMl34bFsdLUQuJji
NGUOJ5HNUq/X3L+c41YQpxGS7Q8uBOis9x3eGP8Py1LBRwmRPPAogx4/f8lKz1TSDo22MWCLyyR2
ZrW8S0SUNf1tD7OrzyTfVrUPn0ExyYOHQxXwmOG7UlCZ17V38u9Jlkp7TnG96HWBQPcpcizH3fbk
QVDcc3RFJA8MTfXe7s/7kMxSN0/l54SxpUaYhQDMCmDYFXOMrhLxsbHFRnLY57t5mD2wbZxpTJ0c
HQws5pGM7ldx7XbejfssVQU0jHRr4mJbNSjxcfpWtoEZhaCO7hkTIsDw2FVH1CY4ce8RXWm2uIE3
rvOtHfXB5ZtCAsFLLvUUklbqmGUO44lCakpASj8RU4TdrTi78W33zdO5UfqSI/4oVnYOx54ok7kk
exj2HCSG3OvvvkzA3U911cese5F4XmFjU4xazc8c7cBHo0tIdzkNg8GnNiJDPDkuhX7Eqm6T4mqH
mchYVdTa7149SRsXpIzd9sRLdkyrmSobTNi64PdeIj2ankxpeE8IeByXSq4O+8t8jhlDG2FhAbfs
xiwi60qjRzeayByy42h6e/i6yklL4QrxShTkmS1RjpgdPXH1BtP91QMKka5SLzmMjl75aJGWhfNE
RaDfigu90+pSZqpTw7t2J6DQ3n3XVEolnfWAbMgX8w2Zuh8qVNbPeHTB3+Ke6IHNSSbsWdv3Kp9f
NcfYbW09ldryz4w3i0TcRFV5m9fyDkTw2XGI3WU8ovzayzVMBg2G9wzrEDOGTqgySjKzPVhshUm3
LlTuloGRlwwgt9ev1VfDg+kUGZBP43vjjBg1t5Tm6uNPhbVRRJh1GFvwYwJLraE7lUjJwp0RxVtV
uEWT3Z0j5yjA2dUU2NRLbXWjOWdXz+SUGsXSb5UlzTT+WEofGXpGPqhvBv4CTJh61LwAHs1+tHdm
lfd69Sy7u6xobzvVMdsUupkX7hEhQkzoRvC5qSVDJBqkLTXNTGP13TpQUZhl74SFcluGlgnaWkdQ
gqLyx/xOlFjMKhzydy6COTvlsOPyXa4s3JZh979eNzQ8Exk6QkESq3qbebp1t+T61l8BSdNFjJKd
0SxEjO9/kjHg1w5GGFTEzQziury1+wxVio6mzTzuHJkvVuyOFcnGEOhq86dce1FFZ8PzWH/GBtUO
6VDdU9Oe0J5Q7b2fPjreM28rRor85hh8OIN/oHB2OdNACnS9pRb90fexGB8STxtg44t3VEd/q7zA
IUy4O6rmtXkcwmzALT8oLUbaADiYtuCovnXBh8FS7YEttRF5pbwkXnERE1Ui0ZbHYjE4O4ObVWzd
HC458LJcPHv0CxIvAIUfiRoSqnb6VH22DwBg3IkPyF+9Ei8/uM953QUEEGbLvUCHgek7oSDdu1aD
arB+grxQ9Q1r434fnCdfmStt43kf1TkVp3Z4tK59eqNgi3/KobHjQbQhptYxNuh8Xn/vunGKUKqY
wwt7kDdgq5cLfJ39bGWbC+hLiXjh80htuN6sARZ3xMkqbIwKhQsOLljun+rcDrrLZjq9/opAVkYk
sghvv0/yYE6AlDtrDM0Y6v1colPfGExjKmMFPUfGrg31oYH/4YN+ZkqAknBBSqQuknCYIXaBxDi8
icABMOvIDIyvhb55a8QnVInPH0fi0Hw29WrcfdiaVU4UoxX5G54hTGxB0A8e6GLkKsKc/r89tLC8
ub8V18nqhclR7/rRkoBKNErwlPd6kwEHu4X9FGci+SfKM42Q7km0fOGKjh109thuccD7vROK9zY5
SMdT/o2WdUOCFtvzO7iBkwbRhiKNIzvUTwbReT0n3oirg6YbtoSwmMJDX2nRsM+Zp6/5Y8iOnXas
q8Ojx/u81eKUsWglTl54c/R6m9VZt99msUHHb7hPkimI6gFx3MCIhxhg2eYXvAfrAV4Gvcmz0L3u
l/hlmXci/+Qy1g4yvmSiKA0drtVJ2/1t7kY08twtz1wEsoJn7OK+Sk9wvSb/ZEC9z26QK4jsfZVg
25M7DlfGl7ZB7CdyMrW2aK11NXppzSQmHgnuG2I0t32KGuTU+bvr1rjnRLnn/momGjAF4m6dk4pa
eMp5wgZTTHWc5vV/b3mm7hk0nLj1V+TQAYmThIVHNe9O4wm5HzXcCNlD8Flvz2Z12u9hnF/Fg/RP
HX9GWeIbgDgUS2faEF1XGstGqUcdAro46x0ul4lP5dGcKyO+CCiKBMkW76LGQVknKQO+acGMvMu7
Y5wZaPy0Jizd4k6FnjyJqBt8a80ithxcd1mxcQtQeyx6hnfQb2RM7XaURl/lU2RmTi5JjL02nSX6
mdbTnw6C4t98TuWucD8SovP6pF5ct81+ryuJZDedr4Zhg/OUwVoAiK02K4HH0tWJh5+nofk4yGoc
RWz9M2gojNnmpy64gyk9XoUWY06HL9xXyn7Ju7xK8vy3Snn+IU0kcky/TOn5ZB0u3IW5c+Tz/Uk4
OV+qGPKS3EVU9GA0xk/6+zQf3M9fgZf1BKyCaWl4mvx11RDal01GKnB3eTksBihhLgh+gHORqjKz
WOyBOWl39bHRhXsg1l4oawWTgCfae6Qn0DoSss7xJP/YR345GD1Mhwa2os+5PbRPr9z4ctKGfjEi
P408T/96aXMJwkftOz+2pMHyZdrsez5Es1PzhDSe/oXbBMkgV7mcugbfDJf2+3dWnpFjgUeyYkwK
vz8NyYnXUo/l9M4qXGT18Ukc3c2liZ9jrdP3L8oqwE4s8LCHTpC5vnXw2YM3iCCkpyctqIVRuEym
Oj0CMLGIifN8j9LoUz4bmVNsdd4ylV6qitPMdTS0GlzBVRu/yord7V5eefgU55vrWVgpxnf+qAlD
LGyjs433Osi4N3ll9onXyl+j+CPf3NHrFMQ7ClrRPWyCIBCnhbQC84jK7fkkC6J0ghPNjtWXhyFh
CCMhx+2bVNfHvZdbqwwgRm3zQSE2JAtktCXb0xCDvCmdYig9wFNejQlmgElxu75rf8iHXH4ZFBZl
Lt7tPPYCNQ4DNYYIrQddDkGeLRunExOPVArVhs7ENn72gIXsGhcRpTb4ry9PyUkrdFZc0aqpzMM3
ndvyas/FiBDaijf3NVZX3AmlJRHhjicUMWwavTmz1/vG/M0cEkcaJUUbFAnk953r9NXk45LuK1kU
rwfbxVTohkxXg3tuZn8A1KIiVVGSaPmd3EyguRacwxkZ4LItOmT3ueaU+pbLR9lnfQLR0+pqswdP
L57hnymlVwpfjGfwDBUMAFq46QuxUV/EtNFPUpYSJtDXkFzWNlD2m9UowhNmpRM2qGo4DEYArO54
xpqQ9eS8bb/62FtnVV5o8LavXOn5C14Idx2ZLIhregNU/SFI2OqThRWfQNeABBTrWvH+oK66got0
DBkkQd5/mYJfdLnYCyPICiNg9Bmh3xZbMcH5m9t8mtVk2+d+7SrS8KevXdpoGdvZskAXFpY5uGeD
kzaFRnLQUV4hyG8Bic+ykJkXj4iQikYkLIa4j3zlZxvmmhTM2zTpCP1XcSk1FFGJJL7jARGY627E
Efyj6gAhNziDOLwHY6YSBn0y+KqdURHFaG9Jlp+7PMbNXP/EtzVlnZliIkkKzeCqqZmxQvzbzgZe
PwTjoNGF/Aij0uQfLu0wxfqI8b+vknw4/RrisaY3dtq+PxZqJuObn4DaxERyJCyEJ212WQ7djuCX
hit1P6KvPRqAgzbW0myAuiDmSl9it6Gdk0fk1A16ISjZIqQla/lK0eZloK+gN80dh4csiSVM12jL
Qg/I1AhEVQeX3zh3FPM8HhTVFBy3jfL+BN2Kvy7kkdcvJs/vQWW+MM0gWXMfBRDrGSt1FkVhAWLz
iqDAbQEugcfkAKCl4V2tuSx6YLuCSlP97s6O82FlLyaM57PPLBhQKhuq0yN9CWlZd7g6LKMzq7YY
oD0F67fRb+7gtfSUKOd0JwPi+guA+3GY7FPuoLq9I2QMhm1JN7c9STECmCbM3dfLx094LyuVpaCV
FQk5cFWmESS/J10z5rkmqdUJfll9HtN6PVHpVRmfmldH1Rbn8jADWPxXWA+GZ4MD7GAyFO1+ctrz
ReGghWCz5W947ti0h3lRsoLPltpQwOk0IS5ylbeQT7ObWVmC3rLXF25/gCxb7JWW0in50pXOLC3h
sCQR8pZazNEOXY7nEE0CEZ+kx6elR25ZE+/Ncrasvvp3BRYLWTRIFjs2D9U2CCGW6ox04dt4SYTl
aYNWW8QUXLfEUM+aH8CFuZLiCWIJH6jByF5RV3H2fov+SQlGbFAbLhgQCqouDX+MAfOJP1VESwJm
UBV6ZHQpfBR4hfvDPfBXJxqatvCFx2kuMdrCuqSYnhRe52i66tTEZ5llQoKe9mFt5jl3jCXODkMt
nnVLWPwojY01ZRd9y5PC4OuCPVY9y5nFW6aNK8N9Jf2X0c7biE4ZtO1T1fNIp/ohaiA5uLKybEvZ
XfqKwvg7zi/KSdWrWy77T45JBwp2Nm6tX/VtsbzX1BUUVWbeY1Dnt5Ewxk7ndYv15r3H6G1oXWs3
/AUuphPj6qh2o0OzdfFo0fuhWXLWUTPPD+CuVxZNk06thRa6U4UHUecUCAZZs4hqXqAACmdLsAbr
fcYOhr6tXBTEUkZIDjpalvYV05dX6FOlH9+gacozops7HYsvYh4sxNnKhdnsv9NSvV2VxrA1KP0g
kJ8jCyohzfTdKxcwdFdOImBMDQaAc6c+daTg3kDVXYTvDTzkKk2SFCaNXZzPWbYnC/Hbt7nF5NnK
uDC98JpvsHKerfHJVF+hDvqstTd4O0yiH/h8UScBaxIsZuEUrTJfsri8UzZ69IJRrfBvnC4U3+Qa
HMMQJ2blw4gFRfeErkCbHVQJaNKh3kDtywMKZ+Fxv4/7NE5RU8z6uA/umWNjVR+NxgY9pZil06FE
xovBsx16lJO02TYeSvTpAu63QN6qWOlydSe87DsU/lsZ4E5PgJlVqrmM/KjcScwb5XV0LvaDOQ81
WYru696+BbAXQt9ufjcufXa5gplkExbIDgCzeQnQja1LuuD9s2Ytyrmq3KTvkFe3HB1MT0uohJ+4
YS8TcZY0QBnPrss5ZTBXWfuLGpO2BLL2Y5Bo4mg4xKDaG5V/44PiA3TfbD3ML61MjA2raorKUd5F
LYngMUHmUCC7vrDIbhurtqxuNFjQ8gRRZPmHoHmJ1JrsS8K5K0DCJucP0rzW0Ree1LRZa4th50Qi
PbH38UD686IUlsZ3CNT5Nz24xAAdQ7R3gllNAl6eAhumZtcxSuqDFpTXn6sjpTL516JUaqT2wFdI
E4K/z+61N2x6BPiWZ23Tv6PXqI/BQDTqnyZjayb802N+g3MhixHqYiU2f6AWgBnI6aIZiqhDjdoF
EFr2mSVP2K2ceYKIwiE7LRSJAOAhG/yw0/LoWr1iX6LebogFHfxuui2zApaFSU4HqroOdf5nWxGC
rP/kj7iv/maxoZiZZAbKklXw2xTigOAJzfR9b6/zgwp4Qkwtg3hK7RxmrqGYyVMro4eOElv6t+lW
fv3V2qquSKZtYElF/lu+SB5KCENEyYZrmQGUcDepVjQA+LICS1ED9Bu7AaJXFQHoSSE8hmZYF/04
qmopznNjWzfhLUn4FJNB9wIZxTgFMbjeNfql41PBxVejs2ZLtLqjZbCZwvTqUukxEwszHIlXVmIc
wD9A8+707YIC1aygOcBa1ryzKy3bDLGc1Gk5v620HeRGgKVXDsNLw63ZXQJcrYsh4/HT4FkDiCIf
SpzYAmSyvLhwKVSoIGDMpHSh87uLfszgG1Rzww6xxHj6DSOz7kPUB2DZ8WFsynQRNpy6hkAWDyOI
Yz6ouSWXa164wOeIDx9kbEI2JnUAx+pdnss2sEeJM4eDOytxKJ2LSg1cYYAiDjJ5IwQwdHo6my4l
uQsuwd/v4N2cjs8JEJJamHxc2hGwJuT7UJ89BqstLHDqywusaTEstX4h+zQgVm2tx0IAdBK5zlGu
KabjAMgDXo5ltqgIwNm4NeN3QmxKscSBkAPUlTAKaMOuwy49SP3TZmXjI2EEIVuwebpYUASSaUeG
qnWkZo4BJcejblwr5DOiFCtP+ztOA4rpiSy9d2Q7ojuP6y6unoGtdo+Wqy62+OujjXuD5Xm4l2SE
XIU9kcgbkQrtTbG31frWsJJ6H2SGF9yBQv4t6qVZfmKQf51z3K5aa/5LHlsvYZl/ms4dRbCpUw7c
9L2wOpsGqII0w91JoSt3H+tue03EU0w4MEJDUPUHizNoyf/JNx43VKDo60xZlryv5zKMyft6vPVC
XQCShLruqd4gM2Lf/GiT/fivpam6mxD2mXWshmO3UKOCro2RylHS96mcIMHs2N8TFo4SeZ7FSzwX
lOUfAEb86UpE9tZ9m6PgXKmJ9z56evUaqhbKt+LLMhwkAbK9W2riRj+xaOWaRVIfBhCxK3bViWV8
LDq61G9pGQYDoyRf+M1atzcAqJlnlHYQDXrUeg3w5sv25kk69Rjq6puGKcWaH5b0VlE1O4slf8rT
/5rXmeXB5GqQpWoGU5fsZJWiD9fmG7MN6YqaNA3sKKOQTDDGeNLDZasluQSCtFD2HQ7Oo7chZJ6T
/5pCMwr/3kkdHnhDUmJAuZ7NszTOD3A+WmQIxJvpU4MBt0DuUpeKCclgukEGeORNKcdU2VQu71Ss
mt5Sq043lL/J/m73avzh8NIUR14skCUqHtgk5oxrV2rREsX0iZM8CajCb8ahAJW6vmDVNJ39kUUn
uIW+v3FqXrucPIg3XmISdmUwb+BKn+DQryHYe8OFyk/8m0vFsox1ozUo/4xgOSPqqRUy4bvMjmn+
W1yrxD+PTaxlLMr/5Lttf01vZIj8RSyt1K+6xH6pYXsIlJPz6cVKCwKSKPdp91bSXwv2qfhdxHtQ
yl86B6yZULpadE1f31IrqPv5ZL3VHsxPNrO0uAKrnRBgeiScu/hF68eyReQPnXeQsWor1umUXxw7
UN+O9647iVlMuN9GHmon2Kk0Kt+onhjWLFNTkQS8iLyJNjp2Cj4PreOmS44/gIwstSvfXXQ+Z2R0
HnP927a6IJU9C9bV63X8vablzrXUx2KsqXRyPluStI7DZ+Bfiych1f697GyZLzZd0Is+3uRUNocJ
FEBLPHopuM/brV01jtEW3BjLkLXgfdo711G/ZePvv3DEGSn4fhFfYu0PhVsdgXYYMzfjSuti10yx
GOIyhZeKoRrZnZgvtzaD3FVneEklHHveash8rL9O+dme8RW9pBvO9/RB4mrm+fIIRoVyE8vgZ+zu
cpEbIMEG0kXkq19nvkV2NoBtdnS5ee4z4MtIylK6b6cxv/Vkg87EXGY5CqR3XIyW+Yof9zLmDKmC
IzSqvxT9Vb419BGMe8ds6kwMrv3Wa31QyUkvfmmen6xDLIFmInL+Ou1BQlRzBtUvUhwHDt7X7o9S
Ih75161doEmMB1q4mfSd9D7eIh9jrcOziM4xe41PTrRGDj7XBX3rf9bHB+S5wNkP5KZloyCvBGXe
NO1ElFBxiefHE4uAiy/uiO8t9jmc8sDexBNEg7Gx9kf/TUohpU6PdZIMAMK0mq58mIivYoKanXNC
oc7GjrIweB0d+GAhVw8x5N0kPH+S0VooOKrdsbiwN4Jpg6wiFpJgeKunfvoAhnE3zF1ynOCffHLZ
1nYitXJlvseVLfvIxz01KWIhm4seaGJkvBXuUcyomDCAcVMG28Og+0wCEKn9t6hv6wqd1MMc474P
6wc1kBcyiiQfjAAVbfEQbqVoFazluxzLN2rztjp/END4vlts8TaAnCIRDll0UKl++/l/i3tumUcU
mKmaVpuZ75ONZJydY6WoMdPyJd1iB0Llh24un9Fm86CpfI8VFEzURnrjF9g+wOaMNHGbAYMek3IM
Qd597C541UpcQgX0jb0iBQyVSqrPjqdsonbA2s4SisdfUOSxuWcpJGtzYevOTHhR7wCbVh0Rtscu
YZJxogPKJcpaGxm6FRCiYYHeGCBkUnFzSKzAc5wpgZPUxAeo/Bx28Yaav0SlFM7AdM5TqOUY7ybM
iWIP+WE6hdVzzG4ay+euorfAJz+kyRFdVWgtKNepjEy75OLHltW5at6QVcRze2hgYwiDYtmexjMg
DBXHKcUbcplTN8eqRi7UgmSFGXuA7bCFngUlXuXnVmDMuaU1pKh8ytgYaiXyfl38DLz7NDNAasLQ
bTrk/w9L2z/nnS+ri3zTHkU9cHdau8NknSg22fgVDcwxrmb0/HAn4iPXYnUt6s9AjVBHEUxOfyPT
wzpMBA9YbplKDOUUqcZCo0ZEx8MsimnX5KynqbVeTAsCKgH0PHNkbwYuUXCsfZCC5PEWytwXUlD+
CT76C/0NFwKeas0dEtYgePG0ICLdRT23qm4/4+1+G3zn78c+/PEUfZ3Wd6dj/nH/Xs2FrAxTUaNl
srbAH8wx96jxBHOvObFoBJHvZasdpXlmppKAwTJc9lSiqdOtBvGBynoMC16VKueTOmJJX0flpyet
OpjFN3DSHwYZwU2Hy9lRi4OsjrrDCjUgPLQBJ6tpAcsbOvMn0Ul1JGYsB3LV3tOyhb+KR5JOAqka
a+VGbMYDyf21ApH/baj8cqMeb6CJaWMsyLooTZo7d4qA6+brs+F464RN5VZ+JL7UCa1Z4k/4bzlT
heZ3CCUYPXevQGQGDIAoKoZ0PjamvyKbc7AUUQHzw6VDn4FrRpZiC9wV5Aiw0zmhfg6zXcBdqti3
6YdUXCmMuMrRPw7Idfy5Oy/94aJ5OqxrwYXvwMwU2NAqameMzo+ImxPM9yLDzK63ImsWkoczWgLG
O7BNo4zhFPFoEyvSusNuT/9qP9YzpVm58eltCHv686Vt4QLFhQ637olkVtiGC6bBFhSFJ/jyskss
J984L9EISES4Ru65WbF7LugfEghtF7r6le/CJaid8rkwVeehxq6SYWc9tRoAoZU0ZWN9UTKZKJpz
zRY/d/CxUCfHy54tbH4jLL7lFdEIjugM1MlMydETWXjLYdxtppaKlp5+Ew1gXXCTdMAzVN3SqXHL
ehICShsrZQpGsjSjosb4E0BrXO365gLmGCAC5K8jsV9Ava8UKl+h0Y5RjP6ywWyLuR1yOnmiba8t
G5/OMJWcVD7H9SP2ybbagT5zs2VzA0+NJCRE9XvKpaInRYeXfI8HGKOrpHhGl0/H2ytLzK82hnSV
GJX6+a/YneS3D6OQrSAWHOcxoWdBto0Cv7uaN5JMxLI9IBsHsNjrcDtgHGXkHfZjZkgwUDlgBQbU
EcjZT04fqMNhMHqexqocrKmYLUSGrJ4Fjq4rb9L4HdfZazlmPlzJQS8g8h6c/2oU7h+JD221TWnG
cASxEPejUqVN2yXzuchwkmE8q7gsNXyI93gsixgnut8CjU0WgqM5bsZatmIk9+IkBoH3vSoZ9eFG
BcQk5RkJXOFSNDr7TeM/8meRy+1Bd0WOzGjwrmYQpxLukQ9ho9g8IvAowOpne0wlFt7pjwZ94BMi
jGpvuyTi9ODkM/HLkbbUNxo5XGE1/b4ChhJmnUoLLSjZnUfaZ1bLx0LOvxQg/kUdhQaq8HvqNE3c
r40k62/XhJ4x/vHaiGFouf1j9otgvj8jne0bD7Yp2VrL5qS3adbeHqp/Ga+/+0KiwWCtkX+chgow
rGzygnoVM5ztfr2EMaVi32S6tqAF5YOKEIRbaVywRcJySQbdDAt/EV2rwr/KHpsg8cwXg4ISdFDh
0/EOkhZMMlymnJUX5olwCdfk2wYKEqLwvE7JblVrP2OYElZwIHnpUGmXazpgD0TT0d0FL1/d8KtW
qluTiRNJ2iOvv8RMV94cCBfdVUb36eO+gNl/juCh3ClqGDwmsMAu+FbTQP8B8Y+BIdZibHqFZDxF
fTgnc3izoXLcXGSgcTWfbaB51Z3hgHXnq0DmtMA6EpHLigbdPmED3+W6lV7zgJOzAzbuH95qoEBb
YuDqHEjq7wTpJwrguBxXpa/IzSuylWe/8YHrJT0TM8vuh2b4rcJRr4y+U0aH+6QbYlrlBjwpeSSp
VYjA+/nCyyC+cQ4wlyHQkE4BFxFtpnREWs0LOl64YSxl+8epQiIWO1EcicCS73vx2iRBPGdR4KDo
cSNlU09YmVTV9iqgXfKdyzRcS0AQe6mHWhF9T5Os0fE7wbnLFg6SLWS27gIIDn7FRytegpuDiTLZ
wBEbpTfXa5AnK+NqXgqt5VnftDIYB/NQm1HVcg8+4kqbVa5qB0DQEmyWqKhAbJj704wG+0UCFJGx
ekwwOlnraNmG3MSSL+4WwnTRJ/9508QNzbdF40GefDlvr5S4na0gApX4b/DNpL33a84zPFcZrahk
WwC0Lf/lVNUXPaoYMUKj2SMzLo9vddIHOrVVTFKiqSEMEY1F8WTzC2KOOOQWPUiO9LTOlqn31L3S
2SxnKnn4P294ufbzjRvqEDShRJGAtoRuCVwUNLnwLMCUCjzUvdeLxxrnXrNS9NIGVCW7O3FqsGCr
Oi8AUyOBrysKjyK9eR4plmU9Gw0j4silOBD+2o3XkhUuqn9m4sLWtpl/SUmfeM8Qevl3O1K03N/l
xOiU50OjwlQHXKzBHIvBYKEqBCBWpZwtRUKDwRK+7GJ82JgsXWYRcYd9Jwg2iZ158XK/mVyYbbH6
n/4tJC3D3lSizUnqIpQmjpNiZa0kvZXbrNvyzi7pdP0YaWEs9qUTo2fXEWdTl7xhvfMuig18W67X
WRRAgHv+9Z4PcTnDSKirdPhfK4tx8zq+OYVfg0CBllBFPGuWUjZF38bsO+K5I/pj0nfyWs2eTpz0
GSuHIMHHwcq/S/wODECEIOE7qjQRop3hCFdgMG0HHa2LUIW1c678Itgp6GQtPaoN3VHdUqBasqGN
7/L70Uk2Z0JuonZFyEcVkLzPwxCyVhWbNk8hKujytwea+YUNM8bnP6yJ3b1tzzXggYqdqOtxMs46
lVTfS9N4GkO2S3xrC7YV/bV+r1geBOmvV2X+Lr6FdN1JyR5GGKkhWD1R7bTtumSu8WNCsacRa6EA
TwapDMBps1CG1ooxlaEd0sXWYiDAS/aBv2PDRvCCEsqn/dhCwzVHL279nNwR6+CGwY2f+xjToD1a
5zQOuBehWKfjNzbLQiHa6E3DdrzEJt5qFV94w1Ew7suUFsgTAxgEUoUVbVOp+xGZ1Jn5chA9Dz+d
CpoH2a6B7q+4/3QN2LluQIh6a1zYwAuC3ndZJgWmscnjI6BefPtUxmdNd00JlzRwjq0rbuhHWcKz
RM78rzZGzDoQiHcVBiEgQgYHAZ4t99o/8Y0txWEQ0gf4GKnk5soL0aia8mVBHeqPfcgzu4kBl5hk
tiuBULPAbOLD1iCoFrA7JUzM4DXeICG2XiRxjh9VMF+G7VB7KemYfWB/ZPXclxmAAFpr4hMwiXRb
DSRSZuFwQWC2sTEjE4qklNROfU4/OJcNVT2baJFBAePjRAa7yy/tGAUhc3CIQbnAUVLyO5vBW/83
Mul6dt1W5QFPARjBw8El1Wc00/6ftLFrxIk+iyido9kHQ4zWfZ0MieqTc2hyqPKsIax1yRDQtpyf
g84l2PgIgWdk8hvUkVScM1qohRXXWuLSKB7q/hsyQd6wyqd5ir8sZKwLJwwAq+Jk20qD/5s/TCQw
4zw2PVMDhg78LhKfcikSttQHZvl9C20RZ+Wb2Ob+2/ONwLZOsxEHHo/0pzlMnPW50VQ0GKmQhix8
zJ90xoIg6sft8DuoHSA1qBFIkGWD2SJsGdydZtKNoQUYdJKsYNg0cE2DUaZh8ut2/UARqVYLjA3s
Ax6NrzvXHGvX4Ur87ppV2UcRKjBZ1gKbFWYt/cxGCZpJD9hZDkQOoZ/jbbFakDbbi7/BXuC3GSFY
oPgiKKwK7KHlXhCdZHjXuiRjMIuSnWioJuCviKMmMLGvVm0nL4dyZAAe3wIIk7LJCHVNF1LUwhT3
RLs21/a+HBRG7nrND75ezr4DA7k3Z5flByaChn8QCw1CP8hGB6kAz5WGBRDQU+Z2n7QiBSwCiSIo
2TsxBBWQ21ABe7SRcy8Y94fNcJQRC+j2SAedOufinx0i9x8yTjIITeOOq3wYWgqH4JdX4YvQ++pc
/fzknm0GfUfzJ45lWKfWID2Fi18NlweFmkK+nmsXWymzfxYpaARHSL5TKAl5eAzbydSqgfd6I/ow
KUNX5oyhxXNQpZ2xKPnuIbLBT7R8GON/nddG0oKErdCyowXtfqrFglvDuzj05d5Ptw5Jb6aGcH7U
2+8Eg6rFeXwAyNhxVLJBfVd0LJvbOo41f32CeDNuaytnWv4I2Mvk6D1TAhqPfnct26seHmy2Ski8
JXuf7aEwPxGMwtyzmgeJTnrHUQGG+MC87jnACC5fEVbgTIWAZio0dsimdgx9bsi0nPKPuzWnCeke
Ds7mr2pXEYeDK5iMspPVlheIL1c1b+m/03sf9pKZraSW/hcBLr6V8r78dxYxGp3msbywFQpN4/ES
UqqD3jt/XOpKadpllR4qWX1TBhTmhmSKDW8JRXfN58NEwdMk4ZmvGO099xgajMBioaCe0H9/YJDS
4DiBPAY98rFQdOe9DZ/xKHbCyxyniyM5JF1tgCmJB0alaZllrlGaD+N/Uc8EUVMXSt1dcaSnEc/Q
c1yUj2lATvmzemGJ6SmrgXdS1r2seGJcvBaos0NeY8fA8l1BvNx/IFUnO5VJLnD07A+yDp8z6T5v
MhvthKLwvTMDQPtuxfVP6szTfG2jUkugvx0xrmaeqUQZnGQMV2HqWVtbAdycZ8ZK3bRaZPc3AzKW
YzfibY31Wmw8XOPzDM2F0w27sEFDMVLw/UYKGuEX+lzrMR3tz5GIdEgfxSh0XzLAws3aLB+oW3Kw
wwKu8KQO486v2b0Z3mMjQBfiWNLDA9dO/uawySz1BhiIgv5kcATGzF5p0hctAMwFpRS5EpxDLNOL
9Fz61FxcLEwy5n553BDCLfD8XYxOmq0+IFRW0lLosEbQpIn7mAf8+9R3ZQUZWzvbst/4ZyeNxcQR
FFmoaPrBJake50x+30Ny5mNGww9Um6FxonpDWtMDyG8shJy3n+g6Sr/Xn1OXmZu58m3PlmWfOvTT
os/5RKQ8Br8Ezx988ylsv3SMG2oi+IVsTiUVp8/hmUOSKdLEOr0Bj5GvAC5nhEV9IDdJJ2pY+6UB
rIqLg3Xdy6KbzhsWndpN7pvKlyyzU2Q1uuLrs2ZsZVaLLtZpuHNQVBS4TysFbq4GatSfm8vzytul
kzowQCvNtTnqVRUaQlboqnaowjZoj9pJp+Wf/OuwYNdKfHBisRSK+AmDhK1YzNouHl70ATqL1N/Z
wYj98gvAv0kkik9dgEjpWwWPr1yQciCjT93+zNprmMYfRm+QVuXwO00Guvya/MHC2M6H5m8mVAr+
kczg6+Yf/llBWM2R6XCkslTnHnxNyg65XlTYh3dqJwKHyj9PwXJEx/IoleKGDW0Bw9aAOT/H0aqP
DEgBrsecFQcCz3R+K1sWjaD5ziRv6X0JLqWjx3oxfo79LiyK/MyN7YgwRE+G5huPtxPQgucjbFS9
DIvAtsPJlUxsHj0PwBdjcN6aTBG5DYnwBw3JnnFqG/ZNRkorZkcG/LHSULfzX87AtZmZHoDOTq/r
R/Ugbb4zOPEzrdggU4fCh1HjbYoNECb2/biOwsZYCavFtgxYFYQJQsqf7smXfuutu4dPGO41OFZg
DLF4g85JMeI1Oav5OT6HZy+qvWG7f48nDeyu+2kjqy0WaU094ne5sQ+9WXwX23sRCKp6+o1v5pXr
YWE871lXRqM+BiCmAFiWaboICfRXN9zRnvSC2vVTA+vLFraZMcMqQ6jkfsGCA5IfJ3RxB86CwZ7P
x//kskfz8KqE3c8AbEuNZLo2kylCAZqAuCNMX/exvsxXVqR0YUUCfarkJ32FfN2tsgIT1l7jRi3j
2vpStNaHPvY+tP8hK4JAQL4XEJKfU1F3kSNEf0/4vN0BOwsSI1FRlfw27D5fnV2ks935slaQ9C/Y
wgCBloPqXinQGmd0myCupEUhiLQS0cKk44OE+1YfCbPScGHTY6Qf3IbcvA90rIC/cFN2yqefzJ19
gzy6y+hiyXNbJaZKTvNK2IDFG3zCNxwOkm1OiYFp4MwzU7RF+M0Acx3DI9IJVCBdmClTzhyYWd3i
ODAO7vfAJkA5Aqn/B1nAWPAly23gLVrldDK9Fhu1un5wMj/tbnjlLc5XT3INFY3es0iZi//fUBLG
Z8SyOxwvkH0HVBM+g0e5eovGWYgEOTqZot+SOdM445mHyzLLHda4xdK60w2b7+HKcvxnO6em0eYd
YtI7ok+FOr21TbGNFyjOf0XbI5inQZhJH8Hwt8ArDAoGBV6J0+RP0KGsOLrb0qKsK4aR0SgZKmB5
hqXWmPeu2J0thpiDR3Is2b22r77pvLb7IfrpH8MveuWLkM5Mf2PqWn9DWi08Zv++l0LNc6fQ9kJz
lGuFVBPaotQUQt6BZQlOeCX1r8HpjCn1E111u385Oc7SQ1m+rQBckuoNVn2FpA3At6JJtLSFOpbE
VBb5TR9hrOfvD/r0yJu34BPlqGhjqJ2TT/bEfg+BrcrnvPWO9sjeuhwu8I5nyWIh32SqDUIWuIMA
vGO+ZOfdmjnuRVbe/Axuhsh/DzBLWBnnsUyEYiN86laS0mth7Gn8FPgJ/H2kjwP+f8pccWmsKywe
xedUHMDDkE3cXkcYfN6352+PAugAjs/RGYSpifTN/RrVC41lfEHkzp38zWUhD/lysJACR8r/GiOX
DNbZoAvTTXp4a2u3hCN+fQJkJM34VHXezDwINLKAsG/cfSHSVuqeMNB7kOwjEBTZQ3CxChCJnhoW
kHP0cBr+i+St6EbAajo4thXxsxfC2dyW5qSildludCS40iEbZhQp25K5Bo3wkqkUSYhV3TR2sycy
U4lGWZutMSDFG3l2kpkpYgm/guc8EXXDzXtOS0qJ4eZMvuyBa2HTdQ111qUB6uEbFu5Kr0a+OCXj
XV2ezPff7rPfSwJgc/zwIRgPZxceS76jZPhC218TcRhKT9vvDCQxzlPYhh6gBKa815Hv/wooJICS
zOF51x/79WIe+Fxz9Gn8fcOiIRLMiewWn/jX2d9VtCe5MBNx7G0zE9NrMQyXk2M7kbcec+qIrvJj
0nKgWZHDVBKp3IXsbqr+G70aUqyVsjkb0BIypiGkyPOov8xQa1wmDZXls5xsX8lm4UvOiLS9qQSw
24y2QQFAD+8yPuIZlNHT9BRKznbhnpFDKWd7ToWuOIzRRn0vGEseEtSm2qYQtFkPIQJeH3v+ezNX
86J3d5FwmFooQouey3YMzNVs3PadNE22kK7Bhs7dYZAiEl1Du+TBbT3NvqaN3HUbfckH8RTCOj62
x8sDCEUhL8wI4G0iYICaRR0rZmp1pIqNaxUEmmQcmoocnty5xZUFEWHr81IrRGuOkUugXjdF1sJj
/DQWPM8LTDVi0tNRtQEOEK3oonsQbMZibsRBov5OiKHC301zd1YIRvUQScNOd2QdijPLeb+auPKy
9z6sD2853lcsMQRatzA5WIOgaA/hne91uRZSXsWGEuRmLYN+b4qiAnsZ7+rY8eWsVjsBQ4q6750y
v+VK/HsCtfiNPbvBOT4P1sFkCehLy+hXPiCocY7ZQgWTrtRFyHyAsrNqCJJfdv/FeAfE1bTh0bKX
WmdWq65sTgR9fzGy8P+7ufHPEXJ8JMEztmrd1raIpUAkccQFxuxDLockiwTHAAZsUl8eNUHzZP/Y
+qSpiSY7NvUY/06POgREeuD8MVXKGbbcGdg5zG70QOFmbuhAYZZA6rsr58R5ssVzHdkpMZ1dWJtP
BpN4KoYtRiiQdehYc93JqQNasjZDx9SHdPpi1StyolmcStnk/xW3WiiQU57T0Ua+XO7in1BgW0uN
7eqxNaFshRRepA0wTO8nMLv6Kt7HGmtGWmg7CgFVslDsV78I99pjzk2wjKAMAQf3MjBo1bSp3kNa
fnIUVIeEoEnbyZ5DkTnbhDGQfAPjthDiu5M6tfuTR/KIosTss6bhAOqn3b1R+AsAUGS7WvINOJW9
cLrS2ZiMYQrE05sIfbsAew9/RhesMWhIeJ5JkhAS8XgaX0kQzQX/naWdoJhCOyNNw3Lm+vVdCSAA
yBcqOKcn47H/9xnHd4btZ6nTIq+T1zvLh75iiJEYfl88/sQ0xTWTlDC9NDkGM7TfrSC8Dq0t+sxr
MsZvyZPHOl6eBSb5Vk5Xo+CadycaMngOkJHwlgyGNf/gFuEgT46luKcQ5A0AyJA0ujoIgeg287GH
5i4iPfXiR6ZHM0Zc/5i/sRP59GudWOZhyDLYKRuA9EFy7RZt/RG51fjinMjBXIkYbfcKnQSNbQcV
RS5eDuseInuPLehUUgmQQCh/QpFYABSUDH2xnYPk0diu7u0UKIhGSO0mgOU5kmFgo1KvVPW+fjGw
/YpDD5fS5d/VbTpnZ42Da+D3HMZLeFdZrOSNJ7XgzKBI0dHJ3a0IxaNcZ76/yclhmFrwiB1Q/164
tmVoawC4rVjd+I3iN8N+obQsNT0GSRCk+ZtNa2d0mpQBgy/3W/dzU/vqurcSAlh864dBvxFgfvjN
GpFs5NyW76288JjikJ1gXJCE3WvOibQorYpfNiHizUqffQNcAKg836omyDx4VJgyQgHcdxNjaZIL
GGBmT8I9xS9jfel700tads4Zhf2K3iOl6P9KiRR2QVJjNHq0Q0bd+/qtmGRuZs+vFD3PznfxubIZ
wbsPvpWXH2E4yPf0AiZ+ZSOWhDRzLNBtLGkFaKB+bQLkLEXsTpR/CWah/sMEiWa+nh2VyaEhuqkq
6QVc4X/n/vquCrPUMsNOvvsL2aDUj6myhErFqqkYPpFUGtrwDGmsjh8G002SEWKw+vh6j8H0HI+v
z+eAqxQC2Q01KhU4Jxc2Q52JSIpdsYGAbT/La7+lBmLu6K8HEUNnhIrO/CeQj7aJmNFI2p3SdjDN
nB5loMa+XT9yxMJu5put/73+VKrJEBZEy7GjTIhl+MQAdXLzpYnSL/qzuMipTmZFyr61oAsgcBqR
TGTKTI3mIz1tP3ayn9kbcLzQHFXpFRyIBeWKp90Oq5e4E63rDlZB+gzpMILi2HgQxGwySfKtoLOu
QAjl+WjFqp67NH/yRQC5SgUuLPBqOHVUvNwI1Q0lkfsmX6NOC556Idp2Szb32pMZpqbVCBJxwLRk
Jm0ZukJWFQlBDMVKoG4X669u/o+fYOOp9oUZSfKjSVHQns5yTj0tBf/mhJ8dm7wLpwUe1hc+mjL8
OYKmAZ94MB8Ho32xHxQ3nIsadrFQXT7+QQNuvWJpvUgiaYXT7zIG2TcooVnnvBt6R1vRPS3ESf8X
RT8DKazLI2XagDGccKrCBh/XV0KUNBi6MULU3NroU8r0Rw3iRnAkhUWjVApUIQNATE2wB1odZZE0
4OZYrNQrjS4BeksHdLBnVgPKKjNlTuvPPL0vWmdPz6lCPkhlucA9hzsdWNtmFZ+klgRr+823vgGZ
Mxb9fB9EOBZ8XynghXY0jmQL39+89I/6+tscl35HyWQylqwnEMkTyPb5ZJ9eG0GPd60f/Dahb5Ph
R6jirtYdZqtscf9I4RAhM1REKfIpTeohsKxaqL6uKGeJM9+Cr2RHBHo8cYA0eAu7pO/haXyD7i6F
0UuoAWKNeaZEU+AVyCkuSvT86308KM4ePZf+OTGNXE9YbK3OiJpj72JGtuE9dIrUx5Ib47WYDTHZ
corFY+3dBBpqaviThnmyBu6GWujGr+Srd/vY3jlvXbSA2KQTVAcPU62LzaixufUIYx3Nb+Kzsjbz
7RRiTmcUH19OddLOKNNE/Go/9EXPiE5737Zf3mXrpaoR2DGet8EbTbJ/3M/q0C0V935nP90XRqJz
ebPB4AkISFoPBbNDPLMqY+USJBLfc+AsnuCJIPakPUMOtOmEIrr79w5vFTTGlkNbr4kjHvACdYEu
cmBfBE0wXsK/T+qg/+b04cdVdxFrh6AFd4UKs/xQonECQkwtucqjqs+t/a+63rwRjvjh3I6bYr37
cckYhhnP4iXPrW/s5HsHxsXlOcrSc3/i3OH8bvzVWf+j9FPjLREcNccgvpM/sCz2r3F1Xnj4i+/f
GhaQ5oSNfHU5LFLF69uePjQrgAaT1FH8wNmI5ylUEBKMJS1Xt0b0PKU5Gx8mQi6l84mdSFSGd/yc
3bjtnJ+cF8RXf8w+Ra6yr8wGhSEWVNg/TSuoR68Y8scC1SeibrL2vX5e9nuFaP6sHYNSIHEqPnFj
NQJcaF4A3A1D6rv5ey2FuAd29zfUSxObxk2vvhjeGxOk4oWB1xMuz3zywY8P20hwoMeV2xj4DnVe
IyFfa7YDNNKC2OhCaJVpmIaf8PtLE9vulxbFvpyAgoUd5+wx5aZXIF/taobulGPyBCqqAKZmr+uR
MYKg5hfeRjjzDRq1aMdgFSkx7s+G97eknpyCdFLL82BWS9eIwcANQPPo8XTIPJzrpr2WkhbeEja5
X8MSDvOykYENWFz8BKv0b7YzTtR5ffG3SAeutDEGfo4SUHfQM3DdWT4GeZt5hDuYPN0quHvxekS3
cSuGQbV0BHrWroLxBKqHKAMBc+BB+y5wLj+q8KMsXod0pdOtnpSkquGjKcaVFLvz9M/H0S3h0wWg
3jVWaD6uGfL7JF6Cq41DQc92UBECTNNl2yqXw95eVYOV9aUtcZsY61qCX+w1wX4bC4YrQHJAT6AT
ZCE52tBXdC5XyYBYlmHYd6rB2d6pzwjDXewxHFcq1XWxLF2va2OR2OJbNCtOdoIqRiKbpZfRFgL0
wDA4PG4kId9Rg6tjnNaD9GBM/rhVmMtRpqByXQdKoAZQlxyguOLGuY38MFcbGxRyjPxy2ZfRTxHV
EHcWGpEBbWMaPBbBb/XQF/REt+pGM8GdyLpTdUtHdiJxLR5Hl0NAlAYwkyTG2lMHx2pnjSyO7Zdw
LPaDU4GjYnhJt0293S/UQFN7Bi6ei9uwlF8W0L8Xqynvyrlhk6vC3MesNPxZK/lneGr8Jr4fpHh3
roR+Pli3kWWY7gS+B+KoWdmqc8H94dVL8zfy62PwZN3Dp1GkMUihAI5GkSGnwxzejdaMNL0XkrH6
D0JmvX0s5ygKS3SwjYVJNSPIwVrwyT4xY8QKyayFGmiVR/1oHazuYZ1bp/In3N54xECDBS/9fUCj
GLV4gEs+aFJ85XJRlIF7jzuPN16v3LE6WGhqQRSICExMY62IWTDyqmkxLqIZiBxaCjq+Jntjakoa
1BYm2TLk7olBgRBA2F5e/DVN6KvlsnL2QhFD+rEbv+/ptVzVhdGHsOLmQLi6KgvhS7L2N7uaDVsg
PH88Q0iv16xxr0gc/sfOZtjRiLGlIcH3yCUfwiLIsZB1gjb7Mq6/8bjrG7phWJAQaAlhUY5GWYLh
4nvRx0GRpUdItdFHdzu0R0dGe7FPrUUpjHcmVC1MvbO+s145tVkIVJy4F77ZXIJb7JcRWYivhv4R
1ncoEeKO6oQQ+ryW3DgfeSsK+vhKZnLCf7jX2VO2LpNtSL+Fh/pU04JlcA5ftdudplUF5f5qJHwv
pFuBhG4RwQ6sl626q9GUhFm3XjkO1StkXfVMAfMHrENoY+rrJ+sd65d6MflS2rJms5hBv8yhetjw
XUsVf2zEoz60RO7V4sU6NVWVKzykfgkcYMuvG2pDpcUIEUcfWHX1cPbc4lGZCZHLIPe2bKEeXn2x
fBUg8JJ1FFY/ljgM2/TZHDyieIZYqSCSjqozQauuSJTphvhaB6E+0oPaZs6Oj7+GdoO7nmYAFAkE
zRMFoGQkaApZfy4Yu0lZp6jE7vN1aZ6gnlEfK1iLlNMJ5cUyHqxKJS5hsOMHCxpKnYUmoYLySLI2
BGeU8KUatoXtIz+CrY+Aavc/EjXSk4SEx0fw84rRYYyLExU+46otrsCs00EwXchP8d0C76Paiu8R
/5Cn57Jphat6V9YAAswlNdHAckfWRjG8RAoIolWlBB6QR8guhfgkgOAPWJabMIayna63DLoG79LA
BO9F10CWxhcTF9J4/HIeL8zz8K4E6YDtc2e40RwCBwoGIYBLyerlQrJfmLICo2UUOxRo2qoj4Kb9
Iucyu+1b7Mf5Jlhh4vcnpkeQBVHC0WTWmUNNzqAqCvuWz1x2nYyk+pBXdsRTe32J0f0uukOyVKVN
WXMGil7jS4LP8/E7qPNkZa4GqxD1n+iWiq2W6SmDyFdN83LNKfKB/RCh4qrW0KGhCKC37Pv4+DW2
y2yr4t3n5MbtvNo1uK4Z0BSC5r+uedxb7CedyTL8fwj/lb0nqfocbsybj9J8SrSYzX3GiDAa+3nB
RNwE5CCFvXS2kfaw6buOXMg+uoGRGL3xtMqqhAk2qJ1XceqO06RgzUORW7K5dNdKbwnHxHaZQKee
IL0IisAp0kgHGpwx3KcgQng6kyNKvK08vhgpqYjaldA8jqlOq73wwW/F6zP4PSbAXHBrjk8JArQT
JAGVc5vITigxoVesXQVJrNNkMbrfvqZWSzf03sO8voVfwjQhm5PM/6IuWJ63PHU5qGLldGxbwEWr
R08WnCiFnP3b1wmp75E0lQ/qgOzsFd66R5nvGXUCfvqiJ5Ral4TCnLHZBWARYkdqFa40afQG3AfI
s7zQUFVgG07ERtfEreNLl/kUxGFOrsRP1xKOfGaoO+o0ucAP10Z5gIHxKGLosWWWAdY4CGKPg673
EOhO9isELIVynk/nirFFiXbwzeiujFBGP+3i6euDd/Yt1KWZMrC5Dxc3IEr/AoRRsXaR32pQlmYT
7sXkp9rY8HPhA2urATdImuXoeD+CNFYvPbUuqRLIRqDTkpUvQdfY/mIBri6WpkqzQWWkVCWuKzlO
dAnKtXWTtjHQ9akSucUk5hCBvuMV/B8VNNwuvHh4YOIGRRViZuiTnkCceHJoO9vnBNl1Nj25twmM
pATTtvuI8iX0pQRgvVCQ0N46unpZ6ExtfXHhLLbh9LKQ52XsOUTthOEWkiHzj2D6DAGWOxu8JYZk
lN3V2qo/tQpGJOf6n0/SRXxoMPBuGkX53k9r/8uVuibnmqi6DTtHb6O3ewqqGLYVgNtDbDwexu3A
7HfrllCzJswM4bJU2MxkTuSqqTxxjPbxYr+xTVia2dMtSBBiSzySGEJdlBsEzApJC5ta1HzTm7/k
YRsOAFxiRTNqObVlfhpuJO7EvNJm4WwMOute4EwtBPLf9xk53eGlDk7iJX5BziBiITPwImyfMPH+
ZXp63g42KA0ZrHXxSBCSQHnZ1+E2cSNKFfqZOag7iW1vwXCklU+UrwkwK5mMT34VwwyY5fUymKx3
blOtifmIANj/SNigNhUhHqYI1bC0GXAocHdROmEPOEPsgMXHLJXSOS0PK9YeP3Pg+tBHksl9+rYJ
Y80o1TUPmBNzUYYaejquS8xgDGNObg/b3N0kxxiosn2Y8FVg6bD6n/gMXak9kbK5Hhk5HUcYZiMO
zr/wQwWVAdpjqXXEaPn4eFwZVu3B5LMuiAqrX341ar4zu/HIWns1/hmjHPyK1fx7m39wK8Jzo0Ry
2W9d2tyFu/LFAP1sv3bZm6c7wSfWSajP8K0R9ZKFY1d+ng6ItC4aeGyxgqUg9X/Ci7xEUtr1NHdj
2tVdAtifNX3GtOXXMoJaiAJ7hE6MBFnN3YuCfSXG55Ow0UW7ekKqS3vYs9Xoe/XlpN/KEK1113o+
TJgdOILy2J9+fZCvaNchMOpI30LyqMTUGPfJPwPUo8Qdx+3IMseTi/K4M2vMVGrqN1L6oMgJMy7Z
vn9Uehv8Mzby+tQjHXglNyM5XS4Ue6/fKXtFIQ59cobCALF3P2aQrFkOEcnt/EnUjs83STvnuF0n
QNJvS6xV2kgAzdVJVT+azqQsLO+aqTuzXfzay01og1ZHDQI9AJxllNllYBHB5mJczEXJjCgZoOVS
oFCE3VXzSgcGhqem0BP8Xqc2ks44xtYI6NeDfkNVoVExddyoUbLp6H9HTcjrtNaawTaPgnQprTrN
5HZWpeueEuPNq3sc42aju7gJikBvCWz27fxdROZimG2vkztwvjRZXPqGJz0wrGlwcTCJismRZK3k
CMpCwjs2ktO9ukqHGTqyu6/qQk3KipUHwhk6fWDKcx/AAcZoEo/2T00K2PuJLl4StCEB7VkASntH
TD7sTC7qE0Y0cmGP8HKd3cJ7Jz+9RwIYCu3w2hxePlRNqq74fFnU69Mp3bT5Ke1o+dkAnT5gxmpG
9LUAK3SrRNMrocx2Y0asYHJniqzkcUF0ymRaXQfct3y8nY+ydLV+eaO2kzgJ0bwDJyRkHbPU+2E1
IADyPkeJOFDqx9olDBUE0aDnXYNPmLgs/QKye/xawgKRDO1IfiKf4xXWc5lDifaPtVxnjknHKiWG
T+Uce3JitNSntC3VF1ZPh+3l7fevP2Iwe2tcFUQSeXyG0i04E/gjantbhJRYPaGaE1SWS3uzjiJq
ZmLauE+N/6KH9chDFnpHYDYb3x0nrpkkqXKQggo7eBXh5bSegsIPdQ4GDBPvc4zDIjvv+WIvyUib
Ra0VEJjRXkSj1LaDx16KWigLatxrfnQP8a4cvD8P7RuX0y2BuDVbcM/PF9BhjY2XxTHp//K+syoA
UMmrKNj0b22ArZu+Q1R7M7b7O8yg2+N2saHQMh8PzykltA8tO9xQznZz44F3kCGGE17l3hD3rSho
OiWDx+CTldUImNawmow3e3FKfTWDJRpHzDYmECqrSuHob2iYwZGPuA8H4FToLcdckiTE7x+u6hlj
tgnde3juS6HBjFd+q0qT31BB2pwKWY2i+jpqwu7AemnJtHrfQFqghnMIBiNau09UsTLwPXn50Ysc
rRP+S240Eyt0SJGU8CGCh1MD82REXVx979yCTiLyRp52QZATkKOPJLPx0Mt0dZeg2evgoj0qCsF8
tyYIkdTg3+Fty+bbjLCw/e91j9Y0H6r1UYuckP7GCMBgcpdv+KepBG47j1T1pJ19uch9LKvwnElx
wD5EYS9+CG9O2mu7dlWkI2rE2b9HIiBzvDtfic7HVAbr/kGhc+JjZ2XC+c1moevDwE2C0CE2thm4
e0pSXYkaIfs+XIIc/3dV/VBaQcnC8uumEzN0IMtVytRgp6q+CRO/Kt8bJ95tfOur1ueNDu/BObS9
LrtPTZ6CdaUGxFTsmuQR7mZ7rhi9wOUzpEb/Dlu89JOMl3zaxzsWhhvJdjwb5Q64kxBm09Qeg66+
K5l1v0MRKQmVvnP/VT/rNhd0kJtkdQlIv2HfBsHZ6eLDI/xLS7Kdib/dhbcJb/4F8CVZOV1o0agt
iNNshDhsbHDXwJQ4D0KqSkvsSdIZZMkSSYWVCSa/h2QGQldkISizxK+3WU8y/hz7kJ3aUQYtihUL
WsUXc7zW3fZitmegIyTIer4FF3oxwp2OsKfNYumu0FTfb6uhpbrWGW7R8H4LHas+WNncr3eLCqCt
h49EDvZqgKi41h9IpDvj+53DRoqV/JhQxzeVG3tn/dr2rIe/q5o5tm1zU/mPVz22QEksKqF9aHe3
SPweg1K2rbtxVvP/stRyatSFKaQ6LokIhn3WgJrS+D/DfuUAYYxYwd3IQkwKw2ViXy6tnlV/Ahxg
zBOBs6t0jc7ZB39MKPMkjHrGR611+YSDJe7SLpUkMgMNvXxTMgbJWaQG9+nDsry9IUqFqvRC2w7+
63Q4J+RK0zV12QEOd6RcvTXrHdWNIcAsqSdWM7x8cjSSQ260kStINhjsxbAUhTGTWV/TvFj72x0B
L4o2BiBJkJEXToeJEpGWR1Dghin6hefzi9jUZSNK6IhvOy5L2yq5S30uWOc2Fh78UBw18RVcITG8
4CF12PBS+Aj3nq+GZd4khOJ4jVyjl6WNNqQNdlbJfr/dvGqLAPcpPKdvJeUp6c0gblTI2NmhKSh0
gzjvpGPWDY+Qq+9c+uVRnhFtxZSAFrQJQFzRDzjK78Uf0Ix9fLgmHN2cHQTqRVASPzgqeW+h9IjO
Y7Ybqv3YbCLAys7o4+VP8D3wYgOTR+JEH2ceHt2PzzqbsEewRt2a3aY+Sq3F+wEMam98TNKOK15E
UZLS3SfPoIxuMTrp+cFg9ItrXIlWetcF5xvxl/Qk6QFl8oLGyzNo0S8tK43dJzY7umjxgWx2fzxz
hHfkcyfF5VJJizOpbX/NqlYbmWUq7f/h8yJ3cjl8q4SK/vQAaItIebaoeHPCOzoW7A5faoN9B5Uk
GRAPiGzFWthGUaLq8J2u25WC+EKO7q9oc3A+g/PMiwJxjBr+74CyOUooykwWN+x5zHmclTPu3m3Y
67Rvz/Ty8Loc79V++T13iILzLsnOp+VE3QfzjD0HLWoQBWzCf4KEQxDG/QEy+CU30QE4WeRzlDZQ
Vh5gOF7iYDqJ+e0QQvgXVg4sMzd8kMkhjJTdYgddzuRMqOUSwW+hAGmOqXdNlHUcR6CSVB1wAN5R
tsWptPWT0mDMBY1CKbGagHSAPcF1hwsd3Mhsgs94X1u/4rCtwgj0dRaUb2Hyc1hExZC8uoJS3ZPp
qBdaR6mBXW8RwhPiqV7vauOhzoFnGEP60889hawdHivhMHlBwORvIQXryBaK2fQVk1hlrDvW4KVU
PbyRysptcXpF/Srm7NZrrzL7SY4PqLpPsFcclIFGGRJ6JXCFVYmHZh6Lin1nGLZjwU+KaxfPidIo
iR1y+EaDSgaebIghdM55Ro9yq1MQWcHZ6/2TKvwmIfeFbcli/h3kSNvbzTMBQNHrm8Ungy2C8nlv
zlrS11bHE8Ve1Hc/iiLQ+OgpPnihcJNce2S8Y/5lZX4b3/0bdwJTsICjLPmYTvzbMKSE/ZlzbPli
ODtAKirzdzv/DoUzzZ3fD7qW6KCOqmSb/GBja1w4EGn6Z5INUizg/KbH9z2f8dCq2zEznCQ5D2zx
KMMDmjY8hJq222ySt1DYphqacUF+gKc98hma9gLatrzXL/bdwlYPBXFL18/+pUGHPDegGG4ijWJ3
AJYlk1L5yHUf0zPQsE8fwnR0FWo0gNkobj5YuwyX+dzogKS/k2/M+e+AV4ycm6KQgTOg6wVnVxc3
vjL27p1VW0OsdnC7pIiyjauOP7eEyksJwBYaKAjjYiizjLNURMeISwHu/4apC2f1bM0lh7WlJyH5
SsE2Qk+1Dwz4ZOwAix2FE6+XgWubUqjqPR1390EsF7FmBE5miUT/gs21ZgNhHsjncxkOaXx7Q5q3
GMYKSOm2b8Xfy9OVWUlfUWUMaxW2Mpyxu+mlRWP1IKsOGsHzw4BgbOMjeo/8bc+FKKx/A/Bgmjvt
slg6L3nqgOoew2TO7E8rWC7ex8IduMwp+mu3cbF88taV6U1ntS5WOQe8Pc/1BkNgSgp6YDUOr2ZW
iCLUM0P8NC0poMG3jHDqwAUo/PIBV6+Z2n8lntvZg6z4PQuYFNaIAntrQUNv4V0tapfc2zdyDsdw
jXRUfat+jgAGj4xZLWCVD+h1FBN1u7PAPMl4eOe+feNHkGoCyhFquqFiW9jLyGvOe1KhkWUqYEqv
coDbgtH/5RP16a14rMoDoha+KunO0ZH8EazFeR2xIj0Ko+E9F/zD6oqu9ste1ym5r6vGvzFtX6g5
ekimp5B1Rf5uXO5jVaY3FEZq/ZnRTQXxHlEbyd6ogDh9O2CRPZUQ+PGNj8aYFBcz8EIXHK2goC9u
cD73ohrVNCq5AEzYQuuxzcdAoeRgLWLKEYt6jLTEnE/dGXFq3o6Xj1WdZHnJsMIRUwS/29k+MDaI
7Mv/LVR8uRfzKPY4e21f8XTWIvd0S64FUJ5TTn/1Hkwe2pIoj70OPFjian9ASeSiydIfmojeTfab
h7wBMeimUxwY68lbRkHVOjk5qbx/AqPtB+hkrXLba2Tdx/3ILbWsKzKQbzoVVZXCQ5O8d33+xdqS
Rq5SiGUpWOx+Bhh38fhP72uuJZyeuhhzuPeS6mH64MjOzsXhqMBTndt8qmb18fqLKJKD71dPDYZk
ZVTxXqEWi6osln15JKtJrZyl6XEyRe25ekilzicB0lLYmKw33azOH3n+VCquLCiLh15RDf7f/yxv
QEc7GSneiGSATCO7u/VTudrstZQNRZQhIszMe+odk4Bo8KKvng0douQUms5PXqXTuOGvmF9y7/Vs
m85yEWr4KcwmbqmlohMpuovDyq8xPzHt02UIMbxx1eBaQkynEkRX9KfqMkHKeVC+mb0UHCzXP7Il
xqR5fO8ARf6YHNrbkZy0i8x3u27WmdIpRcAanSbJSPk8so5raqK2WDCVty4FP3ZG73wyePtcMnJK
sSrvMJX8hcCBRto3xyyrFYj4z6p1hdPJA7/suvhAlYfEEdQfThxIe4uV8x4r00SvK5T8gUZWupQS
fJv01cIc7OmehVzQ4RL//j/my6A93uJY8zCXjzXbk0EaZ/maTBkg+DuX4/uZDuB9YS4QK7BeWoeY
Bdb9AM1njyPMLFYtGaPeoIar0ohFIlkHEt1CqJ8m7wwSEuhaI0w69DQGGWmZdR+MJdQ+GA+gSDF1
LSCVLRHlfLkvq+iDX8VRV83ESC4W0N782cuuvhUeJDgtaWJf7bEL1gMMMQGHSGNRiG4A9DXqANTY
rzolgUPpwzOD6+oVOufF5TEu53eMAeZOzYa9xQ7LSECh4PbeWmQlMywvT3H/2hlkZ4ONvg+I4z/z
Tb6j4eupgfO550oZ5aN8TwItnn5bFp5g0hDRu2FjGs186aFx/dDJzE+68ryEmgxPJOGx2FEWuPnm
NSRsXTestSR0k7Vnd85LgnZHot3QCtWhMf3/wOcDgPP0j3z7Xe+KphXk39n3UV1piyCcjACTALI7
NwmZzvgSWB5RZ2Z1vJgMz5v8WjCgZFqcjsmhHgOwJPcwgJf7MJ5R/Rf+6wo6lqCzA2o2XCotsUxq
NvHEGreFmqVQ8JBmlsJedNy8ncj4Cm2Nn7UiEG+iiyGc2RdhM0/v5qvjjubzF9FBFC8+Rpq+8ATB
kYk8M5+q/psybWPo/NzWR/rxeTmJwvdwX6Kpy5MYDgoDR3gWweLvddW/mlI/Xk2P8Vabj8niUkvf
wOZ12a/6kv35Z5QZCPvBg19XrHDbE7uQjBjvduTYBvPH5nHII5lV5zCa11V/jaEEXkR2kuzQxxSK
yczoTJdrUkJOeKCsBCO1wG0eITQKbMtkjIbUFSu+dtmGxzsY6bojc9Ont9RK6M8OeI2f/SunCl5q
43cmif7WtNmzxpyzdFxmuDvuy22mgMAICBjp4XpZOoRSd68gCuOj/QTiLjPy0fBxQOZH3A2KUi0q
cOeFhuw9jHs81qJYMbBBTyy+Cang2elTshc7P0kM673OoJB+WGTAkmX9OeWmsDiGD6Boz9Xr02ZH
CWgvDhFe8hXiEt5btH6VM3KxOluQ5TzPtK8WATkOoDu7VxcuXjkTu0Gp8zcs8k7E9YWCoBCY4ET3
xTaMMCPYLHYq4uE13hIZgcXvGkf5lLkTjlbCi8YSO/hgwHMwHGI0GBgxM0lJOEe/KruQnVFUXZd7
L/lpUXdu7P7Q6uSaRmwr62qBjvSm//PRcjhdDnkvTn4RxC+lkMrE2tzPj9LNQTIadycJjdp7LV5w
bsnLSqlyqXO+a3juvzGyunLfW6irJsB7t3GQmYlBYHep+jV+rwz716ofFo1yX7UJeQO1TsaVbAfo
S+GNHqENBJ2osyIimf3sPmUj+kFIwq4XFAsgIEWNnhC9HclArCZy+lbqOo8irBalrNxDN6Jpiacc
hf4DpMEo50U5oGSwQJ19LCw8AxuclF1B4aMVys+Z1U/ET3+GMCYf57SnuzMwf31xNRR8bZZCrtOz
btU/SmcqftAxO48XHDR/K2e3Ju/6smdrJ7Z7XY0ZjLBdERc+FfXo2r6Aae1swKLl3Di7mo2QiP4N
1YKtkyE+rNDFCHdiTQk6uT9pIE3n6yetDYnQQ9+jwQDUlE+MfCJq3Ek+o8jj9uVkZJF0mK5IFMno
uGVE0OUpTV4pV/VmM13ZhV0th+XrY+xIgobxzZbZNChAgK02Zm+Q7Oh4Up8jWMZ2LAaxyAvhu6rE
Ayhf2LZZj++Vs9+XVkyr1m9glwM71vJemyaE3kOpJDJdrsUCnA2Uu05ZXURS1v+skrTWxy3s8R24
uhvvZbXwJq+HOlNq18eeNoA5T4MhfYLjzIiLJvXbdK7t2Xt4DY9grImGNo0MQ7bKhyO323KsFcW2
ITcs+yd2fyreu+URL13SMoQE+RzTJQD6x3fqVvPbLER6Va0+/MpVfa2Ozikree0XXmZPjg9a7vKt
LRmd27C+CGusxUgdJ12TAKV+ThKU/E72Wi09yZXzDz0Aa0GvSOwILQYqFdbowFeCb/MZoFUk9/qD
jKSZhdEJYew7VwYuX6lwlPOAaoyn7XdxTA80AuXZc6fybdGp5AasWLNfEQOPhxqTI72HSJui2xui
waNUm3eKzy+2kLp3OCtFlKd6fXxenaUbtz98dEJG0NLhoEc9f2E4kCn9KK5t07B1JFIoL587cyUu
AuEirQJdG57dg3UbNftvqc7Bsgj8CLVRrwTCi/bD1tMe1PhZ69E8oNOmeJ2DTit1L3lT5a1FBNsR
/BWbdaSQhSZbo4JEEj2Z5s5CEtO/5zYxH37rGZ2quZp61fMYUqiJ1Jhjp7i6ojbKUrqGqClqwq/l
Wa0QajB8wEm1sio0LrZUEdMvxqKEtJZJtkA3MYZ2FtxBSYxECI0DZkMWpvpH7d03cLGOkQlVWmAo
p3wQmT7YtsKpwDjSM8Oaam5rp/FLLJeGbrCGK1V25/neF7RextTA/agOpH0KDdAwOi8JpPcKzkO2
Gcdl9wCNzj2sJjOCBvfnz1S3jRrY0YFNi0wYzY+FqgWn+Szp/OQbGtp0oAwXX6wBykZ0ot+ucGA1
vybWp1l6gkFj2PnO1ON4cUL++jkp1njsLMgb8vw3A51nRtMuLOrOldS5a7voiEVlAnCQbEGNgW45
V1YeNICcK3rNntmJGLj+uVDCKaxP7fj/lnYF2wYkd7syxG3dyc7DcxAdc4V7uAo2ILhY6wp21XNZ
6VEimB/k9Vymux4F80InjOOurhWEMuFyY7/3hJCVqDjzjCvWK6npsBvCQnbDrxkB7ayQQnKcBNnT
NI/yTcQUM5oh8gnqBvZnS0USjbYY0FW5/eRxl9Gb1NakkFf2UU9zTj2g+K5VV87mk6B5RHKza092
IkzmhWwDde0IShhxv+TS59kwtse95BWOkBYR310V5xnGZ+rMsJejx7I5cEBLVhMaNmQv1cYwKcPL
o2C8KVpzK+0sB+ValUwkcE+Y7jWDz2FUfhIyvH/7pLKDtPJsy/VaE0/JnDAajYOsgpwWNp/s3ldj
qY99wsYKjXTubAbOAyaRWtxHCdxdtJkRy8iB/oB2K+4wAx7QwOXqqYI1hPYPoySvDEumcjUbr48F
0jN3H6lFtZW5bZLyDT7r/Vu1gm98lHXWFqrQ7gtAq2D1IGmmolpFmIEcPGzqd+Aj7eTtKJ3Ct571
hxAcQzgcIkMaVAiModMblFCb6ecGSQNQe9DBMt20DpQHNlbxvXaVT/33fW0+toH9a1j1VdgZTMmZ
uC/LNUeBjDrUZ5kLJFMvlee7555iVfD+mnJ6xTfyi9lXZbVxpiJLwPV/cbi6P0lrCq58Dw4EThx0
KN4BUg85VYIdO05Gtd3mZUkYQP+f/4i5HEk1O99V4dRfAskw03jSdQnKC8nmosxgdZ1zzXmNBcbi
teHLSDgR+QGfCVZOOsDwpuAp3JzbCc7RPs/8Dn41QxPHi3WIa+klfGSxXL2p9pSLd47hyT3ju3tb
g6avQKvcaQ26hqQkORL9y2ZU+ybiv9ypa/l+JC2K9HysrR0mj/e4iSU2j+y8svgZ7Its612Po1HX
2TMCNK91xZfdr41XSKtFnN2ThkTOAqY9wd7TAXQ7RJwLxpuxNUA779Y503jGaCqaIhwdeDsGTuh7
AHAZRh9GDs3NBedi5n5133+3Ry34apsGIPfJLOC8OnXT3Xb+UrpxcqqdT4i9LOrZzF5+lSriE98B
g+TRTm2AHCHIF6JZ5+HcHe6yVC/GfsQXSlg95NuZ6odjbQpMZPhP2jGZhXRhsKJifKhXKyfuA1rH
uTBabH3EgJ8yX59Ks5Xv5zDydvikm10Vl4tpcuTnlIVwyLysioFF1oczGym24J71G+2nfogHQWv0
4LExkpZng4pvHvfbn8lXMwFViiEOt6StEMqUjm6CaPJqUJ6L4mO3i0koKQMtByx4vlzSCqUwcGSe
LjX7jl9vGMMr/WFK6JP9io61pE8EMT/nkdlTXvOrBb35Fuk3JBewOluW2JH+sI/IXwZIcHFFc7jW
4MRWS7gdzPKL5kuR9qjTyFPkYDMYJrXL794MFqvMFMiKyu5GXgSA2Xi56HMm9jaar6U1arNCjVps
GKf9iy1l+07ena9rTsgjwGX5Ta2oXBf/ABKNIaHvOI9HOT50iHznx5n9jElgPkszLFUjFOs4f/rT
T/rMvvFT43+MBXvZHM53QVIIgEfP0z7Kyt0shSnRfOEN+j67/yFCN0szAv6S9RZFOdz099HGC4yG
hMSGmcqHr6NdQi2ROY//dHzWi36RRIOBFhvJAmCtj8APXTHS+h4dd0gA327QxtyFN7xNpfrnF/Ix
4VMss8yBf4vMqcOpknn0lgEBknw2MmAVBuyBqGLJocYCvgVOWKdRqMsNzlDsW01Y7DxnDQmk+ihv
hKTopex6QmUNCRyAjN0jQQFUwDihHR6ts2HozersvnNtA4iaTsTCFRLdLzhuOG+mSq9Oi5O1AKLT
gPZbrwK3vzW9cHpVtWshlr/RIiXMrG3bf7F7KVpUGPP8cDuH95riSKFuKNKg0eGYCZWqQH/VSHRI
f2zGn3mNqGZlpbmGSLmDzjj5TSnxqc5CryStP5MAJ5rHoQOfFi3ttQCMWAjjWcsXT3BoH/JrxhPs
Er7NZ6MLcKVQMmBiiuOP/j+lRK2gXY+G/WrpVQvLV9xQ7dL7NddevvnlNcMcSKGUqEcH/34FTakA
n71YkzJJvBDaVwQcI78yQXw3aKgq2IPEkCFGqkIR3QGhs/DCxKWvumX5ssdUqeSWIpyTxv0K5wMv
zWWN5f7quYtyScQOOL4sqAGkGuL57rc/I6XVg7uiXbRL1BcubbV7sitO7uDtCx+Jf8ZLqxXXKVTl
tUkh8Lr8xIxS1gHx4MYoXCNoVV2+kcqr2rlOcyYXkee8BeECPrSeR9/t6x0Q5sdCfAtjNDA7amiH
Z9wzka82lpMT2p07FrYpfPXYdJz2V1hnyqLnC6NeTpJt9QZEnsrsRuc/3pI7GrQGdwF4P9hiaLXF
Fuy5m5XgZHfBw7IM0vqL0z2mG3JBio6qzzgsWThGhshUkzLIs8u3K6t6vXD6kGkoNsA7Ft4UgZ6b
efscduOhrnogPlFOtVt49/Dj7BEI0+O9gCbV1julKY5AQAJgmJm0dmeZlmjl5f9CE58MBPtPM5+6
4WEV2tmPaX84pe4Rc7dbEAkz4ELfTTE1mQ9if3j1n5NxUMRL/m2KUNC2eYLRJwlLLsflTrq4fhM0
ND6JehJKzf8CZe25sJZaX1/XKsL6SPMecsRiKKVtWapu45lyfWpATpMDjm7zu6UdbhfUJmLKFYAo
DkBcfKzyDqk9bMVMBUzXwySAAw8Mwyk6VeOyQYoFbLrDZknsEQFakNLahAcfu459k2zwqTMyAEAV
Zn9K610Xwbuv7rGZZSmAWBk8kYQMMOVljPF7AXX+DRaNpvq+eRIv+LqPsVepQIGmsDu+J+jiXl37
cAUdz54BfRroGAbjfFVyKT3Jz8I0t2fNU00MPBeU9tPjySMkbq4W9E5AeyytWOK63yj70cxD8Di5
39qLGQxLwQqj4wH+RaHCagHd+zdhnYLYnDgyboAWFa/yigjMwFynqy8S4HzjFWTUa6TUIgqBnNwv
ZvvT7dUnzn9EMeTVWxre0RCmZ+5a0obMPF1alcBNJT/xdGNRFEdbWV6HsfxibJa0rp+Hb6UzJXLV
2edClmNoH8yWzA2oVynEFb2VqjW1gZmtlmuuwD16L1dUhcGfzrZcdO+I1PfZBc5BoZliQcxYEGUi
ctjqSJ1T6F6E9zsY2e+Mc7FS0TPKHHlTiriutA+krzDpqBszQYx+PjndVcMXKOcaa6SiONhykngl
ezL1UN3Wy9HBofNJ0oB95ATeI8cnmo8fcYUeaBnEqYWib4U2RsojsrVHmiyd/BXUTVA7EGPo80R+
sn6dG8TtpEX6lJoC/myRowiVZBWBpsW3qSeL5xFSQLIAr7BJGqvcJrVMT2DXpScHgLwnTFfCius4
V94po4htl92gvfA0z2nh07H2N29OOxlFXdHtdfHum1fYArtZALiOFhv3LbkL86jcegScrhSz6wwD
zjZJdWZO/w8YC12x/megDZWA/DO9JL/3qhMnjMyy5KankwejDThyP+m5copjPgJzsv/wR0Rz4qwr
5Pjg4qqYGI+P375rxqwPX9PbP24tmL2jzkFv+ZAaTufbN6P994C4eEx49agdVTXTBTHYHvhKeZIv
mWAenr2hGVgmF1Ed7zPzQmYzBGQ2JmTBKftbpWmVOSedQyDzs4HQgW+WvIPbqcpejtXOYblneltK
TRHn2iMb5IfRfftfHiEMNS5rS/3pNbwa2bNql9xZnyzzP95NOLE3RY7uDLt5Rz49GA7xVXXeYdc4
i9/zsrj/WVeZMkjEtXMu70sF6V/qqETSCHQmt6mS2MSONwT1gTXk0KkNd8z+dbcrbRukOe5OpEpW
7gMQGogNYbVpqxXiFisDtNyaBNJQHSHqBSjPL3fIuUO1crzZFnBdDemWF0koMeHjJxHzZxs9Hktj
OP4GEcejSfkmZt15MwYZEJpQzvmlvY+20ABeEcTBDYTEQrOrrQBmdN5oKdpwBl8dsrmbJoN1XEIY
SODBicXHsuN9fkb5Du0h7T0qEj3ryMSahULlcwFeqpSEaj14BEtNJMsIWkdluIiLeWORvhSyiyh3
vaeuM//izLcR9iJo19D5fYOoBaI9FM66YCYX1XtJxGaFUtxji8G/WDHn81Qp3SZQ+ny9rHne8GSK
eE8k1xG1yvLannwFdPLyl8ikduoHzU0nSrYWNznp6zloB2Pt9DGp/x54CS1Jpb3guxfkpbu7aQAk
y4UlMAccAkaculK6qN0FWRz+il+W0HLmP63dnW9ZxEYmlm5NCUBFGvO/zKCESkR3AmjeMgW7Twug
BKSPty+eCbj4ZrpW1DQCBxpYz5yxZ51UFxC+sW9DedlWkjdTUrMiodrGjzWvfiMkSmRoc+Ycazlg
9LRsa+vTLcjM9uaqtc3Ga//KWNhCHmm8ZCBgzJyAvLy0tfVEKplrfhEu8RY3Xm/haGKOjnpkw9yT
ggYESMHgNkMLIsUluvpoyKLVd388Lrmk7TxSImSSEdA30YtMGFzJ+HUJNfh2juSyXcRIUrIXTNLz
iIlC4yoWYKi89ZWl1RPLA2FPph7zIS+3UkkjoFVuyASJUJUQAenTVciDe+XEhxNAjiXeuXTqfv+c
6hkBxUSUgr9dMw9TNqT1lZYY5odnf692/ow/wVtZVqajGrg6+kZyLdYanFjWwKKEfK0pc9rIOYMN
ixWJsQoillANkHMax6xZ7iFIDm6HDbZTrYhh66GwDYJK7+Sp6SMalCES/kmgX7DMlOpsAAWGoFXW
hCqNuTWm2nIDfnJ4yz/HFL3K+aa+rW51DTM0d1y8WUsF9gxTUOXDaVjyYWDfJ8t9s4BXEVgLlWdz
6nnqbSeJOc2Ouh09C7FDr7i9QPKi3lzgVoZCPN64FWlt4xcHiTjeOqA9oIN+x7DasCdkl87nrnsE
HHJX8kn0W5Qj8YFljIlVCw03RNu6/FKH5/5vOovJEavcvClEw2O9L8T7HP7s0Eff22jHbbPha5/V
A+S0AgKZIlcgZK+EljMs2YCsdNkmf+Fx+HZWRh3QA0d3DzC4CCMZjvbkjhPKrEw7BgmOjl3ZAKbL
TyamRmuq8AHa8R1A5jAuWqJhq9N3Y9TWWD8XoVWPPiZpUuN1GzkSg2KVBxuyBUSzb1skLwi+Z3r/
u4ehhHusrGq6x1uMYDM59UvXuNXL2HDzgnFENQ8xf/oj8TP7AT5Q0Pm1KiYBxLVvz5GjoBU8ZqCs
UULNve1g6t65DroiHPT/qUjPLRrKUZfvweOpTKByHoo59mNifmVytJR09yJbpHa2XJoUu9uFHDks
3NihW6K4TGe+j3Hh2HIIcPwU7su4MTXvqzMJPS+DpDG7yG4/IlDVRv8NWmkmmtEd77IRs/Pbp6jR
cw6Pv/VraqIsk3k1c+EeVqBvu4wpD8zVjQVxvZGrDVVtkd4wxOGavO0Rk26GIM4P+XIoHFx0rRO9
aMCGiw8ej+vbkUmd/hVe3Dw5StGc5xar960JBKCzcbvWLYPoUxriOHjbxThBLkkobRQ7chYNN7zp
e1nhCq4Z2h+8Mhact+efXchcaYyoSYM8+61P06psAJeTdIMGMMZDe2CtJ1bpGCOSedowQH8d/tFL
jHeBr4bK2oGlC1+qoUOzQ+DilyggHw2x7u2Mfk3rvpeR65ZF0+XvocPiQpPOXH3Z6o85hMxYFjnt
h0NXmM1cVt2IKGymBiXuPf8ahpkoivmmrUPI37a4PcUk7HB8hA1XvNn25UYHrXxq8tzGRGYLNztP
eGMLc6FheXZQW3uGK5+160fHTkq8GLfNp1rCBkR3fip2mwaKXXecx175Oo7z0+J9Jkj5SD0WS9N2
aJbDkSlCxN4GoUn5KqR1/0dM8xv2QqjrKuzO2b3v1LdeejUZ/VH4mA3LmvEBQS4RrzCjpjYtZH35
XRqcNcbF2iHUiAQNH75pi32yGrtlmatCLLYwgmrK1Pg30PlEZAtpNi7uK2urn4RC26eZ9pKHlDhM
ZF4mNHqr3Dp+iv5kg8th0kTUpsnv7+bMBk+16ptDWWAJegKbu8fewfE7037FTI6MydN2qRlQW/sG
TDVxAqcsXqGPcsfNMAi4j5VMNqVHlZTE/vVj9t8VckRYBZgIsEJdcLgougizhHwy0Kbv0o3uLLq5
X9U9yZ74fVgMaMCfR3aWSABvq2kc2YVY9KaV9vjohhyWp5DStpXf68NxEqHkQTOy6ISsqnqxvbLV
h6B/98WYd17gIA2n7sSbAlYhq5W5XS7xyeHhJqcXoQM3SLJHloYbO8O7hIdCejWJKDEcuzwcjWI7
0asYK4d+vHW8WAc91SLQ2n0miQejbeO7WgBqonvCuQMk/lvNj4Gkh1b8AU1Z3T6i9NlVE2yZ1FTq
GVEqi+CRabYUsl623YeYZZoWn0GCYhbn/HQOfIg9ia71jsl8yrGELMMzJGdCJA33s1LVkauQXfA6
n5YD0LvzdDJ05OCV3BaOpebx0DrQ8mI8BtVnhSudN9g5WiF1eL5Tkymqqs8zfMzNgLklSnjci5Em
aFj1vk0xe9vd0IEASy1IyeA5uNKqTHULUzL3f6Cx1HhITnDekY65jwO1NTptLJJRfoaXy0fEEk41
9EsdfjhZSywXQAbRq7NGA5aJVPCbI06YRaTpLfDxi4YpywD05QwouePnd8DDtWe4F9yPyQVGxYxI
IMxE+ovXeV5UBPcnBL4p8tfl5OzUrWc0gs37zgXpOvy407yewmhpP8adJhO4qLA7EaGoyn52bB9a
gDk1+HVkouJcDXMcVb9uROoGB0NAGbr6yFMFf90Or2mbEmgbBbiEd1wJ4xwU4TvcV81ESPD21x0w
b1NS/OSpKIYiZd5flkAfb/Aog+Pcny6OdpypEIGRNEs8okhFK+iZxAEXQ6F7TE/3ocDvlpi3M1bY
KBCZ8Nyp/nqYQ1qyxtH/KpgS39zSzVgI1C1VZPxvj24J7OGTWfmj2jEWA6L1AdSf5LYzKlsrQSho
TrIJdU8e+nRkujnVW5CpJYCrNF9C5i6QBFlsivwf4l8dM8/bxE0a1dUVQo9QDk2k6aLcandY18o3
f4SOq4hJPcN75fZe/RLKoz/XOO81HSGJYYfPIQMwj9jsYhSbg4hWL3w3JjQYzVnikxsPX1aCCHfV
oVSqPiWd+Q8Z6bap0ab30WOaMG9oqM4GyUgVUv40GIgeZUHYGyvoXIxts4qIOjGVonm7FzYwuC0E
9O53DLNH+A4EZ+tXp5+gm0b+/b9tH3SLj5eDMrHvbnR/5jxMuosrutTh77JehiE3nvZehMRsZTg6
2N/9CR1RNOgQ0/QgoAUp9CeQZd4NuequGYMLEMR+OTRxNi2UDhnIxpaSvJ0Ih1wwjdcL0s/Ris8y
5NCc71CfarrhMssHaWP4eOR2pjqzEFIXB579F40wObUd8RfLGdKW2ULn1JNv5j6konmS5GyZsq/K
5UDNTs9nNQ8+M/aWzUKnyqxOlFfWB1KJsQ48t9fRpycg+oZd8sDirw8AoI8TCfuvwqQBLWL1ouKw
gt2/0byb2oaPaGm6sysrefwKwpfP6HEMA+YcK6OE+3R8UPndbAtNAr/Yi2FuVeLFt87RKf5GGHtq
1iIkBXkbAre2KgbiKc11sZAAza7/OdLDqRn+CVkEipBwedVj4iiTDZDp7mLcM41a0jZy7kuHYep3
fonjGKSv1+3jELN5HwZu+FwoFngKnLVLHVb0K5qr4YE6r7w6Sz+mpy/ELoNvmRSAQFudJ/jvL+fO
JiSQI2STxkK9ZrFD3CeQOFwMWTnQaxxt881OQ+Ep1Iq2WurrjcWfcyF0kPKT7IXPx+jDRXvSGz5a
GJenjNRH4SQlwfz47CY2nQ0njTX7F6fPqVv9jtqlcz/1T4lURR8pZfw5bu3Dd7zDsxBkmuFvrGfe
0lJLNPyBLpmb78MByrAI01JQA5iHNBBcAGL/sjEU5POzYE0QMW68Re9y0IwSHeZ0ZduSQiYSTwUS
L0DmhgG6U12oT86L4pfrzFYcyR5GfPNihP1ZPKWR3SEEvSs9Olipqx5dlbbKQQ/34Ze3CeOPgKGl
K0wFBPGUICqBCDk3bR6wiR1FYCxLleoVJTk72T5buzcaLASvfKiNDfWnOFZzCgy1rhOAny3vy2VK
9WOaQGzJFzFD8FW/LBlDRQPY22kJe18niipxCVK4kMYK34s+B3p2tO27YqgZkO95BcrNigvvoCo5
3qI1vPN9Nhl7u/SeC4OKc+MtdBuf4tbEfH9yx6kUa6YaCEAHTApRY8diukdNT8NRNg5iX0rqa206
fZd9/2dnZzgO+aTGrJCfKs6eBt2zc7jKeoiRge/Z7AguHSSQVwaedqy97hur2v2DyhSDHD2Me5oO
sISgoF3kYr1mdA/YygRtxS54KFXJHZF6cdqTnsT6YLJILvzVDO0HMq/5DDCrOnyIDuDi2P2dyFUU
mxJZwg45LRP+mgEt+wTh8/cDMyxmhyAq+52NXhuU2QXmTl6+6b68YRRd9yfKpRvBe5fuDkwkQdl/
ZZjx1dGp0Xx3cSsDoZw0k+vbGZ0k+G1uCPsA+l8ZEFpHgDH688UEcEgePKz/ToXWPp40koe7Hcqj
hw+drH0hlS/tGFyk5JH21X4AuNnaJ9bU3OAWWFeL6FHOxK9+1LTDnRkp/ctw3yxXQbrLwFju8N9y
kf/2f/2Q+WmR/niMMFFQGamvJBOoES54Zn6buHaxzl5V6LU7hYIkpESoUITizY/kIqNRKoGX3Bwj
t/1BnNiBAMtomoHx8uXJ5yMZmUhxP8tk/tN9hxi+MMY7TrJExsgekrk24AMAi7QIlQlP7dPUUxIj
QrPlwlthopmH1jld7QBrbpbxtcwgLHiAmFRl1mdCV3W5eaCsV3WAQYWFFlg5FA4S0Nxrd9kRY9zg
80CIUUczNWbGyMwHkOoZwkB6ieMwmOGrXjCQf/zGzIoG5BQ+vvgQWhRXtKmxyli+MfC74XEPeqYZ
xnSO6zGUznvrZNPrpi836VIIgl8bGWXtHyzi5g2iz06arfYJ72C+8wp9XCCFXWcP0ZKfu6LXp73b
aJD17QiWQXs/fMn7mK8pyvKG78GbgVNZToDqgXOa770jSNMYIw8fZBKz5crWSkGfek7+3AxePOdK
XR+ZIhTGpthJojoy9JcnR+K0Y9ygWPR2/dRX3ZynDKDvItmQ+AO3H8657YMZhA9w5nLGZIcSpxtV
fGSylCzSik3aC2VuzxGZWZv9aKZlEYS7ErRSl0YK6CYnb2GdRPdBGVYefFiT1IzVQ6AobxWX0xoY
Bp9wdAEp5bjnC1bDrD8daRO5niKeNVjks941TGMFmiOgjlQ30HFBfRtNZ2Km6OU30dD3cieGyuK/
cvijsPIrTmBM8yhkEKdbgOPl66tf4qax0eGWrANfegbqVDJzCDgFGe/vAJZTyoguKZUIptdGrgBI
6wENCnj3ouF0VOjl/zXN95N0R/taqdSczOXWstUJBHS7wv08dmXbHWk8iEp5CuBI2x2BbGBgoJ8t
lEChjfe6RbCswkvEO0D4CChyxk4VZoYr4dFPSD9tiUFV+YWefbLenp3S7KdrkM8exsa84g0NqxGA
AwoQ1oTel9Iuz+oteqBjKNdVY9PDfFAzts5FJs9HZgeuOKex6JeNno/7qI1zAOzdAXINvhxFxSQy
QoEtoCnzy7j6voJrLNE6zGYi0yDFz/t/yiUMo0DhxAZiKKIoAPpPEuEh4iTMPrxJmsP3kYiWMV43
RDL0ErxaWUFL+qDynFWoSxl3iXfBv0NQd1d0XAwKllXO8n2hWDZDRAddpObdPwJuZa2D8hHXG2f8
ZQ6NYsO5ZDNRNNvmyEmgPDQ4Zt1T5qTmtorFeG0aSCCoz7/f6gnwLj5zuVAA8piKVmIns+kHe4RA
L23+seYgs5x+qYV92SkggEtaxR/Ua4/aMi0XQl6Le6A0jBu1lSKlSHM35D2mbkMsDn9L7TGLFfgQ
8HS59YSDS74KorRXuffdyN9at5/7471RBg0+LPqBSy3IqDOsvAuELFWgGyRLH3Ytkmnm0gz+P516
IZVXdg3sX+AFQgKqphyO8ltoFkevdOry/Estqij7nzcbFcE/FxgZ2chCT3V6ySbd7rLF6DLd1EfZ
9Pi3ujc38X/pqDVOmkqWp//6FjF6Pf91uyxdUsGwlXO7raX/vdU5RvlYaxkvbeiNrwDKl32mKYMz
ycq2c93gTZdnTcLiBjc/ZQR41pdjxYtayyvfQJxmnoARmJVPT9g5kLiuP6xdFYTiswVfNLkGgG0S
fA0SYVQTOTix41gNavQQweW2xjqLMxqpxfg4wAqXCDEoPto5c5lPwzFAVn4yN3wsTdingAAUGDg0
3s4DEdv0VMcwRkOixLwLjC5GcLpbFhTp7F+TkCWxsmTOsaMCLRus7phbPolamRoyU8+vGUom6o6Z
dpqdk8HEFW5IvzpaNeq2FCJz2o6EeXwu1pyPj8+9S1Z6WSD0kxxGlY7PWLNzJMSxkyhc3Ap3UWc4
E2PPgs8EdVDbywS/LEFmvqOBSl4dOUFXGh2IP7+Ep5KFRPAYWHgTiWUdeW2BqEHVFfM48gYxHD56
B0LjyNlGeJy8f1owsn/KXBuuAUt4SY8DVA15VV3+FEU0KDRfJS1wxVSVhuXfDEDLS3umdV2D64DW
jMRJeuP7puW3nDcMB6o2Ft/4jQxaanmgASbC+yIUCOTRYf5LiMktle+7SOB7rOH/74ED1+l+7Nfn
vweHa8735iv6pyZWkFTjdVwf9nEp2vp4OC6TVcUrntaiOeVQm88pQc2j7GJb8DicZiSdKtdEpAkC
H8sMEVbpVx82ir67hDQwqyVXFbGQFVOer3OnxEBPMlAS7B4e7WcCNTgToVBQbCcyr4aZrTUDzG49
cTaqKByxrrqCFeDDPyUGKGCroo0t7UxF5C8/oj9l1np0vcTgM6aMfRduc4TVukT8FzrSrnHf5Ums
FxMnFfsvVcVAHkZdvaCdcwTWt6z4ENdNYB09LHGj2r7FNo9i63oXjPAJmsSwzGoxmM6m/grAEEQt
0To0+5CGi4+iaZT+mhF4ZcAQOqfJgjz1/fDw+UZ12jXEdUN8Jj9ea2dfGZgE2ecGJAky2ILysV9w
4iHeLaGOnRDj76RUHTSc49ejZ44PoVFrC2oDtJ4fDnB1cxk6vEgPwYU+BvGPmV3wmBkdHoKD91gj
y1F+kOaakPWhPqEgNof4QYvaExuRZIf7uRsR8k048vI4wVxYgvFoNOuwk2PPn/w+8xPKwfe2ZV8V
Qpo0VK4ldctf8kHK3p287AV3ECw1DalWVhus5p3LbZzrFTH0h5R7KW4uRDQcWO3epzNoV2M4/MQQ
n8DSGpD+fma8Ejkdqb1w225V5QrwJ2ImLmKvZ0TbJDPUE2gbFE887ksM71ewKhjO9snbSgA3qWiz
eXyALMURT26rZYSbgN5gcWIdFFfGu0eZ2iFhD05yxrgE/Fx6Q3e952mT22rlCl4E/RlCSuZojSDk
EO+Q9bJhkusmhGbDKsJTgUGm4jXfnLbRk5jfy2WAWvfY+UbgN+A/8IOcz09tO/zyvtMcx/mffDYM
gCJvtHMMkL2MH4CX9Q66EBEtFl0+9Ajsn7thaVHxX70Op3FVONCTN9Dn9NtI7gsWFjoPu0gK3SsG
otIpaYHJuwWo5QbrPAkhL2bcYJ7pUbecKBf/IYZNlmjsezL+SiYxSw9Q3jqdU/GIdRDNGxI/Vet/
guMFLKye7Xvgg4qf0r9jHv/HoX4Im72IP1R/GVaTyXaT5GgGetUS7s8C9qULZPjQiR2uP0sLIHW4
v5ya4K1wYxLZPHhqXL6F/RiuayUHFdEjgFRECbtoHxZfgEElEfTVNgyrkJgcRT3+e/8fKQYsOEUd
0Gaqa/OuOFfHhIOSCuCutnzEUE8rhA/H4/YWDKLGUD1DLcNvlm48+CVNPcrpsGyEz5GJ2h6mTBK6
3wv9iBDmH9ckIycuUDRIAUgvx0HvuJVPV/nDrSFaqHak4xqFYHj8Kqz9MXYeJ4KAEYR6qKa21BRp
2jpO0mhOGQm4LzF3w0TbCsGNCdeI35Ami/xXNQTHJ4gJlvlS39uSFPbnab/yv/doI4tzXJmk3rU6
4gcNaF55y/gCodxx2Lr1FaZ1Romwno0zKJFEyijtFMGOrRCTgBwEfRe30pt1yTXPsZVAsK7hRiJB
44VeR7qTInZzt0Q4YSRTHpKbC6Lsw2XdqoR0FpqhBERZUfxLW/5bCO5oDUcY5cBevjuLkep9p8jZ
heh23/IAIJJMZOwI9cxDtlOewSJRhqRPKNJsktDe0enXNglLybAS3JKCFndy3KIuK1J3RCcBz2ON
IRqovzwn6DTLxfgm4GXiRlGEVVDMWjR1Hc7JFIVApvvYwLgPitugWi7Bo3GuGdkSHaiHN6dVfYdx
aAR75FwtcN3rUKrRjBhm3PzSPQtUQoI+kPHb+AfrK0v9dZnERO7gDGfcK3Qu+WfAHAkMB/vSoCn2
1OlCNanrdfyYveFusVS9Cf+DZZia30mxwUdn15cmQroDbh8hq8v66gVdWtuesgi0EAQqt1Ngsfue
/LacU6ZmRaCRX0ueYg4W+zJ9MXSV15tJnzs3jvcGLAG72c4Z2mrQ9dY6ebi5EARylOYTVlnQD2bB
K0A+m1UeJsCCNMyujlYQmsQV8YJKJEvCfK+B8vnAM4jUUaz7Xvy8OY7sEWhNROnoOw1fAJ8SrIaV
Lnvi6buIQakBp7yGSmdPS3jPTBlqmc7EuCLFcA0uXoM21PejpnEfS+KptdQ6SazeCiOO9s9KhSZY
HAlqlvMJQpyCMdq95QatHg6e4Qu8V0tdILBbZ2rt+2g8qVqyUlMk3kHZ1fK0xVTiQTrb88IkAmVj
ATeD3J2cnh0+6G3EbnSnWvShms54LWjCx8kvr5Uo66YWDGRWjw/OdQVZN+M3Bn8xh2vyp1jmb0Q4
JVpTmLUx+l35trU4yrsTpdJ9UbMG9qnL0CC0eODZHqm5ufxxFiNC2/DMnqzdhJCcyf5HFqaU2VVm
redQSSdOnlhfw7vMbuTpVHIZ/qvhEBJyRj8zO34PamM/c04ZasNVoDUCzN3USx4JVHDfzpno4bMo
aaYHSVs1KmvN3QBHATn/0mXHkft99JBtRqD6D5iZWqYtXzMGDumsrOFOUZpBPbeUVY/rtv0rO6v+
nTvrJ9puvQJSpWqRwGgJeRdQdmsuU9d4VY9s+xAl8Xeq/q+odalTCHXJMo1Tu2TZUXDm26IZZBzb
Djhn7RDeXdP7p+m2BmvBhBZUwv0JdJBBTdzFpa5MC5zW2dUxv+VBKsdIEC8B709THpPUqpxJU/zQ
A4ewskHrRIBpI2AkMrIM4ClTLWcuT1AWKD/QJmYicIy9GSTfegci4LndPK//Jcj0OfJsH1Z6xd29
l2nhe3zXsmbAATKRkyK1JuYvAhxu8/J98uMcmAWBY12eu72ce9O/mRPUkWfmW836WqecE2Hs5edQ
v6E5Aw8Z1/dkOui7J6CoIpHUgAKHLkmSXxg5MonxTTUl8D2pgL+aV/5hRJhT078cwl57Z8AUsMbY
c60JHMCJFa31iR2gXd87ni/G9xDogatjJ7pKsTJfoG5spFQVgsWhDgzIXgunnCbVu0/65QtkJXiI
wJNB1td4dr6KfOgQhhRVKcg4wqUXeyRI+E7VLSc8VlFYtFCZkPGo0MGjXd67gn4ZTddG2UlNmIOj
n9dbTjD131zk/jgPEv3oKL0Ur3oVxV4xm7iCAQFEWVoqEOdc2+HZ5FyET6pqX40dM460N0Npi+YD
E2cGkD0vIBE8WzkpyER95uqtPbkVQebDKzNlieIi/qC86cwwhYbfOn3Xg0j4yPWu6eppihuHLKa/
4ujSSSs6G/nsFdjhW8iuteyb59/Qu9seMet913EKVJTlBPXhl5UJuV7Y3hUfDcrGhOdzDAy/jxBK
/QQL8WYANqjQyRi7D0k/tVAGDf8vzeQHjXdwInX9E6/9IrSuNONLvdo9WqF31CS/uUxef6zqzvnF
kj6D2w59wg/dpo9r2lO69juIPzaPODD06QHbMg212icZH4PxmMfHNY3QNxPpGb2aXwdPrKEER/8Q
1MB4yq1yNR5m0GqH5Jp0WCN240ckr0wcIdCkkMHBNaBVoXQAgyGeOYt5eKdRvHcZSc5ybKZdH2o1
zn98f8Rsf5HA/xNPEQc4wLzNhqBObXbigeeZIzUbDkK0Y8Zq/k4haO82fpQg+s0gTjbK3oFWZ3oE
hGexx+iHIt+qjRU68zwcl4iupT7saiaI6R3NVlgGwn00nXfpp+cI9N/kHqJZ4Ry/Ep4vkkLMSnxo
7nl0CDUmEBHMwTv0+9zE3bPhPD/slkHSXcSPgO2yaVFtl1VfNFBfjgI+2Q5d1uATv6fdbeBSJ0xw
1GnG/N8n2F5uSsiAgrEW4TBh0EGkuY7/JHTdJjxpZd/ywtU1v9ZNErJEBsP+cllp3Ledib7E6OQf
q2qtNLqJC1Mm1MB/R7SmOElpOCDbnrZ9IUkvVmgcO7HMbJob/bEursCzkO2LK6elb+S7FyZgi/k0
v+Rk+GR4rAfzBvlguix3PvORXlNqhc6oeapj0bveixkS3GXS40utdiBZ2YnZ3rI8ZxRCNNOx1Jsw
5pkR4A5/pTK4ob44Cx1DUfzw3bM1cSc9PP1wInFPdB1YlzmHUxUtjSOp1vt3543BeOzqKI0yHuZt
rtgjGHOnpWRThGT8JYDzF1ZSlb+q4qF8EdjsO1H1Mf0I00Xb4/21aEfrifY9FtbB/CJx+uEDXekr
+rMqecClBanctJwCXgDyV8dnZ7xSEZfl6zJojW8W/amjCUx5BwlUdncdxdX7ypNaayF0ceCXn7ge
Fs/SDjtsAERFPri/wnemcvnI1sYGlpErnHDKyBsCL6fHwheb0SqoFsl4o+rijLGmdCdwnm38tife
g6llGBt87c1LNOAqX9Uo6/hFr0A/19mf9M0YG0eAphtKpVniRqW/j51JsIuchxh3lY38o9cyNT6f
ezJ+bzoUGUpUjueQhhC3PI5UxPcj7NS63GEnHSZGnxB3N75PnvGszev/28nT7Rlj1qQ2fDnUQnpH
xJRuPxfKp5eCcUntgTSJpF+n2w+6rU9smrBhsUjq/vkQaIzWmNLkqfIWLBHHTy+RHBU/tG+i8wtZ
OB/Y+0JVXeFD+oPaapQmIFKOL/u6gP8hA+4Rzu8rclviw2jkn7TPNayFdrwWoDgzj06MhUIpGjdD
0osQpPUkoYYcB8s431vtO3dxSNwrXtek8raAelXf12bQwpOegxAPSlV8WuIzvmlSuZIIXTu4ixwW
q+dEeqTgCAbq/XABm6uu8Zxl/jQglAdOFPJoFWqwc7+ikqjsDKABrZ4tkzHwYVUkyvo0obiFP27x
0hXyCxgF7KscpmeerrawPpuidWVNh9TxYaZx6X3ZfxYJtjWIzn1EfyOtgGcVD6HQSVWqFBgP5t5/
xsN6pesq3Wh+fX5xd2yqCUHytmELh5xT6XPzAa4cR816MK7wGPtM+Dz99sk803csS4b9M1WlWfaR
gVVs85L4OGnthcA3hYCwz0VEZv44iqwM0YyVIDLJZh7spD8zB7/ew/M6qXhmW1IO/HqB+9dRAb5+
IR3ul23rRvGJOodsjsmJf9cisEOkgNwEpaJadiwuWxwNIcKBO9gfDODKNrb2qr0nCVJJJnlBheTw
E71ZIJaq2S9bSX0CwZ/ufAKPqmKa+m4NtuCJVOyZcKcGM17lTiEfGh8Xw9NQVUeoxqAUb09IRStj
57+kssbzqOIgmYVKs7u0eIZTGTzls+4D2bntxdtf60/RL6RLF6UvFPQ9qNrc+7jlvxeOezjBLUcV
083/VQH9rnkQdTUc3h9Frr2ucp3GgSZUJpFyPUjbE60XRNZymQjfWuPGdf/tGXSCzGml2XtTR5RP
7MMt6mRmCo/bSAtMHHEfDynfyDU3W/7JOdz1wiDjcKblM4RkJinO5t6pSdObT5u4RYHlqzq2Q2W+
xmc3/cK9ZY9EO/1i+sQAWbi500RRqsVFL8hRNsnJZlHOJXsrkbpX9HDfK0Yexo9KO1VcAZnHk0SY
O6r5ZLQp1WJRnhAmgfdw2JdKeR4eSILFNS6ZqRZX1HYjxr/+f2mkz0PqF8ro8Psv3NO7niK5M01t
O/3c6Mk2IJSDDFQsbDiL5dLcY91R9y/cYnQU1f3O8rNpw4cVtoupk4Vwe26NqIlBcuIXMHevyWC4
/x/qx1v34vXCvvpnaApWmNkiarzejPrsLrqfGfINd8TRW9hWEthhui91QCviwZdgI6oU+6lY2EZX
P/hZ8K6xUU99kGz8z3Rtoyp7789j0Vq4eZEepI2ZuhGeWtzQp7TeAesjnwpnoaRCNWolbeUCvQmr
QuQEkLNoagc5KTU0PHQexH+rDzd8UxhyDobpo2FBw0qZjspowpOPAUKDP/EhiFzaW6SYumafTJqA
aJcrTZhxqtz5XzjWMiPslposiUfe8AVIPTQ6+USkiI1cA81KHKA8N4LFaBLlj7LVLE+5e9NBGK8x
4xUwuLbhYeEG2tytK7vt2/Lxf2LxRwVo11GHugkETgnOWNNqxax1UbxWXNRt3GAK3QlQtWsSB6ro
oFxKceb6XFiufAztXTAJVaxPknwCYxnLYsvdhXYgCv70w+eW6RSlddRDIlO/M/O3+jte2KzKzcJY
fZY6vlfmyFnZCoJ7mZizTnCENE4wIHyWFLqNdxrm/ROqEvIxk1lqELwUnIqXWAYL5vV7dprNL5r4
QvIYBzUaq3Us+R3vgXo94htdfY/KLQbbFs1A1X81j2vO3Bks4Pc16huLxjIIomikGx6LNBhRa4BI
xIF0JR9kw5VHOxx+FjDRPj5sBs4edME3TV8Au3FTgf3xT4mZRJj+JuCMpe1M2CUGaQmckpsmR5lv
hqFxmfNUIn0Yy/KBTMlSGy5KorbF3l9OU6OezlB+VpULTdGkYfPtEEQQcT6t7XJpO+evKW6ZJFGY
t9Wjf0q1jNKxTPe8AfVyoZFV1FfsVIAGDJ9dWXL+pslWdIeIt60eUykLHfal/QFubtuQlVt/ERFh
GWA7dqUY4tmr5+5nHGEWRDyt74YlVdZHIj9aFlyvscb3WlsPexvJIqO/uRTmqcnDGDU64AGqMknw
sN5gmFe6j+pRXQYfoxFIgM3JL3snnic5ZOVwFwsEsRYC02ghsrZTxSCGYHgvOwsImIlo91GY3wp0
N/QDjN25sMShmFQgwReTWkwvqDVLTj0+SUr8qbY/5l2SAiyDIWW6KDtg1qiAVBNb7RUu6dSAODIi
PB4wQB6v+em6C9zZ0ICxO/kY0ZNnH64vqHqYRTclHlJnFls53hqzuARXmPGnemibUA7cJ0jBdns1
dZ08G5o6jAd28eASoT6HJokvEQdqdWgoH5jkS5m6tcRzrbCgy55gmS5p3IFmlTQdZt+5PCd8WeMD
okoiXhpC1yOEkCZOPLX3SO6KA2p+xe+ieM2/Pc45PlkiGBdg1Gc1KG2MRkCynjGcbCe72lIjrDmX
tVmc+vkOwqjq3huherPFUh2l1fae5HDgd3Vatcw6msC1q7tVcoMrDO4Xo7q23mJdw1LH+wOX6ewD
ger4kQXDCR1tqSL/zgDRjZXxm2xLeRTvP9OTCP0DSZlQpVOi7SD+A5Gk16IWKnI3m1P+4WM1+GG7
yedlitFxGzbToF5pYaYwzGVpKjaxRCqcqJMJFEfSjYXuL9UTaaAi57n+ttL0HPJQzv3vZ2j9uchD
0bmifdDqT784eFURZ6jO2asFgO3e8mc/7jSMTLajpiSxtg1JMaPKCnjDoziWk4UPHWuBYDvgongY
p0GU3dY3i0aa33VBsmYuk19mWCcODHtxS1MusnLyANGfcnju9in4kOqc9WQK6HUEKgEdmEqFShzy
hKP66+WK5R65b4ytj4zzKiajN9vH3vy2WHoKIlPXqzPsCuEAyPa0pH36/VIfsw2JNU5rWjGDVICD
ElnRbyNGY80OAktDmCmiOB/ARO4OKbZAyOoc/l3YnQx/jkflqUPc2krrEOJHYXoIDP7/E5yXRzqz
Ahm8cimhg/e0YG3xv1tQ2tGjsROMFIzzBoZ9ce0ey243RyDvo6RQlmFadba5rC8QK7chBzs0r1FT
dySZc9vOSsq7Bauzkoc1+JJ+pxykMFD0acWTq9d8LPZv1IaEMezm0XkmXchpjmUijd6RFvGYFdjd
60vkwkCfdDmEbYOQrqZQTncmaVSrDg+xsv7h1AI6cXpJDfk/SgjT/V7yv7OW9e0wlSM9nJWbGclm
vpvV45q1dR416SBZEO9staKwX1w5TcFhO+iEoi55VUrw7APlOv1L7bUlDre1ibIVL/aJC5uIShPG
ZinzbRLBHpHn2qdRXJAXKfg0hWVEVFSF7DU0vvFtMrG8jx7xOIfCRutTXPvnR3prTyg9Rw96A70Z
I0346rrYRf//SrK7wGLMP89gjJ0pJwrtxMLDLmtGwMAUQyucPVi9a/k57GNOEQmIK54paa+FxVsB
Q1JuVO6dzT+cFHJ4AP60V3P7+LDAw1cCL5oJbRumQClRN4U7zVS846G/t2S0c3nQPJIczHldxftY
JRUWAyH/4wtw9sj/8WQ5xBkI9vbuJCulc9plKufGSTvZNK8dnmkUEBm+EjgTat8cBPhu5c6IJsXQ
DPXVWMNGw7sGvvckLz85TOVRjUw1+OZXNeOYDelnpCSPBrp9c9q0iPyq7QFhjwEt/v6bYRABgx9X
OHQ31jz1m6ATANnDPMNrI1m454NhsBO8yrw4AYvYV0cAZ7uX5WUtXi+q8vWv+H+X5ip2H0j/dA0z
k2Q4w6LfoPOTrJ8j6wm6WVQ1VRs4zIXQQo8c67fC4CUQN86mcmd/DpwlBjgpOLHKSmKoZoATU03u
G2PrgeCbuYvR/HcgEoafq1nnkbs6DzwBKElbdGgcKtxGO74gzhiHbtR0K2UmumVgI0ik3v89BbM9
K2J+xlYGCU0K2RNNAkOE1WUo3/SRCYOlkZOGG9Xlzj03xYvi2Xu1UhWZvgZhlkTuz5SD+MAqaygM
4LJHQo9klSSOIkbsP2jiQr/83SISM16mhaHWvEPdZtoHBcSFQ/i1+pmpvL+Zf/QiJdVcVjbAXPng
S47hL/yF9aCTAoQyFxGGI1t36yWIiDk02g4cX9r4RmoWd7Ijx06g8FzBtvIqVUCDfZKfiJXplgDt
91dBty5tT781Oo4ic+OsrRnzzx5bZPIKagNgzT5YB1XVjskp+YcPbj78BsxyWhHOHrI5E/bL3qES
4kumC0kgv5182aEPv1e1fCjuXFSBKoyJscNLhcHJmTczjw4SlGogNb95hIqWzLZLLvAWLzzbgfV9
RiUV8hs+kYrk38RPWTg9U/DFR+qkrtui+wN7YEhnTRIXNbbvXpQB8c19lf8mtukOl110kRAz5G9W
8/NvvPBuB5wZNlx9Kr9AuU+X5Nsz50vRSNUCsR6S/wT+2/HPlzfG0VZxRBI7vccAGPNsol4Bzxs3
t30HMTwqDs7H/bhAsKveNV1EENAVjEHC1KqzQ/iD6YCrte79poS2kNOpAA+loEgLHJRUS+s7HhPh
fTLyYydDBP4907ZrSznkwShPJSR9N5uWmgVaFIlv22hID1z0GYEgXFY0zl1bRblHwKqOgSe0kkKc
HkjoSezBdJk0IHYLccEtEMnVmf/LUn7G8xba9Q3UeY5sv19JqYpuosFkXjl/eBdwye5PyHq8AXXG
X+BQAaP99O1EuGA5pqbhD8aIY30ZZQV1lnH8m6pFBVTBw4QMqvtW7TbazL355VNib5Nvxi0aD1Ro
6anT/Z0+VqZsdrKJmAuvsQ527E679GOXs2zu/RuzAQADQI0ckl7xF69JcKqekDpP+BBChjAFooi3
8KuwavhNNn36q5MFf9Sdi+y7WyIahGCPxh1egucW1dFPyu+5pvUDIFOeUP96QSho763YJ/4B2KXA
82eEQixPJXIcxv6t/L+UMlGCZcXVUTSi3ZAJmyGRRRRg+KQMGBf8LO/X/IbVDL5xsqZ4/sUh2OhB
Myiekd6d8uEoX3+exc4yQ3ZHnCy3NNMi7YG/JTCjKF+pRpv/Cqy1MYrKwA3XS2uydwhjOV7M2N/B
Yfdi4QNfRv95bhQd6zM/Mv7Scyf75YAocCQJxdN3nnOw1UZ/gIECFSpfSKSQFmKE/Zq2+BvO6PV+
R/5k5ZKrmgFVVc6EdXwf0WIuPpYRNNGE7HlXCsbSHoEmu+WVshYOdSTEuQOfP3MPuKip/ODmGPsS
IusTIJz4AYMA38kHhkq+bgN5E2xcvFOP7euDtq8eMOboPR/gMv2NotCN1mceRP4NYEOl5fPPgBIi
iQg/jw8p7/v3HKBnzQHScbGkJaGFPclVzJN88SsBmOyIYbFkq2kIFRT3HKxzEPh12u/+5XxR0A3J
nWh1+6B9LIOlsZB9lLTbqlOYZ6/CMjkfgXnzD2hL5+wsCnrhF+8V7NSaZ0hbWa+zGxio7qWEbZuz
8O/cCA8M9fyPCZq8SOFeCCVciH8tUHOt09IEyxvzEkrJ4B8aWRTn2uN3xDdA27rIDCoV5oX6vylc
bDi8UzmNCxBa+LGFQ3p+fGgrajmK867PFxYOhDnNuuHaiucpqgndL8laFvM67uY1SdSQhezPxhlL
ALZbrSaxDkb+wbxIExdNhSa5nxSWsGM28mc2S6ql6yLoezrjnNYq8gegueMTnNLU24vPYZxAG0HF
dF4JA+7mg3/4aMO1iaJ0WwHlk/6mBOBPqlzmYbJenOpLiuSCpm8FLnCNK6QyHpE/h7EOS0VEKCxD
Dy3j53RlPybEY6l/+Abu+waFiOydhwRQ5o1wI7LrrWOFG9VAt0zU8viHDb5JA97y7GNNG0qWNL/Y
a9wHC0b7FwGVHRDEYNZppDVBoVVv0dIro9da+4AdrJ6hB0KK6CZ9yiy1tks9ztuxXtryHCkOyjbR
NLSXnfCK8AqtN1gPgzT92RM+in1KCnfHiOwLFdqLwbnZxJTy8RSfuCIODRPGAOKKaiMzWIgaQ8lA
f19ljHLrgpairetRAi/D1Th7xxF65Yk9DcPNUVqdfItJDejPFsji9zRZ8OyYb1jj26BGxxqUiXxQ
1zJQklNVVVmwx/2cwEwAGApoe1/qJQ/F37Y2ACGky9+Bvj2e54pb402/u7oJABKQgOGERxsVPenx
uDvgM6EEdrGutTdkBbjN9r7HsLk/4Xr7tXlddQEsJhZmD+RE91NEWJ4HLGlUuY/O3Ny1MAeD9hBG
jo8lzrgZzaL5MNY2C1WTYLKwTCEq+8A7hibvNtGpEN4i0yg+0vLJARlPlbnlPeBBD4s1SmSBfzvV
4oHLhQ5jRk5PUyE3qZLvGBLwQ0t6MJ9aDIPKiUwxA1+EkCxvLzmyGB8XSqS5npqvJvGze6lCeSQp
DwiRcQO4saZ+vJHYmGgGDWkRW9LO9BFPl9X3FDAGerS+F8OZ5ZPSMGMSar1Ck/+xhqdkbHUNfg7U
MqG27qBN43rDo2Fv9B1dquIufhf4Syfkft0ZwCjmh5LSgoPLgPJMiCeSEi3ra7oXF8NtA6W7EPkD
FDwhhDddlAJVJviLHkiw6yyUZnkuW7DlVezTGvBV8Hr0F8HPAc+Ua6FRqRfZM7KbFPnQKjGlcw5L
dQIp6tU7RqZylD26URicrUlR9l8rX1okJTTiYThD1NmtPX5lHykxxZKxxKgg589JtifOP5H8aMgw
P2zIf6GYuka8Lrg/sRgu4R5UAxunl7dDdy2wI9hH4pPpEAjlauq5jeCa/g9ShmDrzogRetwB72mI
6KJeEbIeUJuLjEva9h0nJ4Tt7dC8bEc8GvM1twe/7HueikR/Ao5FZC9Q0XzGd+9iKz+IiXsxPXf2
/fBN9aCLO2LF0m2C3wLZA2nCEXWse2or0R245YXXwvkVWh/pthE6qDg2ZsNs7eADD4qNsTjWVpdM
1PkLQbDyKQiFRAWX1TlmadQj5SKMKsUn3zhVE+79dYw4YraB5FTkGEbKVNvMIB2YFxmNyFaTPd2a
NdPaEJdWVazgfvLQfySaIjVmqZSY3W/S/nYZXSTxndYWuN2phSXHVHBFAtxazAekoYfF6jKic8Vv
rTKZHU4oUV79rDT9wrI0GM5f7chHggTICQ29SOGtc+9lZKx+nxUV3BnMCjXYqMfCT3I4S7TLX3cC
dsiW1rZPWgdmWKQ9cvsDtRroiTJLs3X1vBXyCG9FqfWFsdYDr5MJ07nIKvcqeK67OwFjp8noO8L1
iS7CY3MT8SHgcfOPuSt8DYu7prqFQz+fLkr5Nz6qoZfG1+yzdXWc0RP6sAnCj/hfi+xaGNaUqa4L
BhTnCs8CnhB3ALqMF2dPcWdQ54kgrumXm9McxiV/Do0Stx2+g1iPMOMt+g1DvWM6+NUIavvxF7I7
dmDxxdiSHk+cDFDS394UnRTedpXkhTmTJ8hnWOaEelOs4GnCOD+llb4JQF6r4sykhpc9WeaTk0Ha
FTOjo4uJXHAgq5cOw22+TcJDBtbZGd8tCHccgt5hrRB9tfPBdU61JQ3sJqIIYy9sK1zMeorB3yL/
7PBvEGg6IbNT0LzdHDxLL0l2nqRASWvWxkdgYe3K28NmFia9l7qskNIqcvmj59FPh9QjaKA3+Xo6
Rn/llJ3nVaUC17L7OTANp/mEjPFRntEyXiznM3OEvYzKYscPoBIX4BkK94emIofdVxk84IHTdGZG
rE++CmDImWrTdm261pD1LCd+aaw93QcEdWzYRq4PP3Gmfjb3a2XW9ErmGd46cCuttLypHKkaCyMH
AcshKPyZUKp563hNFeYVND/EGGuELYsWWYY5fxCA6GsEvCA0MydNoOkqc0lC4GGUqImKq53MW1ya
RMe6iVeLDs5gYSomFzBNr/cFXmuKKwH/wNP5J+bZx75rGFoDWqHg2GewvE1b9YLWMovZCV7mcQb+
ly77/9cgw9lp2ZkfmztJRPmkvgR3rMfSjNd573vrtzLaRahk/kjC8oiXttT0NWNRtqFBmFQhJRsm
+zY/3SotA33C02upEGcLxo/fwQcLQHIugNrp0z+TFLvMGvVkF+REzmHY0ZSqJeevQIVI2KAB/HTJ
Z3BEvqzcM/Yn9T5/37vRHZa2BqvVD6fBtULSdTGA4QQk6inmpgwBPg87m++C3B+fP+Qh8frFSpFq
B32iOenu3FQ85rT3oFgYtcskqXwGo0Mm/cgBzrmXI2V2VKmlPDo+ayAAn9+3E5hyeI1X7DmfsSq6
0Mtab06D27upr1tAI5jYraW0XU7SDUD9YXTumtwxJ/3AL1a/rkK0BLFHAYAPMnuQoFEdytSOh6SP
OHm4cAIyuhVSUcmg2UrXc+xoPrB96i/ltYDQW50Fi6RDF1WAY1AkHeKISLcwsqCpAOa3EsvXYT47
xbCR39P0di2jNKLvCQzhPIoeQFVSXzMThwZe675tm975ivqJ7P+xvl/3CjMat6nm/R14JVMrTEZP
Z0yDZORPeQGC9J5ykt7E6NcfAxU3RR36BsUkI4vkIhwNVuZPWHJdihaf7YJf1+2qxV0yggpe6acl
Xpq5ne+7PRt8vAwQU22ix+caLuuJk1cCjvbZhuKbqc6YeMvZYob2mBFKHSZDnpQQwSgFclWO2UxX
K5tLLmYtAlZMaXQkjfmxBh9VXiE9ftN4WoPInh90B79OYY+gM5LKfFw0/siXBJhuNzkPyH24mZr3
STxhPitkBSr9qFrnRiIp0DwQZZNywzuO8U/AjnEpPBh5ErqKdpBAH3uutYMFEjelFwa23Crp2Y5W
6+7ejPXai3BgpwE/500e7hZwT79WfU5/TE/BWTHQhilQv7mV+/IcN9/L+3ZHNXUMBuUxfmrwEU7g
jwWk0srPL3Hn2c7oGjipEO4upJcw5ze7kMR4grSqrmC0HuN2cyQnrmuIwUO71ItAwBGY//dNB2Qx
vzwMCcmqcQ2nGK7lvQS8YT7msKDhJgCKa8/s9/ex8TZ71WM2/cONMRnS6h9GVACZrXanKpYpz9Ss
DsAqrDZS2mVP/heU6aFmaER/Y301uaTr8xHIn1G/lWoxvIelfISxf32heLJdPL/e+rfXNlb/kz45
TkA2n8lukbg8knmg0UuJZn3EkzrV8pno9T/B4sxtctQvEbZhSWNx9Z3TzFhHvllVYiQ8yRapsrHo
FdDDJu3jZyXbsaQ1xK5MVT7u8jhF9mdWw6Bd11mKVSYSu2fT5CfKSS2e9RrXMS47ZrSkU/4hezW0
m4HZbUipgUDgQ+MG8KIiCqjeIxovEPl630tiuMwbwkjZz/SyC3rfH5d9BIsoC/SCr0m4BtWZ0mvV
eAwZtJ7wTWftcL32UhsUwvVQZWxB4yDWsLkYErqN+YUGDXDLYgITzJ8PIjp+MLM8Av9wwFyv98ep
u4FbXdvogOq71qwk+DjP1HqaUiHwQop1+DTfg6PnQTGRhWf3WXh6i8LJTv7eAuJrNdTxD9tLbgax
Gcf7RH/NPvib9/K2wn9XZZyOkqdY6QStaC0LZWsHtTfhVA9JjtUSXYZQP7a+7E/gPSOJ5b+PfGoM
XXmtEMvqbwT6bkyFRLzfPgP+BN7hVogMBti0M2RK4VUMtN/I1zaj8XhMbDqP9rsN04zt0CqAkBRx
Bggh2Lc9cpu6rY62p/iOnca+vI5CA1/5+vo3+POeazzLepg4PDjWPDHBb5TJo+YKv9Weg+IdK/JY
JFysqOWz2kOJUpeZhBIrXZ6UyycW4OE4QttemHF8q85MRZzjWPh2bssE6UGu111xhEDRTG/imrm9
8QKJP7r6FkaaF644g7MEWADNJPI5fd8+O0eRRBVmAqufsFsqE/aeJw2UQMbOZLyudXA4yODu8848
NlztOo5BOEYl8egaVGOCEMON6aCkIABnFVBlHfYqEjOM/Cg1SKsW+mB84XFfxh+TDBDrn2gWw+Vt
2QWODFiRHVuCzvak7ep/lMebzVSJ3sHi3D/PQWbWzSLmOccKhl3AKH5ebqihLLKqHqBZvdNWL7Uk
me0ncGsyWUe550eAt4EEAS+viu2r8/w75Xuyd9tKRc9H1ipL3bnmvDNo2E7Yn4hoAIbvFVQN60HA
ueMyC2RzuaTTJfEfUxX5qlrk8l2ZzCG8OLSM4cRB0n06gqgIqdTUvCRQCKtYYFYvnugLEwk/ZxXy
obV0YynbB0TI7cIlrnBF8ncgpCXzqo2hALm2567LmFzKaGSb/oNfYM3WtgodKu/mUm/xxF/OcPBQ
p+WYYSlwxZ06/4KzOSlnr4DuM4nJij+5qSmssAY2k2W4UQk9hPsch/97tUXidraIwABQA+nGLgW/
13DPiUY/p14K4AI9ADt4Y3aWWHymgCCfPY//w5OZbghqk1Dq2fHgWBwxSr8K0jB2qremfuqk1WJE
cjdM5cqZAbLzpT4i9CBheedDBb+Pw+RxCc3lequDMrr1o7VTaYSXCNUQ4Zndbuwfx0pvtWLnQvzB
gZ2wCTD4WzmFuTm10HPsmuWhBuZGGTPaPpcZRd17MiPCJHLZ8gOgnkEgP+G7y3BNBckNOjGVDpr7
sNaj3U1D5WTBOQrnlnJq6gQO47MhYG/DMGwyFVTpPfld9SyGn5hrUK2S+LQ1BDPPEN+EU8CcATyd
/5TpbEmgG3pZO7Mvqb8jcFAa6KuJu9LF/JhP9VMn5LA0FjAoIvp+DgP2RwKQvkRew+ln6RGqhYJD
7KSseT/CrtnsmMI3L+e6Tm5uUAPyoDHgSJ+HdeCFBqQoeDhER0udbBf8onrKPJhYz8AnXG1DnE1a
/knSq7Z2RNGRF3lym2G7j6fsl2Ltr3Adh6Yu8p4iX14qLsbQYxneA6ScDl9gVeDVftvSSdVPz670
oczuA0Pf13FMPx3yF9r8VOMh+2V/k2/iSSTuVb4lxstmgD/Cp/zuJH8RHJmjtgqZXWS86Odj7JOb
TP39iJB9AYylT92s4JCywpMuguHj5/spsF2/EOYHLh0bX8ti/GAfPpDZFWWpYKmiz8xW2geXM0Xk
tjI/TceB5MLpRAlFer9He+3UfD47grbq9wqwhGNcnLJvStJo4og/PC/LL+cF2/V234AMy7TyDCPf
uyvgBB8iGa+dsQBR9/lr7PGKbdH2MLPhoimb9yzlwCQsOvTrhc8V5UK29gTBtvnbL6dt8BNLMG75
8vEkwfbdIlGo7HDkaHgQH04TYWEgMsZ9eUS7QicPFCGj4bn2RuecWOutwUKI0TAVKDK84S5IqJUD
NQCMHvFIMdoT6KGbSqepI79W8dhlYFzT9rnrc7bPwYjIR/cErLa4T2tm/9wBE8uZELokEpVQDA3R
E9XLMkcnYpN0KW/rTESKUhg9YjzreOJRSFftNo1vV89GmaS48PYqAKx3M4rqQxTmufN8FZEN2off
tTa5e0rPQ/whL67yR8uvTp/S8sF4r/BuGzsXTR8Bo81LA2h3pyu20nJtyxTE5FOfW9kF1+dGsdLh
BgPy2r3m9pHujrA0KMCb2vIPhwmZpAdDavBA7KkEGRE1RJFTqM0n3IgWri/tBjC+lVSwrNm0jGGY
QXUSMkChFfwuh/+fSXg0+gR5uP+j5y7JpiarwdcZ4wjzw3aP+KI5TXS0d1RY9gSfre5CG2LuwOCy
Eve/zYQYmMTwzNXhJOKkLgsYULxNnZ0e875UPFkq0vKtejxNqLNRWJOymZeYTopcQZpI1kTxOZQ1
GrVCdOoOLvWSFZW7L9jd4X689nhB/wBOCio49zrMkZiM+IE8aVqgSdhuDr7PZPvQpANnfP6UmW09
xvC+7Af+Xg4pjJUAc/g8eCHaJVJTAP+nkPabQZeQVnHUpkCyMHhkANbP/DA/yNSXGrmJAr3vZnrp
AOmaHaU3CQlKn2IMqR7Za3E5hybZgtcGHXBPYUSYouSBKv6OD8nuDTCHPxMdKOxyH8iANJTFN2Pm
ar3yJqG7kqkVev4xOzNtCeSjtzIRU0aLkQXu/tlAuZMoVsoosM/Yl3lRG1xmnu91z9nVeScMXf0A
sqtTMDnrbrfCXsGqvhBie8N+cGWQMFFita3kCbvXQ/rzCMZN+V55cG2XkSjXGTJBJjOTo7rpI8dH
CB8IoccVujkVYLBCrWa00lfzhzDlXWxyRgNKIF4xjO4BS/5vSVmDwNjzBbPt40mGISmjm2JnPbAN
9jkzmGC/jxIw04zslo98/iMlN2sTnxxHUmxFWrld2TFTt4zFzHB8Zwzt1w9zWsiTSKk1UaPaVb1h
SJUVictxj6pI0JR78co2AFhkkDv+AnWJUkk+uchCdDd7EmVR3wsHxjPDf6diFABXX9szhtiq7WiM
ULWZ0SLBYYN3zeD6ByzxFKA/xp5yDzuOwOb9R8ApMNZf2MOxYesnj+jnFxC83b08PKDcL9Utfk4n
OkaZMH1FDs6mLrxtr5Ouytwxcz+CS9kXt1LlI0okxGPoBGv/7I6my29wNnee/rlMm6uE0+SRrU/w
ZZC+gD01mSEWFbecLKtOXhiuZoBgSaXdG5A/XMlROv+S3vTFF9lFSJ+L8iCmxLSv0msdZGpcKQiO
/FNbAp++SX51cv4cfXxxv4l8Yk+Bge6nwBCthkTgfQ7dZDkREoe0q3eJDr3Hrqfm8Zb8TYNoIdoG
VgcgkaJJO/UMYoLgqTnCkc7M9CciurbRbiLRGmIv9jyLyCoOqa/jJ5e5Lk9+zqswg2jP6vjCRARn
UHy9S7xR7EEr24Vutp6hShvOsDjXehCd6+43n5o8LNPWAweYWgwLQes2M3P3D1q1sNLsztInhlbV
0PkE9PoCsAv/k8gZi+ZrBfmIPLVWA2mhbiLRCjyraI2Na1dRV3DJHIpSDtnMi4FP9AWsL5mT3dyz
L8A6yAQNnaXxwtPxj7N26u/zOizheF7Wqsdjg78Q4V8D///QPKpIbj0wH1RaIu717f0oU9MgvB5p
oWZJNxnwZMTqj030ISSzJz0LdUlx3oE7Y3BLpoc8ZD4RBOFXxkivHqvGIjxdn8+9MMKNcx+pBXR3
Brz7RgUn+km3JISfdPLq6pDvB+SgvbhEAjZHzxcl4eNcq2KB9QA27PsOkHBenVc7hmilfi3FaVHD
ew+uVwR7aI05OPRPFB4NaA70vyURSuSjZ17CazleBAvAcYoEIZIODQH8JNYi9wru/mBqk0wthawv
hyjff/w3N/uyDV7vuJoQ6e0LcMgkSR0zIp/e80lA1Uz03OIb290MyE4IDXnBEL+K62eq+QI+krHl
K+dq71mKhAUTamgdiszG37C9Vym41VVF3ZYXV7ACf/fgdWg3fcfdGA3mNGBlFayDHFMmffSvUaOD
OCzuua9iAFEPyZsbgIZljpEKPlfQJ5BGcSjKXS+XCYYQcsQX64bGGsEwXu8R0gOZhXItOKVLDdhe
MIitPIbEMFKGRC1F0CO94N+uABygSXkMaatNAr3AsEWwepui8SkbGpvnnyEBXf2kRrz/pQvl7eb9
l7r5jQsnv8Q2EfW62CbCq4xOQyYCcerYBc1Oj/lpJAUE1bFMw7+ltDbCdDlMRCY/QuGbVDy54CYJ
PiADsC6ccEWFa2NrAd7L02IPDrfv6Hn/CDW/zV1LwmwRy2cMXtVyIJkWzhYLWnOf5y2ENCWBwsaU
RkXsrPlNkY/EcXB3hWneA9DvavtkTtlratbFdhoPrCzxYXIkjPgXqg3TfxDdrNcCXZshmyOXhpCk
l9W6vNp3IC7xF3JYUfeOJbpkbXBT4lKYhJSeNR0rOFHt81F/yezi7GXv3yMBgXrsg8qR2xTZX6FU
mcBBQvUSlE+i7bweXOOZlH8gv0f2KzMArv6ZTeXZI+cRTRJjfPVPniA+UMQ4aCuNN0yOS982KXDB
OzbQ/GhLW10wWGoF+A/ENPNG+B3tQb9+RRP0vlJVCWQX3OyDFElTGmqQdRvBxIET2jO82/uUuFAs
a/FvRl7hyNeb1A6vJMIrR8L7c47CyPHCE3i+Neu8QNmA1NmtAdUuHci+F+QGQuCQDJbXXex7Snr2
rE/1VCQrs6rutPS8CawYX+05VEGnYexr/vWW1KBVxpQkaLprcvF+5EVROhnN3C3z1JGkOAMQmyBf
WErfZRCspZEW4yb9D8aEBr67eMD6tB6Xdk2CJQT/gJv/RChjXyP9wtgGWmTv/LnWXeGHJZZM30NU
bNE0wQggqAoLB744QnTTi6Lr92tRD3rcc28F3QwdWuQZrwyNObg6zyuWe9pii3ymYKysnKUqUywP
9I0jFIIlG/2uu3Hpe524ZPOJGBAEDrCF4bz07dmAJy6bspYBBdM2/BA8/9ml9MFITjSIStM9alyu
AQSKKupK8q4KA5jqHFja7/vDjTsOBkhqxOpa6pQInAN2Lsq+ZiN14WUtITXowiwHslL47TdFfFaf
ICKScFOyUQjDPL9L8xobB6IvzIwbWVgNC8dJqjYmevYoYqmXD7ASCi/F9pGV3Ho+qbtPvxl70dp/
PyeQZJFwMGwarcc72otkWmg3qX0NtYxkXrWfNu1NZGOHVuPPuUgsiVtD1YYjbryAHyBr0QBfNhjr
Wuneguw6JMSF8ATJX5yjZpsXXXMY6IF6MQNh5qyyTyYM3QUlMT42SdahxX3+6aEoVjR8Y2wByBGn
3GahSPoYxlkvWtkQJAKw8ltvd8B6SBtzv8KVg22+WZgYC9bObvXJlt7fEM52StU0MW9RNO7agNe4
P5OUdb07tTqJMqi94PO4k474hGq5D24+RBBPJRXvC3K50ZkSjILk+BIfhsgvGEcFGv0IsWcgSQBK
uqRSY0/0iv/NBLVFyAa/+yqxDhCu6CAerRl0e30Tf5Y9KICYz4mbfjiZPEDBg8orV+qXsjyZypa8
rv/i79XRKAts4KXAJzBSZkTgH70Md2C/tM26urxbBoLfIbqmO03a3rXU/k1ZihA32/ykB7y24J1S
aLy3EnNeTOU1OVHliEgK92xaZgk4WggvJCxNzXp6Oq6tMo1cC5pDkBKi7qsq3kXluaW752L/zysF
c1oVUaHxZSQGAbTTdb5MdTrk+SUu/DjZeFh+LGlG0V+mFvukPreiXIlfPfgA8Ls4bM6QEYFRb//Z
D4OPyS0DuUhiNF2+TrnhdGMOIvgrZ6GTiy/AyVD6btAhmeTrmf+KcLY/WrZan+eczTGfFPFu5W3x
Ii5z7NXXbJayhGerc68SSIz2omZRy5S9/2HEzKSdf9MSeedrOhjSFn0RuNkul2pEDOf+SMHZVy25
cxsglOLBXoGfzjGM2PTW+wfmnt4Y5PtajHHCzWm+7+XPm3u2zfcZKnYVbnPj1gslcUQ8PlTunHL8
sgck1WN6gEK2KmgWWiasCnxo8Ae75uOwbkUtA6f+BIxwqSJA82pfXKvsCkteQ5+e1o2DtTvFQsar
Li96WkdVV81z4ZMRClxaIW31lK7n+rB8evaBYgOL7N8WQ2U/VkUS+n2SiRAoBbFoRLrGZ+PkUjZv
9hKbSN5e50SOrJdAXrzoslAID7sZnH2tmtrsm3RxHBRk2PHe40apDut70aAvWYE3E0T/SbBG8qv1
YydPXuQkNEQL96CbjkDnxjJihMCtdCEFG3Mhjd9o4hKpDs81SdxHsEZoMWVpMlBTWKqNLJ1Y0Rtm
fj8xoBpcFFZnMKGvLkOcWeSF5X2v58PE3/0mAU1Xjt2xs50apa2DZYx/XIQN0z808Sc10HiDIJS/
Vna6ID23BJz5P5uEFXfcr307XdaS7P7I5nqPfAJk7T5wpuY4FI2TZewffOi3gKoib7azbnXzwXWY
7/pXCaXsyzicno8ZoOnmj8OryBzm//WMqGHuRV7KvSzp85LqwAa12igSn/kCUnxq2TDMVGNgIQNN
JNiiFFK6y3ekKw99DRY1lUCVdQwUXkw8tVrt/AZYMSyxu8SIYCxZNppgwtC5Ybdlfv3Sb2amgL0B
0LNvhYH8S0g2ZVajfGFCZv+BQvbTnuYqN3RIBlJSrHctBtcNsh9XH0PUymicUwzbx0pGfFHGEtS4
TikBlh7iOOcBUx7M2g5MCBDBz8GfuhGzzIYej9Qj1w4ExYLQ3c+gsfTzOIPf7a/Z6jqoTpo/0N2v
cdUFszo7pBOYsh/sVVSQKwrL5YwHdIc9oPZy4jhWXN370CFZGRJP8pnJ+SU7vdYTtbiUbxvtP3hR
KY0cHbDrbzoElDfyCZ4XWVzANl4lwPlyWOYPdqACNGtMzJ6Eff7/nhsEzACYkNuyHHStWP6ltk7L
k49MpTy5yiGmw1xdf6K7y+JrrFmPNChR9Dl48sh1U9nnQMg0kryydcRj7iC7seO05/+1OdMCi2ji
4xXtfAN5bkQ6XXvJIfL1AHekXJT4WFRA7COKbXhIozLhre4yLv+9R92DJuUIhRx9DY5ohHPFwgCu
khMFTY01uMumlxSruQ+jrB6/d5rjAX34s1T/uZLdZ3yCGrg7Fj962KyJEFSLT8dur4uxekIMSDCx
XjCn+9r9uifa5xCNoHFw+qmLg6+nfYouQt309Jdh2aERG/nBYpBrTq5ngncdY8m4yd25agEtilzx
ocaKnDBFsQlXFGYkpIexnZg+9WcTAxlme0tGxe974N4VpK2AjCYYN/APA/kF852kQ2vKHIfy5O1c
+3Noiqyl6AAz/z4F9j7dbKo5+xfO2RYGe3FELPZQh7iHBW+3gY0Le58cTLVS1gNZmflLf1iMBo/C
ChKO+zNGLCgo0itJZTgkYTTNRyfYG/OlBWP2Lqg2uiHhz14m/9yi9uw0iaKww9e2lwcTNg4vpggd
mMZN+TNXBWAMBO8Stlt4bRN/th+j85DRRk71db3cUV5vuZUqacZl5RxzVfhHQDLFvtIa/hiWMVTJ
nDJ11BaA10RJkwi7B6u7yVx7Tq2Yv524oAr0+yGFKB6xpY2Z6iTviH39s/Ioa79Nepgm23scGLdp
Lp4XJgxUgt2rfP01OAjSFFzDM1QovIdoGxhDohCj77IniOEsh7/feqowPh6czxNujFzpQHfjoNQ+
67Y2yFDbN0Y9rOOyjQHOgw7LkAhVlEXI1zP3UxSfE1EkzdvsAYHv5yWHPH2QLJtT/BxhO45T1Wf6
S8wHhI9/nlEaFnt1VL53P9Fh0/CfDfqkj8Sj9q/qHIII8b3SJhP7oLG36vHzmBEfuJeTnIvREutM
W9YY2PbzshZFFUuN0KvOR+UjfD1Nqfsu1jCEW0msKDGcEH7m3bfs74fpRQywL5L+6yRe87Mc74TJ
E9wTV1SUSGdBBfjfaKurMyIWoSR92vpfRfN25m2dcQCdUhXg9BD7NLVL8jMQt3yC3qCr+2xzB88A
d57dGjAc0kVwqSC0Mgcp2I7v27ypJFIw6RLDWzs6x3SvqGba4ssf8IB7rO0TmFD5TKUXlnYKvH0t
FJGpfzxTeI8Yh2TtCun1VzH2poWdiMb4vM2Q9r0blloVApQDdS2n+cUzalwkRqN4ohJnuiaMrxp7
AmbC3wwxfIHZ6NHeV0XDpSgrjruMqEU+y+5BCGygu+2BHo9Q6RbYmp2BgBh9RvXTvx6itGLCXyA4
57Fx/b3j448+OgxOoU9S/JgMw+ppSqEP4/n89f846Gaw6iftoSzJzmnNMY5aDbdG1Ah083zBxa0F
9LJl5e+ZvZpAoyJCCFUj3+JV7o1Iz7RfLU8IAmD3HCQh5nPHp54/IPWFfVkwYcB8ObD6PAHei9rf
pgjDU12qYn25B6zotgGKmIGTfAMb6fNW/3mI6nMuBra8RrSot7w8zs94ZzIb35G40+CaTCvocPhJ
Gemv1jquOMHnlPEINt+1UtsTtD1KNpQgWOvQfCkCdQDW/deTAL4+CK6JIy9cME7HjoUbhXb5AtBd
831jbSX3OhXUZx6dr/M+6dR1MvvVIIM9XS9Cw/SGdML7AGhv7928tREeLaNvRdMA+TE5htrVXTrM
8wrUDGq5C+vIdIopfNK4ETafihmWnrZPI2B4QGVTWob+EwWj8UuuDmLM66Xgp5Mz0zbtg3uqvlOG
+OBvsmxj+Y4d7m3mcVb4XhqT7Vabhfd0pIyyVm1aG1INPu1cOxSxpqCVCrymbTp+WVXMwp4i1o7i
CSO772LazZhVWT/vWMr7pnj3wOZFlB0B2KXp4GLRruJDpLRgi+xRoHpMnowXLDK58QUozcmBbzJ3
uvQomNHKvyW+L7a5ahdwxUfKtvQXGarVjfskrU2SZSXWPIURjRjwcd+HAtr+1cHw11PiI8QJKogs
JmBBOaD20IOaeuJMEpx4wWWdjOk5i/YYH+C47oU0NIpaDvJgLV3QnNW4wFMj/sMkhkuVAiRZg/OQ
WIk4QrcIxBfxvtO8bSVcIFg0zl2TDx7dfUyp1ZpbJv3h6KP1CLABFrTUkxAwusQKcc0rx/SEW+nY
YTTYGjpxbwmM680C0M8ACq8OGdt7O46iDYyBY8fP55mC0neC6gIRUD+Ox1/hZg/OX8yLJzXd4TXV
HD/MTHGU1ZDXYa5RGTXD3FTZv8FEs+xOhrz5H1zKf3jvlPvYbD1U/+6jq9jznnNqBZitGMqPudtN
+1qdwMwEF310Lf9nxzGOaUsZ6/wa2toyF7t96Bo3vLrCGm6msQDMH2tF4Ku36NKoQ5LuqpaV4SKj
Wi3+X6HHvVbWiOfkRdE+KmhLuZgwLdBFYhoJKN5u+PJmEU6VQP2CWBaZk66oOKK42nnKVyU9Z7Zp
vpNxx7RLR4tZyNfPKookbi6gnqiZRy4ilG/e81ohbuRIkJVBR+YAlMqdADDuEUhVMc+XiaTI6ZKH
a5XC4s8s8Ex/6+07LWLTrrP0EdxNJlilYOj4S7KsWa2rrCCiWCL23438/ZaBPLWyLl2+mvaAaGh0
ZwCUcGe0f9+RfjdULGx/CZDMn1m9M5Q3k8X43iKe/vgV4KRS+fMTPGdRFtX3TkaUfCGxshuAwA/D
NA/UhZSDNy1rUAmdvDSefpDq7Vf6EwpY3ofHiLdUhgQ/8eJ2c06l4AkoqgZVGgJzlyT3kH99yGxA
sFc0EzCWUrfQiDnY6dYu2AW2giKnapiOaeDCTY6u1tckPKF/iilIzW8BSdOR5vGbesJJTzPuQiHw
S09guCkt4ifSNOvjTtvzBXrArHOr+SE0B4OrF/Y/+K2GYA4fJWBjmoZ9HhvvIB1+N1yTw7CjLmL5
FxhTz6lzFEjtfIbfizjw2668Fh+c3qGs1RAGzCUUveVfQYSTtHBAoQQ0KoAIdlcRbjf4gqrdajeD
NKx32IfYE9ZQd3JBjKfsW43DqFbx/qEtSeWzDz4MF9rt/gf1RjXwfZOw8LT1TVdMwWHEFdGlIPbB
Wuan7D+YFrA0qe93OK49zRt8jccsxc4cL9ai1fdZ2uEx5RoOSdGoaqTM3lUZ3VNmpmyWEI7tnV71
ObooX65HkTqEb4ykR0r2vfQrj8tH7V6KrvSMCPfy7r31e/YToP7vA0UoYIVKDqVa5ftviw7TEEUb
WD4T1yH6o/wzYA5WQ7SUwW1d4glYYLks7j65pdJx+RU8h55OgEOJJtOXVxNevkUIeAN4qGaESt0r
wZs82YDkPXqk+QcKOlQkC0kEniIQ2aghtmmfCGacaeDCqGlgA+AGoIrj0xL1O0H2Re8r7GBkFmWI
C6npaXF9chVSLaeO1wIvrt/xpFA4Yp+ZnlFhtp/E241K7cACWj5gLpGPLPYQFSh97b6AxR8Ojie6
RSKsFrYt4IKqNrnJaUYdhcIPWuik0VkSCoNzitzG8EGSp/DwZBH5BK0drN/2wSkzA5OGTw6YPS+b
T1wUKDdZRI1oANiyb2YgErEKt/Wr2V+HV1CISNVCeYc5IqcnaLDH+oLkYYpn2JTsjgNs6gT/0KXY
OZgKLM6KllpjAVOIX8HPyUOEND5C/0T4B1NZPt8uySu3XWOl32jTtiNh1GbnVffno+IFmbS9XJ5x
CRFDmVOeSnEmuiqJ+YQgYQDBP5b3gfKqq9a4LWMbwKNj3htWEHQvGsDVDIlwq++kHHjxNC1vxquc
gQsXjL0xH++6ZGC521OPHeB5R45kLiFux94kYEdhcodsVx3rL0q0rQycwharHzCRTtikMURG/3UJ
SJIg6paa+FrHLkCuuLGJ4aj4jBlaBIl0J9HJzy1j6QoBKSpASMedZeUb8IKhulpKNHj7AQytISoM
Be73Ch702lyNqbx2D7Q13PgHd2j8ZieMlhmzEH1MDH+plG1If7HHOAbZGj5weyVXToZlMHHupH3R
s2vnMlhfLMro+aKWcPYPWGMEczwCyUpXO1SLTuNZotV2v7hHxQTWmrK9V6hNAjQlxLGmbeMelAoM
0YMpINiytuzGmkGTIdN6LSOWbuFi/UBYJFYxGYMyDqrlBj/sXoH/BlKwvfbg9RkEOufuydQ/zGyE
3sSRCCpbi3DxZxXfIXblMkRKvP8/ew8UANjfAnAcAU73aRX8gwh7EiRYLRwBWhnZwf/y817XwhMn
f2GroOtHzeH8Sm952r8/zbcFO9BO58jLi3LvldyHeHFQOWHIaCgNIgSHy6f4PGUvWFy2A5KxdlMz
leM47z7FOICs1xUSU67H6dGohlXIBDeuNJETqBycus9fvzlm/n0HCaWJIjPAhatn2cNYebU+aoYV
LkwrPjDnUDn0lK5LaFZZzUo200q9dVFERJfV7BMYoTzU0trnoAnkE6o/lTtR6jCeIecahB2vYsFN
MjgpgvmQWzBlhKPtm57vlkZ4U/AWeN9zyYdAM8jTMGcgPUrGk+QS54D6z3+GR02c6QQvZpvr7U+0
JWsWhGX389LEeyeblr+4oATAX4VV1rKtGiae3QrV1rI8gKgQR9W9VWozJcjtvRMge74pfnax8hlV
eNKqSFJftAIjntqmvsOlED4ghPRbwxkWUsbtLVSaxlkrXOmKMl077pXJ5eYx4yN9ObKLbJ1yZvHh
tR31hNJ/wohNmmUuONP8DsCYYM4wb77eA02WHPFKXiHJD4BOVax+krBQkFxWB6k96axNjSrz5vbN
g/GBNG96iwuTdyYDCmfrtAp5DCfgVohLhdJIwIeH0WvE4fLmNShZEjecVt0tG7++vCaa5QdxQl8U
dI2LyJdKH9Icqq4HZhCCDzxIjYaFIMU/KQeUswieBsReDom/u8Y7rl0Gwk4mCBcxJdp6+4qqt2+3
DFyFKALAbY4M+kFaZyXwyzRNmsno9Zyrh8i00ikBC7fZd6hXAq6R657zswKPAxfyd4aqjyQ6VMD9
AKD9bDyK8raZPsZixRXPEVeLL9l4jrOTiY6F8K1F7Yowht0xLSdr2Swmm24an8Ab63PHmAuPkvUt
iBiuXFvvPlxVy3UDEuFlxTY3KLTZZd3AWeaev6bSfLido6kA0hlGG5CIDe9Y5i+No0hyWBT7mJT3
AgzeGMhgHigL2lUL/UmWyhkoZ0chA0dFk8Ou4klp6nwg/+Af8937z01xjdzZtiGDhO+66g7nLnGv
PlIKlWIvpwCNUZuu4n1KdbEYgESBZwEY5NxWZ+sy8tpLeGmiKddxKN5QIHMsmIMLd5OR5Zynuwol
Xbn3p88Cm8XMHIAj6RuNYCXDxvD7oOdv1RjuSY88DRVz27Krq4F9eeO9KBeGGzj5TbMpLOZ+ujuw
xy23tmnTTi8vLmO/28MpINh3E9RruiuvvSBrmXhSiBlwNacYNcYBMrMSrSyGeZUCgdrvzCq55mIg
trsVzydV5V0ESYf8ZabbWkdn21B7TnJIKPYuIn8YhtsFNlntbGiINac9MsFhSmAXO2TQCBJq+cjp
Cvz2Yc3Hvq1AGiIkQ+0tV5ADLUgiot2LqknsB0ZrrKTXC9OQqvfnWPM3eOyJeGqZ8rVZ1s1smMsQ
rVt7C+prO2l85/vcgWC1aMuPGJwzk1qX0IlGSUMKyKdhBQZP6+2IGHiAqKmc81TkrY2oUQyy//Uo
VePTj0UV1H/DLv5IhNCDyWp/O3V05Oai3SXSAf+O7Xkw/6Hfc8+cMI1nFXPMAuXf0uIvmTqpV77U
fe/Qa1AmFFDM62rPftlcpCql/5tNJDLOUpebgzrSDQBtiPIpf67EVIueKCsykLEp8FJ1Yz66VAH3
1R4JpddMdYjxzs2yGCEaRB5AhvjiS/AX0TtO2qwF5DQAfmsf/SJ/ms/G6b23mmxD3Cy0raplw/Fz
oChtFLwy1CehRopuSIcKLqYClFJqtXEYP6tgtoOr/6Njm8Yq85ebnJmOj2dnOGfHxjTCqizM0qqC
5kk2hTQlIGEKY9s9KV2evhAyaN6F3f1mia87BWlaSkq/EHXhEJYsazG51T+j23UQE/+9Hl6tkuwK
E2ixJFgXBHkCPK1YlmODazoXfxfPjYaU/tUkf3PNLKCYKNbtGj5xqNYTk0iuEb73lcyX/0IHr9qM
Xuau5ZtrrD7PsuoqGmMg/vTRZhFJmqXB8ct7/63A8/nU0iQ0EXQljbEexJu6FVU9st1MdMVGYULp
IF7x+vnpvwFHIuwKwOvmisH/oVJLOZx+GvfaxKbzy0eN4wtiEn/4N+VMAf7TwK2eUL0zd9rcZuk9
122F+ti3ahVHW1pFGzLmwUCv9/6Iqvnd0spjaWhbCobJg3Qg5t+/iMtnezh1dfMd3vITNIyUvuHW
ljkpVxWiDjK3cBNJEm7tRcE1NalS3CEsPVRRakR11e3zhEL5cLnS1nMGJiID3JZdSnqlGezoISed
xF24wkvJLajKLwGl0bcP1JkcXbQiAzRdQsfad73CNYIy6OZxN+4oQIfhkzo5T9Q+3p9znnruBtE5
zQXz5iUurRnZqEZqRxra8lWqZJEG2FfpkezNC3LOQz3AOb2SOElyoTlq0nOUL7IR7VdQhfq+Ikb3
EBWbS/LtmA4VYGYWytj5+jyysBtG/w4zQceEs1op1ivl0tfGlckXpxUu7LQcPa8p/ha6xrOOLN90
qu0W4VvjnhdArI8r0mDg5K02Fx6UMmBR1mI61CSs86Ympj4FkNNS5Mj7Ahj8L0gFU0t6EOpPo02m
SXgHxsZVybZNx8AqF+tMp/aEXvvOogmvE6VsnqyzsNaYXrkH4FS3TgB3nO0CpANYizhtEKbiyxR8
Ss6rzX1D1xHd27tyvlzOomDxx2AyMF/R1qC85D0PLseNjes71oRZlDuAszqz5AIqTHVYoTgYsAu/
P5a4WJNEhmmWIwltT+HT7DgQOcgGMP716XnQZqMWi2ARgrggOmBMFvGkHUo+reD5PavITB0W6SDH
T/SFlxssasQ5ytFZo+q7Jq18UdCv5bWgMoXhLFpZ5rkyQPXPQd5BF0O4MNiuWo3FaCQJD3K54G67
0CvZiHZiCtIWCS7DEnFmkJ5ueKZ2beUWmBlw/GsFRjY/4JD0B7bGBLSA1bbOEDF/ieBVfQS0g80v
5GFIZZJaqT0YJ+jwjvfEcQ2b0KZJx115D36fV3Tu8NwVsTWdIi8zLJFzNb4KQEv4egX1Y6XndSdd
u9tKNtWgZo9wCAymSLgXCVTukJOzrHqTBuldFvbi4pvuJe6TFeSm9oSoAeEzPNe7BjBlR7FWopP1
1Trh0zsnxS7OtCGAcyqEAOqXg9O8VE/rrdxXy181zicART7loNlEE4g97W0tsTWpbmPY0ADuZ6/R
F1ogSOxKMOEekjwn1aK3aUITmDprULqJAuho0RxzMisDLlAa6JOrlLhke5qEOKPxShkazLjuVaLK
21irR5PIidQ+CWpenPc/0LEiKAnTzWAjh2PZlzmke429qQZg9EtrKzn6RosDUsSpbmRZdD9zhTTw
EA5a0+elZUXxrQYY8oAmABOjMNbPTdH8YoYv2FUgm0XXMop6PA0s1ZscdVU0ahBF3Mde7Zu8eWqT
g/GQbak42Mmt/r0Jw/9ge7FGkwgFz+DUMlfABpvpNP1Pq4bWC4bZ1PKb6Q3DwVCvtAUh6gqBCOXv
2aYbpuIpLJDf3J8SduPNmrIqUs5m5Vsb7AvVkfAyfButEJ9oESjoniA1Tu3TPFVmajUZ+XvKQBgE
w2H233w31WYntYkrIObJCbghH2ojs+jhBG3C9AWMhc6tjCoV2fBXfvEANNvTK9yLyXZqKah16O6L
3RyGQz1C9i1sS8M3P7FpKp6G6ueh1cKXsXNYxPNgc3rkdWv5fJUKPZYLoc7uMIcTOhRMBsQW7fp6
bgUwCx4AV/pz1qfe4lfn8x6zT7oW3IZmXi6JBOayuHIxsJ1vjFzN+2P09Stflb4BzJ0iKl6CzWKz
uvxnGHxXp7O7eVekBThaivDz1ihCVRJt+PUXxqc2EycBV8favLifqiHNg6v4ynTFdJvto1pDt0ot
xDk2xr5YZZIivhdH9mSlAkw0QX/ulJWodKAM2ZdwCHDHVsaMqNeje9kPNDsNpKgCYVP4J5SiFWX2
YBtMqWa/h6/kRgd5no3tS9Zeqjz4leq5XcuSY1D0sKWY4jJoC1JfWPDT/H4jkDlhXaoc780zHbfJ
RmviF+TRrRqrWaehvPf5tN862ZY9inSxa4YoBug3s4KlSX9mCrcRUDZoeHmLGF9P4ptq3jWCB2GI
d5Q6mUqJ4rqoCoxqqRMLHowkRWay+CPq25v/w8VKUcmmbAsIOASp42MPvgvMn8alZC31oP1L+PS4
iknLDlD6s9HK5b86/n2ANPnw+SjqspeJL3TLBnRsGD29EoXFlVPWWMg+qUVRYSHhNV2YWB2lq+3P
QVovOx1AbnRG0qFcusqkQ7FyztqXmGgA6l8i7y0mP0uHV1JI/dgIa8k3b7iJ2FVDsbzGSKKjRgRT
5nok16F1drAToGDXO19lv0XVhVDhY3ubrjBuy5HCKXRFDIA8hE3+jCGz1DNfEbYVV9IqiVFvaYFa
9XVciqbTLeeiI1gMTfFbk5qJvZBR8LhR2QaS0OgEKeIXs3EgMvPBPMCPWkQpdVNzx4On1Pa9AsSb
OyYWt4/R8xoZOrboWvLkqVrTgMef8UfjqTwXvozS7pZqR7bwnnYXl2Ch+hBqmL218MbWa/Vu6WFv
UD+ln9snHKhmvWdmdbmtiUNsT89YwVK12kK/UoUJzeTRV0rM6NMavOBRi5Ed0NT3Kd7TXbK9JH06
aKp1NDe0SqdSx1Im0eWUHlxwNLWodm4c4bHimRr9wqI5yl5yU541+UhdNeDjj/7e9sCAen1Eb/hB
o+/aWXhzhu2yNN1fbe3En+5VSgDfcfuaLHMijRmOjKSvzjoikcaIXiNvHyGMv88VGnQhEmUvgMDo
oGgmTyTZcp3pu++cQJo5YU0IU9czOCx1v2GJTl93IuQlkO26kcQmNO6U2Df7hKoOMCDrhGAs1xzx
qmPTVHOYXmvxe64RuMPpV6+7GuyN07Yg/fYbM6Sv1JhwTkrJJWQ3yWeUhKhPFWGRRiocV4yJIgtD
K+mtRM6UXV9I2ROPBTOfI+cuxxzswl5DFcodKxLbpbPAc0foUhEz5Cdl40z8A66CmymeylnDn6ID
0/uMT/u3bk3Mv30Yq/EfOHogy0pFzJc1Udbz8AQ1enANCLeqa7E1e39Y4RTVjpU6ZGduDd1FYnQ7
8PWKHpGQNW7B+NWtcgAdJ1foz5ZwPobBfk+EcWMPsYga+7311ccZyd6ho6a/m3OLfY3rDxpXOfFk
E5bvWABv5v892PZV2Zi+jWWsqRSUfTTPMZwNby5Q2t2Sb7VVXaH8jrbtwb95rcHcJPBedmajhLkU
+0+gDlFfKiqyaFxlwJfOfsj16oAhNU0LG+c6ls8wFDpVCe7rQMnw/Zv80KPDFKRfIh/Kyw4orhgY
I1GxTPb0CX3qqraOfMt+WkT4cS+Zu2VhJ4DOh27wPgjGQwTjhILYjBPmo0jdCLluLP6PxCUw1f9V
n4KwIDyuM1V7h9niW3355lXzBzN9yki3Te2qvlv88qraBO4uis3jz8evRhscPouFNxr9XPHAHDXq
lQOscI2j+g9LrENlZR3Pxf0n5og17QKTgtseM40VYkjECVDFRmVN1cHBwEjDImcDGtifwnnSpPKC
nXT09PMMgWFaag8j9QtsH3GLo3/xlqIC1sdHmL7KvD1u+mnk9Anxg0tIkGrXK1l8PSkQDYWaqnUO
y4p+/umIjvjY1rAq02Rz/SfCL9ohFBWb7xRqaF/wSpf3PBMGeBps5pCGDmyagDjEJ9D4cFIIbkkb
W54DWZkVa+4TPoVuwYNcCS3PyNR4iphx0d0mmX+Y02TeUOc+9zNljNRozGpnZNBzS5a44BUhbhkB
dMgdeRMkQLlRYIhBPxS5TgtBxkjjnnrqsjhzzXEcDG0EC47i74ClgEBkNEh5RQqt6DfIVKKnZttd
WeJdd7kpYDZsZA1Nd2pDydRrnJHp/rpRhr+FID/VEuABFQmWwmTAlgN+SpD55rYCjWyXvI++bbLZ
Wcn6DY3gHgbSRxz6DtcS3D+iN/pFA0U7CIzFnTJPlTONMVwppp37fbDbFn6Hw/7XxXvuENv4zOJp
LUfleAxdCUoG6TrJxqKtQMk3/sBFJBAX1tw48bhEJHQgk9MrIpu4iqYcmf6onom45GvBwl2VMhf+
xefsLPiyuYfautYm2sMQ9jPMDgw7AT4rsbKcht00H2fICPAXKROkcK/ODG9qW17S5x8S5p4LwKoB
qZuar6OGrUKAF21mPdvxxhTYMiwMKYsWjctoZX4tAzpz+ByQVm8Ztz9hcyTmmvz1weNklg+KC2Dh
x7SPooIKFlAbNOekSXR+f+jAY9MeVxN3SBWzfw1y6dERvAWdypDLycVlE3p8t8YPb5H+fW89a5CR
5t8cYMmZrEOA7yqrhPqa/MUmbBbXur8atTq/qX13CQHl2H+VIl639niYj/Asky4jNjqeSLxsRkqg
el1S+0Vyta2tYQ1SCwUvD+dxf7DtfC37iFL6t8QtLaErpW6STahsGTj/jiv6SRhDq3ffvPVpq0fe
GDax0N4n/6NJVd7eCr/Zj2kxSfbus5jV8JaI9OW/b73tmIcLSiEEeKRa0XdRf18TeaExH9kNO0X9
78VtghxKuF4wEvdfb4oeYyUDWCOVoKnrCPZHmjA0GxkwxMDyMeUv04Coc78jrJxWT2ZqbXaTaCne
uBHKfjp9gH2OJ5zXrYAozIzd44grfLd8IFTu7yP4LhrqSkXii+hfiPMBOu6QEoLxCg/ihU6bpYyT
u7hAop8U87lDQhKvOZnJjd/eUdWnqQ6tn+oIxR0Mff5PgNjXiFCSK2o0/8V9WnALOFGw58Ikhx+Y
V22uPngF5mq7HaUIMZR/P8tKrHtXnjPsVBnysjARt6hEWios3SfmW5A4sym15Eawzk9NL9EHO+hY
HJ0kF2Ux8VuPapOXLbTBPP9dL0Eu8dHE/W8Ak82wJ/p/V4JuSCmJRVuwn6Vnl/IZuAVRmJJ9s9db
pCqH5pLSAR/a7X0oMjIaQNYGwG0bZ+umZOX5+VXQPhGn7Z9lgN7+6ZiHynSPc3GZF7VDZ7o+VCYz
1cDz5M/QzAZb86KQf3QflN8bsY8dOR5YLogcUo4NMAQEirBaWYD8MV1OD60J+PRl40nOjWB96Ncb
6xGgUfepFKfdhrZO9LblWLIR+1KVpPRLcIMf1+5t3lKxm2stucVhTIAOq5a1IfKpLbgPeNlBaI01
4mT0sSDvGVRDi1fSr08IPMVTW8KFB8I8Ma3Q7S4kREohtyFlplXeQQnxggY27nXMSU/ZcIFLmaXh
iqnBFiDXxgskcm67JGJN9LBjEyLB8yZoY07G5Uy4Dm3a2Fsw07DjaAJDdU24dQiVMqGu3JLjNcDd
T6C5JezycYLuPRO8yFgpIeU3qr7jA/eoDbZo+NRjY26Ca8v0NtVGMDMUuxrs+Cmtb92RXvIBOMnb
g0btv5/wYEDWzTW/zi/xmmS/EgaKl3Mbxk6L5MK/GM8ZRRzYLAlRTCbDsEfnvRsDBdO32mV5aSri
3mU1qKslGr4TZLi2qDdNNOgHRiec1hBsFfFp26zi4DujxYq1ihB7G1eHi/+doHJJnuMt928sLsY/
2bfCUQVU1kXevHkZxF27353AX9NPdep/i26Jc1jh9u4ZmcYvm7wjGw45G0dxUQjJcvKC6g8WFHw+
7YETFfkP8iWoIU+PpVHlRK33HyN4yXqZWWwU04jqqxX8rG/XAeoDZKjK2W+eOnSCPqU7jdj55wqN
U4Tf2mdSqoWmEIvmZjre9fUJIsEmwTqHrGLvCDOvwgKudvPpCFtFDHOqqM17czn6cNesmipZZklo
QuqGp+Gtt6Hs4FJImcRcLSMQhsd2IisRP3Wo1I8du3ELChBvrwny9JPxE3vfCPlAWdPBlkpObvil
5t9vr7Vu7B/q8cXJnIDVFabHtBY2INIxtJL+qIewnx37uoeqyLQcAhytvbk0IzvvQzVBvdjjc/Vy
JaNnGWgZthEkhhARBXHNadxBIABAKuFaNrhG0uzEVPB/Ce1nKRUwMzErkYwEWcA9k29cfFDaH/nw
oIIaA7doNhBv630lHV5Ie7JhikK/mTml/tZxtAb1+Ix5FbFVyavO1NelW8N+AQ/kpNfF2SrHr2UU
/4SJYDO3hunrr1HX+cstwvx93070bIO84vEcARFeenOm+TARbJMeC3PPahXMNfu+2cgxiFkKtVgt
wAUdka/n4ExOfkrAf9n2BQ4rtvH7oeeS3rbJ50CElQKQx1XwSKnm7raRR1CYhJ12exH/2TbFd+8/
6z1g+YGL73q8aJu9ZD9ukpUJqyzf9pt5AMRip8PVy2aeUWDNXbdG9d7gEWIkX2BcuMntUqIL13bg
vPQ3ihMsNCNwIvAEdz/x7ok2MT6ST8qH/tFtZiQYIgLh61MtEp6RqVCiZOxxmCk/BmT16mdeUQyp
VtZwEUzMx3964nhYrwVjuf8iLXsjyKS9FSWZCmPJFiT+u3Iq5sspeiBwMucAntZ+GHOYs/gdeuQY
yzC2I8LTzApe7omTkYpol+XHqcLl7O+iwuG0goGR6QUcpY2ZTdbru41heGfh6TWMAFoWI573TIRW
4f/R8mwm+yPew/L4/PwtClEdxnBvXJMC/8mElzqnLfvlhzV/FQiBeBpxgvL5fTG/Ci+f3lG7s/KF
Zw+Oltv0Aqckf3rwErAlZfwDpWspyK0T1l3BIN7FlrIM4k9EtDPMSbPvT4rgGEkKySXJWgq1ZrPk
EwwrJZ3Dr+WzEJcZIQnvxRulV70Iw0LUdwKJyrHslFI3xOoB+AmOwHYoSfjDVvHSsVjI5XCNonf2
x16tm6Zxlhij78uNxoBHDlKGoz/LK3A9XYCxaWCO/KQEtcEFgkb8GJDtuMt3cufW6eQFzdMFK++8
36uME7M+mpcfFyKHVeMbnnQtVPai5hditxFxumCXWgMV5G5j8Eqw2G21kOL+VWghp7t9XA1Nl85F
KCkX5yhMkuzOkSM8PwVnSHWSYvPkxDkp+Ka49e0tPDbz97ak5IwiD09HfwKwF30rFfp9NMDfPzOn
3ld+5JKND3G1kmt7WBYCCx3tsGTlh3EJZHkgpKS8IOuLxxUsGdrZ6dSs6hVin3xYSzZdveoAX+JA
VExmAH7B9+SVy7JUydi5qsI0u00ZBnzdv/g0UVild/i0aKZrV1qoRWADirxgOjID6MaVRqZMqFjw
X1YHca1yg4TN5E9KRzdouCg3Jtl7+JKyufGMdCdXw9UWrtEE7TuQyj2BuGadY8PIQ9XJTZb0oIoe
Db/Tdbyr6mgwvDOhL1OyeqddruUIj9BTpCE1yMQ8yP7Mm1OpWqIA2gXQ5HZ78uJ6DZtZedXhw1ne
dYZPVVbeKRFvc9dN9exfoGuGiIzJS0+uhdN//Q9+dyqaSkcFxU3dtf966epEr72MOX85Kl1FVchS
rOsVUl0MBtBm26ZaicqHLCpTEhL8eeQlpm+FSPhXq1lPHHvtIVU4dmeEbCB2bZRU90bGMBcbtp4R
n20v7IqbphPR985tiPkafenSSw1PcC4r2ssmdUS7xuBc2/bPYxt/1kWS1D5KeG96A3MUZL+IDsvW
I+Ixz/8bnnNupN8vdbuiqHb5YRxi0Kto/NhvZnLVezjsKR8PT/qtW/lXzwUZiriU5lCGtxO2E6em
0B1uT7jHMz6JvS3KNr7CKeAmSUmgVKbg3o/ZES/kafkzKxDpl65eAjrJWk7ZKw2awQTn5qGKfB2A
EsaKFZdWqWwLorBK4dioDdbVB5YqboosBQ/7aJqohuU2VthxWRDgSXqUP0+RCYl35EYYCjS3IIH+
Jv6VpCLYKYCBc3acceQOfBa8pZuyuwIwk2n5IyWgwutCH4ojgItzGE4prglZLfknPV/VEFhOVVcH
YM7vOx2+U+9zBXOGihHkeVp0BFbMrJyFNv6xAxoMOCLGh6/DKzxxVInmeO9UR+pyV0SO6CiNwyrb
2bw/L0BvnoR3UiATqxFUbRtzB32w+vERgqZyRaW4tPqWxMudYODAUKUy8r+nFJAghUoVwgYt8kaE
XayD5IwOt5G0JF2F7hsUY61d6EtdiEZw7k70r/Cki6eh88OFjsXoHI0lOf0AkAt2faktbR42nTWl
yKqQvBFeCLgGFjF5sm/K8wN3e2Hn+9+QD2EUrjQVIXiucW7J5Wqdktj5EgG/3a8m+nJ+zdArTSXB
Biui6s8aT1hsXThQGoDQNrAJGD5EoE180RESecnJryWjNZKmpusULcErc9Ki2pnZZXIz5Agav+nK
rcNaKMFFYbDAkjHxoQCKj81l3/1sVcaPgQpdKd0X8s7rdOJJogmdNh4c3t+rcvtYis1+BWorgvd+
ee6ky7p4gqVMNpw11kLrWlrPtCDB8F3KlHZX0qCkXwG0sseeN+kLxsD9hzf44Fsn/OD69Q7J7wUO
6CR+iLZPmm4z4TpzzKRGP4dtPMU7qk6XXh+UAR9ByP2h02k8KNV1rqHlM0P2AgrA14D6ZmEBjszm
l2zSBFsKSgfHfEXrzqMlX96DEgQ8Po96Vf9Ps/EW73EW31zqJcEMh/uTdtqKaiDw3fDjH3yM3aeA
X71SpGLxBRIzxuG8WK8bnopNcPKGQO9HJ+roFD9sLM9It8V6HTjBr1j/BZmv82aQfUnkD9X0FQiR
1kRaLW3odXzHc/udcZPvqxZHwjbAagrnHhy7E6JGY4cKz7W9KrAj62xTpLGVuOwEO1u/C/JGejI3
tgrXGAnVHj8VPYb/Fuw5d0e4mkW7Mmx5f9NOTcLZgA5DTKdDvI5GZaY3+0KICg1r7UUUDi4/Z2mv
INZC0Xv9y/0AZCZC4AUQm/qZk2nxJOd7GJ/wbBuCMYsry7RMMu17EsZ+b/jDdBRZR4jahrrXcksS
ut2NMjMRv1jnWxJyIzQ3iQwm3I/7hmN6tyY+dYF95f3Mo+8Ii0xqLb7mdIZy793CAB58NoSo3rge
FZyXYcgRV7yKboFpWkPaxCh2AGimX0+r1FuABTkaHGwEhVZzEUw5YywfeB5H0RMjZxAkCj18GTua
JtY1fq2Z0ars0KzE4IzWrIub/1EQRugRkLOqGTE6bUUogmmLdhODEPJ53/UYLCA2bzxl1XjVmRhr
o48ecpDy1yxyy3odQftaQ0BG2sSIHAp9cmQLhQRXCn/neYJLmpNFWFnePsFf3haU6RDGGME/sofd
bQSgnN4tuPFonvC8cwicUwOQIpRcO5+79kXOsak5eehJl2ZkOiLhNBUkE6toufEJX5I2YXzSGM5Z
G6Vw57NWbL3UISWjra94P3KrIiNvVyo/XqL/8ZCe8eu7zlNEjS+Jb/uZaq1KDxmRO1uY5u1/GHjf
7lY+2/l9/82sAjvqv0DjzDHD/43LYdMtzKvU1nCL898kXDBajsJqszkaoRshuJv5UWtH+tF2BPLy
TuKT2gY5f9jCVFy0DP1ic8VU/iNBApSUyvhzL8Tojg++pQNPZegbM2BNObYmwl+bgHjEee8/ABug
EvEhmgude6PGhOVIyDwC+zgVINlnX/Ys7SwJ6xk1JaZSYuv5Aya1+Tn9PJiYpd4i3Yzew2HgZ9NH
h6/+Ccd3LfIYzn5JISICSSemPjeZFk35Z+rxyWMhVgvQsnzPA9gnzDf8APCuOAVbWxwaWxfgjcQr
X/GBTPhV7MU9dYrCIxbUUPv3/j4SnIFr2uU4fu0EttIyRUIJ3pbZrS+V9KpGUbn1AOiiOXpF2QnU
3hfmojkUl1391ge7FinUDdhR6j35U2ijwFNtelTy08S1KVf0sxBTkuPWRErRSXyzWvGUy2QPb3Uc
+DS8xn/cP+BBxfmfe8FU4+w/bMgzW2Imx3s3JMilgtpohKaXYkUbYNBcWbZkH0ABdxB1AGNmSbrO
Qi7eWRc/rI0wcrUlASLAYZIpwSZ7giYDjGMiumRl1aJDzU9JTJIdTvu52fIRaDyGghmYDc2aX1+C
KFf2L6GT5/OjsL8glp38Nbh7It0J9Xc7VGl22G7lK0God2TFfzs4+iUWjemeddInzvU6oQbREd8O
UAc7tWHgJs+CdvnJXFFmvFnZ9+V8DteI6DasApiBKie1C2Ivet5UK2IoiRenVGgn29jNCzGqkDb6
Pu6AUPUl/nt7OM+9kxUdFHctAGORxR0uLFhUy/5EmgbWQo5rgAJLfqAciVWIBchxEv+dhlaDRCDR
j80j3Yf459dqDhowbET3mXO28wQM2RutgFJacucXJEs+8CUu4qdj3CwzUbmnV08F5i/gZTFx7ixL
OBQ9R8vzK/x31G6W4BBhpfqS+cEo70cHl/al/aVkaZGk5kcGCMFTjg5SLtoIIHiTkW0Gv+hndxP7
Ynn/Wn8l7pYkB2ZYNOsKHaOKqWaKlspeENQ4rEzq68lCI8bu2pW5dTlDHQt3OCWeA7ZHfG6+071v
YAalbROBtKOVIVWinyvZj+Th9mnkqadDC/yVBbZHzFCtycxutoh+mvhedxPAcYltEAhel7ODJDwm
YRuSNIRk0V8gBstbJurZdze6pzGr/Mgafhn0QidRB812bLGwKSoyKPjqNLeyBP397oX/rrEohbZJ
ubU3cR3tXSBxmDJ1lTuKaxmuyh/2BEd/uv1kFFd9k4DXm7ahCJRxfBKXgtA6UAg1vkcCkRJ4RNVB
2lIvyP5DE6f44c93rclfnAjuj2ont+cj2/saentKngx8Qr1aiZa4huYtJPQGRVdXtQw/iQg3AOmq
k/vgkAyVGvKFaJm2aayNEIr+M0AuUk4H7f4KonPgV4u9SHMEWJb12yGh8Q71L8CbzQmz81xsFtSR
ofN487OI30cwXh6vRSFlPy31oiwwnZLwrZmvVYx4574+lMcXcuBIHdeWdgoNnedH+QK22Gamzz+S
7vFdHN0mBz2Z6iwP5DWveqpI1TEzuRd3jGQaj4PNq+5L47G+CBvKclOVRd7pMTN7G0PW4Y0avMTS
MQSG74MgK2Ril5oydecz047PZNyhJIp86YdbISDcrhAQ+QYFqZG8goDOh/gb4xWpB4tgVLlmsj2c
WilGZY2YYysn4GF6y4nJJVWOxjLjClgJQvZeGMAEKVRly8IUHWs8F573T9zqKocwmoR5g74jqnTq
uz22KVwjeLgUjx21wDTkH/VvY2DjWSbPQh2IPIQOqC0muemRiAl8DhpWb84MRqq1iD0YdWvNqzly
H9ZV7Pg9zK/EpVCWEylZrzS8KRQ+e5fPQ2SK1vDaT1dFcfiFi+Kf1J8AUVFfnIpcGMHX/0VwH5Qg
Qqqhi0qy3X2XdKqYjquIMNPKMNBR9X8VFf0PVb2W0yYD8yiT8lC5fFn0pPpd51xiYaSiOclYZiyG
uAaLfNOR4zLYZ48ZqyeJO4HMNyWirQBH746kLXXbCIjTO5+GCTwoUAZnSpvOp5++6qMRzihTicH1
5iLErfRUf+N9ievt/rxKDz8lspcX1jzRM+ZT7BSL57nqXo6JTsKXtaaTa6frwJTA0Haep8dXMqDm
fNKhkNLFR4gV63ugofROCzLLut3GQ6Y5dEsMvdr6Z5AAHWpqI+CU9gM+48QtRVZdeqPyAnd1kSpb
05FssM+93vbHYK1kfWUzB0OGrc1fpRkHD4vUqXeJUlxdInuYqIAztJ+bVC0EOj/naFv3WlltbBoW
PpUMj+j/Yt4O9doeaOn57S3anfBOPPt7PzXUr3L0gcFG1TqKdqginn2G7MPFqeKQw++rGY5yFi6G
Fkpf4X996lqjxPKjspdR1MtmcZA8zaYiQ8AJX30B2Q9GIVlxCpGRhyWfp5nNjV1MKVmY7HUz9N1o
DemUGVG1Xeemr9VSgmnRbRjQat6jA/KHojj0PMlZQ1MlWumOWhQUxHKYEGFoMCJvaiTb03x7AiqP
Xg8l0wiXNznhQrF1W+F7aSdEj8o/Z3uXkfZfgWBQ8Fewn4xWWHcV/3UNQeXb+oujv63PAwLXpMGo
xol7KZc7SHVr6ALHQWLhFD3ZAQCHWDvOyzBdkWMUDCViDw9HLtA0oEXx/jTXUyAuNGCqTP0/LZz+
rhP6tY/QSnSX6EVxlSP4G4kVSrWbuZ44jpzoF+xpYVc8Q8Xrm4d8UWI7Tsc9NTs5wjNDVDHYG7F7
NDJZqFG9sXPNSuNzhvngaKcLVdiHi4s+WEtFTCaRRMVoMgpA6Dn805gR4Csc5tZtBeGZ//9/FjHE
D/VZ3vV4iTe6SZC1kkJnJAcTbsD/wzvFr/I39W69XbfYvnxHaFqyZc0GMP8YPQoycocL9p0Mv5pE
KzkuQ4ipkiV28Y+BnWCsFzfwKKvGtd3djoAhgUtk+RlMUAdmZf3NUjhO+XjaQu4BpQw5lrqBf81G
mYVoaGJyu+0/HivFMf6Q+NyERfxUIIUhGEpDT4DcyHnHkRbMUQYQm1WM8nf57KKvuObPFf7x0teC
fwdGfCMUiF3iqdzMS8+2efy2NF5ftI6BHEH5DOzttxPlDi3EAm5AFq24Eoyy54iYDnhhmt28ri+E
VR2jDmCf+D8yB+5yOsbQ0bXHKWxxptYs/DW7DJ/DSgPj7Z6Ql6o27iOMRAJ8dRnt543u+9B8+S8b
zGcxa2GIU/c43jdFyYJpRynIVCK+jZQBu6DbjNOD8ez8K6IWHF2TZIZwYC6VZgVYCbszS98z/Y5R
I9SRtad7CCqgbjnb5nM2wBgayLy0rVQGuPPvdCXvVinA4gGft+7gR29uCAhvcsBqmL5nz5+q7HmK
Yl7vTmcd2moBNKRBiKyrTpqpFbCooFxODhAJ+kIdG8ipr2jYE0gNRYErJdTLY0BQ3T8EZ5d9REoe
UUicSsNgtyF7S5JHEhZ3T8ZPC8t+0ORVqwfsgpFdA0Vh5X53a63J0lHiXdHavEKTtzx6rnhVxYag
9dwxpu2K69Qc2IYUmQB16VX2NOGJyRNPyqhbL+IhSfEoQgkb78cwSBgjE2IvQssaGm+tZcgXW93S
1iACyOJHgefn9pze2GLCXn1pAIyFYqVq8/ImwM3++QV2Md9cuKph0hYEbOTjasbNeBfukfsnvsQv
pAesAQeJdT9PAgqgwfsPKpkicOukkk8v+RlM+IMza76/cu/vxWaTbB28fnHOa8NgkZfhM34q0j19
BWAZ8T0cvFM0QmyKADT+7jIgqyBRlsm2WIBBeAOx3d49Hue9H78QJFLTXUcSpOhNilgKnWF6EIRr
X7wyX+RYBM7iKHniWRN8VQNAZOzqJrdK2Uxr/JZfeyamJFbpkRymsTH3yh1HjMMroaboEjyPAdOc
JU4kxOrJMKTeMiZ0QZoUKQXlOcAub2aCl3I/QpC1Nt1IFYqLn5WY9u7rbqJAbq+wu0W0y2yTBpWy
d5F6OgqHh3Fw4KMpyYqnchw+/x0znURfBfmePBmq+3PU1h2oKuUzv7q/rQE7uHGVGj3uHpyNCC0v
9t0nHH3cP5sMSrqit1+7a4IRk7jYO3RymIJVn+rei+NZ9slKyMTyuGIMJ2f9kxWS+vq8vCY5EGUx
HA+XapLoziy3nzJm02OGaQdBjBO7pG06xhuavPf4bAIB0UsY3anV9CrdZHELaDqysH7p3sYkj16/
WGWuJj+/WqoeV7rOo/yxWtGIvIX7m4pbX7Vfzp+2Zu5ZepFc1B4PF5tSHVGf2EwdvLbWKT9YOLRT
EFxPDhnu0ZfBQzPL96ZvQWH+BuftMgdY9MvSE1AqombcrVsSA7HHhGQh7L6Mo73YiJ+ZYuFlSfMg
05TzYM334KDJpQBGUfV4McrJO9oUEWMD6EB7GICYWTw3SBYgYjAolBy5WVccJIYJhIUaekV0D4q7
voUaBa2V1EUqpZq3IRNNNz/zENeJAGDXs+1SK/9C/dM0dyPAvnMplSNFGbtLSjLeUNYEw2Rt5Rn8
qnM5XoQjQ2rM3YFlFH814b59JgjnCEUmCsx+RPsMSTbKswLDw0mByCDVuh9BXvtFfUoAT3EF/JOR
rijzVDpfv6betdBWCuPJjC/X4ytukJykfySnrAH7d3eop8jXAu3/Ut8giJwmpZFzR9LSvgfdOUov
+fw0iOG3mT66hqWwqbNOMqUug7i8d5EOkaoDEH1Ft7NcP4kEqx/7F8hD5EM8LCqX0Y2WvunAck+6
bZczOSOU4NOH+GP8psTv6V1NblpeswrYCD/YJDdrE7so2X12c/zTHgOb4On34AOa6bbi61kL/cs5
mh1b2zlXf5EVLJIF9NDBE2R7IGf7K7Looe4Yuqdf/6c7crijyT8nCKhqrMpcuT3roeYDSMqSNbqn
CsqGoB3C/DYYLzXiGEEVu/68y/MHkgIKvL5F09epIw/BEU7EVTVoYWp2yT0D1URTdmMZGFiMq+3Q
FqA2etqaIgy5Kq/mWd2mqjaP7TeseG0iS5l9rDLIEhsb1uqYooMSTto3J5IAxZjOTRdFR9RlSsWC
68mTjZLl0RkrGxi/v9Azewhzr5jNW4Phy5hVIcx5D7NsPWnUxD+6MSqU8Ufy1XLhBEh4t5HptJAU
djvRpdYRzMxsI97sz7M9XmxDWicADmSaaoZ7aG1Inh16os+1zdNXwn9X3/m0OmoCG4GZk0rtZwHJ
Oy+8ha8UuT8QhqCY72GEGFTI5O0SB8amBAVFAfMYVMiRMnrqFFE6aHvO6V0PSPaFvcPdov7z5yCs
Kao98KX8uLkDaGEBB/zxsxUNcstnK7/Qp+LkE92rc6ZoFru1IOCfP7Kei9i6qKLPT3ha41rnJkiX
IS6rmiAaKxx3vmjQmbPDc0AjCprCxXpV/7DFtWZNSweCiMJMqCWAXRUThxCRqg5Hm22kP9KOJBXV
A4iDAChVfsnpWiInw9VxVVta13Hb4jxlKqPs6H+OQmuwhTRSF6bFofYkQGErMu0qISeULzPnyx9k
WRTaqp4CNT1z4WQLgf2GJ+JS56T4HdPkAAEstu+iZAAEskjqZe0wWlrBUz5PSFNGONkKwh7C+LYC
eY5UfxRO4dScDKgVJ+Z7X7eEupqLa2lfIAejM5SBmFHlpH1nbiG7zrKcw5cGdwNZlYRzTwLjNuMB
xddnsiAQlz7YhzFBPdU4BkSnLbUD7I+uCnOtkSA5ygvD/Fmavf2ooYnSVACeaB/1Dczhi63KsfkW
7dcZYz/HSh8rNP4FeaViyx/IfMeqvxs8jdGy+M8s6QpCi16cJQVFrxx6w2GsrPaMImS9W3OpKyRJ
4u6W1VMIVHnyJv3c9a27WY2hGiZ3qPjoADGY6uoa/cIyg2BfL1UJQOgEMYEbA7X13/37gSa3ZrSZ
L06x9lqhE7jyAyE3jbBaCGWp1WPRYYBNHHT90wpJ0D1YKFek/M39lWUykd1Dx3KwAVXJy65rKlCS
zrSObxudlaWuTasw4d2vOOsZbRTKNOWvD8yMej9Lye/W3mrwnUXYGnh7k7q+7+2ZTywNoTZMTJFC
v3pC03LmfN1KCAmfS9mJZnigm4NkVuitgMnQ68T+pdlNr4X0sHfwcTcNTdMJ2t03cNgUnFdCJhet
WrooHiFzZW067Act/CxyvNPn7KAkuQjz0WJezquyu/AqFFkMHni8EWPYoKaUZD/S9OI6iy9Dw4fq
3N73W1vJB1rjv1ACUI88l9eqsL6Mu3Sz7tu8N7UjdIJhU3TlYi/7KzVjkYH/SzSV6n+4IuhnRyv2
O06xKsAj4/W8ZwRChtV3Cr2GshDMJMCCOGAyXS4hQsIwKtHZqKqwRKtRwavRKgFET9sBy6wd9u8H
y+uuCEnSYxQ7Wx7lA3M6mZQBkrwWPEhcN/TBxC139J8fG4F+EZmGPxl1DLc6hV9tGoVN26RbDdDF
F7TyzHif/f0fyOuuMErS/v/XIZprJb7RxKT11L/XJ2SLjiOUlkWzzqYlr6a4KvfLolvooTfrtgb1
WoU2nr3zS9jD9iPCBnDoe8tvl7+9tZJHnbRG2G43NwT3QfTvp16nxjf6VO4IaFxzzOHRBRAOocw6
9xpHMA1d6YHTLERNBEOveYtJE5MLUPJYqcPOIQW+0Xic/eePOnEJZEgWQu2JVV3ZCEFVI5aNOAAw
95DEmtaLoaZ4XqlO+RHEP8o3M+sGAIQ3PFFqHu0An4nblv5Ttwuadejc6hesg0xMvAs/Pf9a/0BB
C1b5M17Hm/Pkov+fZurI9JtlSqyzEuQd26rbT79ynrEdpO5HRsChNo5nXP1y6BBAavoxy2qrIMt3
rq/a3rS+yZzb1AflapLvMosWZp5PyRs5zKLcAX6A01QRuZR15b4rnWglIY2lxMPcYCVqGzGpT1VF
TaipyCbYPbjvgdASC5CqzyBN3qFDP6EA2gJtl/JuA2JS7A4k77PhzMe/CCqOch7gAVoUR7F2r+VY
16pFCZtD9zCkwOk+vXZnCprK0jbKWALsESpVvqUsGQJgyA/Q0okrMHPWDr2viY3WtUdft3Vxtl0n
MAugR2oljN6kBkzrq9bQSeEWNN+xvtPGqsoYzceG+55tKPhhVFHfb2v2c3dPN7yUOlTp9hC8tvl0
X5po3zLzS1Bp6i5/7Ax39Vj1v9pf3SJYQVTwOynCLSO6TBEe4Ytfrz6lwCwRRuGq0k+YbZvmEstd
5t0fJtfgKOZkohyAJpHLkwHhfJmo76nIlCYfhbBswXMnfHCkGARxz0U7SMdBirq7bFvllkjgGv/G
xzUcdbTNf5BFB4ryuMDghPdoFh/6itjDIktrnJyPhstBlC8IFHoLRUiED2Eu0FXE/NYIp3GJ/K47
IAU1W8kCkgUF/unYB5a0bN4JBlFIlq2sddaNEm56f4vEMQ5LtWMF1S4/VB6U8U5XAahHIeCZAVqR
BeBQ79pMrqencpTnEhFhDCFALqrL4cyIkvaM9YnngEHsC0AQVPsxfi4QC6kRwcc2KeUqpI0fDyp+
rvsyiA7vhUAwNqgJKzpZNCHuW8d0jMNu4nzzCQ7qfZ4C3o+2jbbZSSrwEDsV4r5XYVfareTgvXLw
gT1Gc2Knit2UhlP8r2C4ZcPvhuLe/wG3GIs7zl6dUydzO1tSOo9uWUeiHkjJgBb4AMeAbjkmi7y6
dS+HChJ+X864hGnW8GSdI8DMztnyLefX607qonAn91RCwoPi8EbGNfGuDG/s5w1HlSzvrSRBr6Z0
DXj8eqW1youRhik0/5e50WtmteWibYr5uPCb/OLjbJtxhKtFwAzG9K0888MgWrZIedk+5HlKBr1f
aS6mfZdHwBuwpOOukP/u8nEvQoeMii+fcjhwXIaW/b0Kp26wubLYfFdXx3qkuJhuRiO+Lle6rL3H
QUTO634E1micDuNqdjBA0g5U86PuLCWx2rqplTgmfl0vSPJnfizYUUaGx+S+w02kBDDCLRzSqpma
zTO8PRp+KKOhd7s+Kg7BG58s1xfW3TrMVAj8CZTBBRkvLlGh/3v5Dp+jawYPODBU97z7nctUIwj1
W9s2w0oH2I7XAuRFkNZG8N6/2MrnygoEpJl5Lag1aAwkQfLZ1FEGAKGrwD73oHWh57zOgzS18Lq1
nvUff3VOtm4CYCZaf/sMmQ9atG8MLBudOjPVmXETkZW1EB0u1/hZJITVLpzDTCzlDD355DLFiWtG
DDf2QoFL4Jvog1k/zVX6nBdncoDQ8wmr5yn0OV6zOYbvK7XR5CNyFczaT4hr7DndxA/dtB3CPZjb
iL7+BtsRD951bMIfn/nxIlV18a/2C8eq0RJnyMyB/wKfVOMu7dKR8I3sOolgVs/4qUEqS1hK4na8
cvEh6gXy6v7zDBSiuq3xKRPHH6EOH6/jmYo5GKetuYTnY/o+/82GL0AXV924cTJAQOkueFpHzwIp
HYjDF/ZcYJROPfWl2IWTfmzNIzuzthrUCw3W92nUwgjD/I9x4Jg6vMp2oGNNkF6IWXIHb+fRFrSP
KbazBcQ+O4zDPAP42EP1nyL//soC+IMXHAFEJDDkLCczv9ahmScN4Kjn49Nk5Up8SssEcAID+FVK
33Gb3PA0MDElcKvuBoPb2vgiPiEn+zY+X0eeOwpIfMF+IZXrUIlyhHWmLDWtxAPnnuCkDfbkd5wf
kv0bu2uq3bVi518GaWjWss4PjvNvzO8vT8bN0zW45MjTGxr0utGlAhJGo9V5Y73PIiOU2asApayx
CRwLftH99aeAQpqE3abR9D3r7CYSlDAhY/dAtN2opqyAxXJTMk881cz87LSdgtmOhEiwqiI1Ua6j
hNOFezzjYvMba4PNrvaEAXbGQoD9j4NmetyEXsLOR4DkCYpF5hVFlfwqtcFS05by4hCcwRhWDzau
1tqb/4SkTVve37ybeKq9jOoVPF1WMJkLxx1TY6ZtXKMAS2u5mZm27TQTzE46hEuhPrOc3nfNDBdp
TMdNw8WajZT9BpOg1Vwfgc263joC6KeEbxjKk/hIoZhsN3bZCrDwulUZut3s3Akewij25SWlIX4J
87i9GCt0voBFQgbd3PLM2rLMaCi8rGt8anfPEQNdWORXVySqExjgBjgYqK7IEltYfXGwyUo8Kic+
a9D0zXl1wuSvg4pweKsu4f1x7wd+kXt7ptjcMWVlbswOYMr74EKZiyydhOL450cNgxqUbf/ASvot
vGtNmzoIWRUPegbLYomdtFQ6H23ToxHobph8bGsy/BN0Gda9wjXHlka+TthQsRBWcuMjlXQtyAih
X0I/5NloOFO0Bm5DmArDRnnpuBqJCZ0K3hTGK9S1yDP2lad0XWtceMW8nCBqEtTKnlIfx2NmvK7H
gXNSJZYcP8w5XghWRFOvA3j7WZGj19txoAindDR2PCX22vVcS6iMeWtu36aViZ+z+sb35z83XAhE
3/anJgZTyhjaT1rhtEviSEAXPWlUd21thakA5gu4ZUN87L+Yy4UPBc5w1bj95OE83js+U485EVWl
syPfdMObqxgHE6LARQGWtV+tBY9QrcIGsnI959tlG5Sof6AvOh2S/AmPjJ/CAYyJO6h+p5JovFaK
KGxC6XntLSjU2zUEbD3FYqBZBu3li19q8k/BIHzw1j5RE27BascXLIZyup48wHBWThuYgH/sLTF6
6ZktehVbA6y38D/JOhKNyk6oE680/IhURVQMQiJuPhySKdqMorM1y14lUu0pw6R5bfi2vZpJ8JN6
6Bq960aO12Ta+/soXU95FUs6awEUmz0yizauXV+YInxrqcfyzTb9r7UW5zXhwuRhqi9/Ve0+deug
FY0YuRg4+5A9q47aBg8+6mLzDi6bmurYfAJMQhLljzcc8qAusTYCoWSkB9BVTX+JkR9U16qyzbcS
bjy/CMEz6JX0QoU+42kyXTVAoUjFOhWZrS1ML/piOr3JiTjtLYnqF7mg3NQ7TnkuOWmqSZeekHY8
XXx2o3QbDsi4iMxkHIPd3jlpmrisWJNRZhuc/W/EKrXpGXiv6hnt+RxqshFk1rhxtIPYkOfkNCI7
khk3b1hyr5m8hatel/VW+VBLRLWXojilXFMAy2Z+9vLyUg06qCPgv3PW8d2KxuSDNwZR7tsiyqmI
Bhn1zqURZaaXbBtk5D/Yw5dsjTLTBCNkr0TnWyx0tT2muTqgqhA30cNBzS9YpRQ8ODgzSeAyg9m6
lhssXcEA4OUx1D1uKYsf7C1NkncOXSeHhvIkWdcS40eho+OgzdcfX8iF/9e0P1LtB5kAhSE5U9sD
OlDx55QFGM6d535aXnSG1YaojYWry+prbMXWIqR9z7dzGJzAQ/J+VsLqI73TnIBVzKpo4lHF7lNo
9rG/IfDze0KgNk+V/dNQfUBXA+XEuzckGpvZsEd3OVfX7zxc5Ws5vCiP0Pga/VX5OCYkC1WDD85q
UFCCnmO/1vRz0X0bhFE7k9pHr9hbLKlacrcJPSmopcsXQbLBYmeh7IDA1DhNPXinWBsg4w1FEFRx
KkURfyyZ+/BADa06amViN7pf/V5GMJesiCgTSR3KazcJlUMQJcqHf3KPJ6K1pAV6AcvGBsg3vdEB
NJgqACsN7HAUKv3c4XltEotYAtovhFkyGbV6qYgcx1mEuiL5f9VT6rCcy2yQEKuVY/D6F68gzj5j
2DWniPhSORfSzXbF1eLVrz/yda98duqzw+zBi+v+CO7rF3fYjgYDLvjOg3TKWzvxCe/UY/5QrJas
NOpyDBuj03JkWzdvVnqFovhTA3iQcHVoQ4whzQu+Il9kI6YAEYeIwCaH6izWjaB9ivwCXE+ywAfo
ikBkb/qqf9N+g8lK1uxhX+f+7h3ER2zwLtNZkwj2pW7ZJ66KZIdloVRT7N+eTeTmKLWu9pxcRvSU
+ctEa1QRITbRpe7hko9jl9P3Bb/PEvSQqSDdDezrC5Pn2v5ahqAZuLd4nRCJfvbiyo8gnrEn6OcK
k2Z8lkSzreUB3nPTbb3f2BnKhIMLU9qbPZkYDdKIkmXQP58EDEJVpauxfg4rR79mNToV5cNPAprT
PDcsKHGKOcqVzXd2dbcXhLzVXIwVZzhJ3tBIzQ51wDws00O9Va3WYQkzfnBOIOM0wgabTeAAoFCL
7ITS4EO3oupWZYXGISDVu6y0WO520VIpy+MgheG587JBHu3iedo/V6Mhh4UBZY/LVaMQlZA+agzV
DPxlB3a+OZ3Do+YaLmMBJbcpgtZb9V5fx9hmz0AUpeqCxune9cFYSriaXexTJc7TNMyRX2rhfSib
3R95zeFljFSGKGgPog0MApBafZJsLG5nJPw+OAWwSYqMXnL3rroT0CpuvkZLf5YWGUIfbu7iIYOu
dSupBRqACHGAz5DGNptz/OYDu5QB0g9ax/vnNktWm48DkpV8xo2L6fijZXwTSJgTaApdxaDp9Edp
pB+4OTjKARukIYc5Yv/rLX9YuRZhJt5uhRdcWfzQUeYHcmLapMaCKY7AsoeDg33D1IvfKAaPj0J+
lmsKMm0eg6/Z2PfIGUo14DUwJUS1khtxlx9tT97ZPEtUukWdzjVRJORi7e/uTmsEXzrl7xmULrfs
Iing3yI0u9dCg9B/BS1zD2YixMlTyZtsv2LYFKQOL5ep9Jlm2TWWeg123KrkgHST6RligpLJ6Wgu
L6KMU2/XKumOn69+ty5OchCK7vTPgjMe8/Dz9GKnVB9QAqANDEOMK2Idgb+EXKOTGz0OYfb5WfC1
2wJMjxrqQ04nyGTGeIpuJrj7XzelTgs8Yqt+vLVM7gmPVBnHIL4x/QXzk6fwXh+KmfCjHV21FsLW
FQSan2AQnVt3osikxYdUm11FDQuZ1GwKoWu8JeQrwjpUgtf+qXirW2Ftd4J0r8XFgjyHa/IPccs6
qs1qRGAq7jsHXja/bzYaN7m7+edONcS0gWHvGaYEZZ6mMCmfbJ9aX2ZTFWAXR9ymvQKRcND9Olf+
rLBT1mOMJxSrRZH3c6Pd8JSFGeGfsRSza8JruE3Ev975Dj6GcMA8+EnGrvfQq42pgsaCUjXKFKaU
9VSuuxxyBLmvhyRXuDbWgNUROnDxrNxtqmhIuSzYAl2PD9lzU/g/ydJiQRrhYJbjcxVhIWBZW6Il
GDUOdV5d1oOeJFWNgu1iqG8s/y6nUMb3kP6G4VtYwlbs608Fs0QZlD462mQwt9jV0dbVsDCmIph1
VGmXy/D+94njVX8Z6QVB5FGu6a24t5AAPzSB4kXdm4w29MbGLDJ+sD8LKJXgs3z4gREZhZY1VJZV
obgULF4/e3Uh0XaJjQNF0wocOHPF2lZ2WG9tX/h/4K7Mx5AzmOMX2ztoTo/wmsoPOmZB6egwdQ4Z
o/Up22tWx4QRRpLch7OL3TOUwkLLpNEm4ssxwLwOrQkWFCPInkFcswA2sSS6Y2uYNc8gd1hLBywT
dZOjczBCywEd+ofGAQJrvwAr7+n1w3vFqhDIrTegGFC9wMx+vUBTREiPEJjSjqWf07mnGftF6hVa
SqxnNgziYSP2EAduKmdmcWpiUzXBRj+Hj0+VFQOP0dehrBciVk2U4z2kNgGyGgK/iDLsDJce4uLC
WbU628f17wVQ7Rp6ooZVBAPUR5+WeoF7pZOPEv/+GcT4HY2zFLWhI4M36wc/MBNB6vErao8q+r2V
eWhjJsaHH1UW4qOOidtZCZX6ij/xkk8oFtigEw5/skUey1KjjgwQw1TpLi1NTeJfTOfQmUQYdJp7
i2hAXahWMGVRDtqnfonNzTTzYqc3eJOq6rO4LO4vXm2NasthhR15mJCSmG64fsUfMQg1Eq7oUAAF
+TmGqxXEeUE1pxH9N+fblSIFYu00ylZCzxeFdaYCD8a9pSSPrsoBI+2KCduwIkRRTMQSjqmJRv8I
WXk/GLZslNRbKfRzVTp7mFROwPiMGAzKNL19oP9wmuJk0Am9rI4s8J5m5jyUSfqBhPMU7VYHoJo9
6MognJvhrMQGCz2TLqJ5KtVtJTqY1iLGyCc4YJxvr9ok+2KdS70baYvZxa01ZDpD1KlrJXxH+Vin
S69V3Mnafn0yn/EeC/bcQTacbigIL3/jpz79CpKo6WkdtruZa1VJgIxRnW4WYEZDZ2KvN3dpwSps
IuiX7BYoKBgJj4BUuWnqdHav3re6PokvSsTjN5tdiWJkwbjWt6OSDWQXsB1h4tmTox4ck5fBot77
3GxRZaSq39v+RvDeKDrmnGFlqRWUQLrA6urqNhDSKxW4WORgaRX5l4GzubxhxkrtrAT7ZUNv7A04
poDR5SRpnuI/DJTgJU9bPcsLrvfcWDzjngosbyWZsCVYF7pSHhIYvzQMAxP18get9d4Y5R+4nLDV
E2KTHVARKobhr+E9RZnfwUQ21hii2MajEEWw9Lqlr/CxXbsOJy/+D7M6hYZmqapkZSWNDGvbVnix
4sxDNR5PJpdhx54aqKEJpgKF1vj7/Ts8apO6V8tHvGTc2FIQ7uLC97mtkAikqSmogRBb1Q3q3a+l
x79NZq1dSjJ/LTCXUIkh2uwIagomXbYHIaTmJ8EXji8+Pwta+KwHXTx171rZXLaLn5AbBYDW71eZ
M9xEu5lLbm55o6EA2X15B/WFQZ+ALH93kznTkSVpY0UWPGNy5EfhbN0XwkzDlRQNyPnajRrynjIB
5LCTfOWDs3DAzh+VmCTs3QBwKLU8fklH7dJ6UQcT8nWcLP6gJ2SyS19eFpYBjLsf9a4BOTWR54AP
4ATPj0zZ6xkEUIyK88+Np0kL22IAJyQyR8tH1MiSCemnY1cGPeTK3Nz0VV/EV0akWjd/LrhcORC8
WCOGBpvMif/57FZk71TqkEQSxsRqnkhWbUP2VLs7iNbBYlTHLIAXJ9G7oIMJy2OHlM2rYiIMDaha
dhjaT3gXrBvtFhCeXKzGGS0DtRBm0miDGPKCpFj3zW0sF/d0q1GoxbC+u+QsVT88CP/5jWQqAm6e
e72R5EHSCmn8kDB816WuIweHBED3gIWyqTsbix7nFegNI8q28VL6fA9k26nQ1yEOU6R8p/Y2teaC
rkFeQ2gJ1GMxOoU7bUvNfIpbt1ZLyjMF+4QpfptJltr4zdm/s4qljX5ttaa4FG3jWmxCgXkEvLcq
M77yO8mSrQI2ggsITZX8C5BLZVmoK0DAaf3HOcrTcZwU/yvWooWkirAspLHfKY8fbQ1SMfIaYhks
5OVktskjELW30yTtGm1qY7o4IzJACg4J35O3lniXFS7lTK0PAg5NjH/ZUeiiBJUmnOYW0F7sIC6Q
0SyqYMiFt46oXi3wOnO/rKEI4M0ZYsDcCsALAHcoH48L5er4YGhohbTUJOwfGavg/CLu/g0bdvhF
5XZcHqF8dujGzWfcWG7M2fe5/kxbY7gvI6H1arHG3oP+ZLl5kQU/uTIoppVvdf3Ryjw1P5ghvAxM
XpI22vlD9jkZHqqWgLK/mt1Z0i8CXY8K6xhBPcWDbAkidWA2RKjPOPFRYxTTfcTaEajjzD1gsBDI
EnA8+QXZggSmt8rcnDRm2w/E1CD0D1gv2dAdrZSd7+C+h1BzgRnqMOiOzn4jCXdGCMf4ozcc3Cha
uM3EhGD3M2SIp4shxb8gQ2IZyvhK6WA4uqvYhYZMul/DmY44P1PY4h36A9LF1KPpYT2/k/xgXXiF
DQj7tcdbgDqK/H2DcgyglskOgE+YqwoyHVJ05JojtzCC+8DdZt6Wb4RM+7D6ktGhg0af6aygHHnh
LNvQifZPukq8HHq2gjS/9sXsMcU/J1ArvkweGPiOCMXSEM2doagyQVnBx8jcu9QjRhPK/bGmkBdN
qJxeX+TWbN6uMX9tVA3AR7jXj6hUrjCDBjyP6Wrgsey6oPRX4HMvWF+VdTVTUiMmjfaaaUa0i+WJ
6xVbwtr+kkXDdxFdFgWHUVb+2xSVzhbMr5zCL1cpP2sfTqq/TOyWxpJDENXji1W4deiw3usbtFLT
1iweS/IgmRQ3sWdgoQ/KZ8rWaT2eqSJktbvqWcEFwAsA273RzwuMDCWZgpNYb+tpDrqKJD5ApCW0
ws8N74FVUs7wBkv5bFR2DQO2hX3xyr7c443eBCPgc73lNwrEcK1rZnC32mljjny8tvPw8NJQVHvz
0cdkwe9DYnrWCHouokFZNKnDFjzJ+DTwyHTMCY+cTiZ6DL56BopA3s/wYzWDecNnwYAzjNOT58k7
1JO1YekCgbMfQ1K/6n9FtjxjfCdH9iVbhQJGLy6xIQQo23JML4qhXqk0yHN3JYOFIV8Q7Dz8U77L
Xxml40j17jQuGlbNjMwG3kxJmC/GC+/8cMybhn8GOZLdy6rauWue1JlysLUdC0Vcf/lP7dOd0eS9
2SnUam7RKqWEfNaZFtP92Y4tGs43cfFnBg/rCXqpEltqBK19/XnHsWk8hcLDNThb++6w+kM4m2ny
WgQvBKwGktWS8b5+ESUbFuncEcPONLJRvktLiXQgzvwLmQ1hNJYLz6Yr7KFhoNAR5/X0F9EMnnrs
SCRm9Niv43OAE+xB9ykffqV/UGDRMoAORFhMdZdfGdxATyeEI6NtKXZHmOkUI+uGgkrgvN68b/Ma
FEcGNhTru7nl5/pcZiAOaxs1YwmN3g+Ku7Vew8Ma7s4SL91nhov2qp6z0GVzu1ETA/sIvI9UvYa6
IMsDPsQS8Z3GpQw/cMLxDTewv5hKi9XyJhhOi7yQjPhaKSwNW7oQw8cuNnTypk1kXEyPBYHX+zhm
e6MYwG0KLlVWU5GTuWOh5iHUiCii2kGWd3Yv9L/PeaROSnpPqPUfxhTsCLSmYnAzn+iP9wPsvAdp
uZWBPhqGsDXwcGjRJ67dLJ2TBxOK3fOlMTrYcTqtRYnGJTckkJPLogQGtf9bROrePnD33xQ7Kede
5iNG8XpMfvgtq+sjCL7UYhNN1mpbAZStkOKY1+BWGrWwfQEI6YGxop89cwIcOZF1mN0+m5q1BDlz
6k4ioyyCJiX1neI1K32xCbB3w+pIWDpbGtBK4Gpi1fS2WZ+XRwe9N7xhQvnoBx3wXk5wmHzpoLPj
7Mq1APDFqN7usWnFwfhOdiYYrrs9EN4FvvuM0NsQMxYBKEV5bBrkbHSsjmiP9RnG3v3FWNWDIRoF
oBE/jdoGYTf2XmaskkHXAYPBJoOZcI8swmR0VyMELca+5+C+ZRmspJj/AV366QHz6UXmC5KCKYWi
BlpX6XiLlnSxslV0CEAUispUafxQzlHJnveeR7v0+q+x8+pbPXwPyzBA9LAXPtd61dhO1yDTvVQI
Il5B6dNoa359AHCe5Ct90q5gh/HZAULJqwQOHqKp/5UcHEYmBsQF1/ItinMIxFbNcE4ELPdCMjhZ
CT5Ki4wa7O5IfIZ7bmUreXH1S53CXeU5UYG6Bg0cy0tNmm8/P0Wn1zkNIh8axURpO5QWIilc/Mb1
haNez0hSRpqP7flTqZZsHyGhlnf4KjI58+iqpgWmWgffKN+6ntvy4L79NVBKoEjNFWOvGTUayh4A
sC8p3mZ7dlIAqYF6jxMvvoh0vNwRbDMqfNOxm78/I9QAG6MUQNKYrswDa5tx1ThcBlMmRtFUT+nF
qgNPmAJ9Ok735hFwNj8TuGTOXpbiGJr5VlbjM74KEo/Vxe9f0dpOO1fErziNWkVacNK8z4/gxSDh
O0vDhDm6bAoU5qpN8Xyutu8hjKGmvBRUDkdXpc3jmUWJ/Cp02JXIi7u2JTY9yu0SnwSoNezutuAc
fcRgKft8AHEVyt9u8XLeIFsA6Z2HEx2B1NPj6seoPL3DCHnZIhsxQzYUk2t7/QvXJbKMV5P1EO/v
a+eBfnxn8Pk/4lDfoWX8bOI7KsuQtv8u1EcimDRie0tSpUrlEgYszPiEYiA4vSRQUDVYo3IgYZfa
NYMu5R+yEIiY0qKyF4dx00MgwP/QZDvaxTLZmossvUL4S8TBk42eRO0O0QHe0vHIH/ZsHyxzpAec
Sl8ETgjV5yYWHTg/MMDq+Ga7dMTNjZtJSOhfvYvm3HgjjdExnVkz6K/RKoj2MPFE9uI7ySTK52hT
Ugmm0bdm/Wv1OYy/RjeHWyfXxPhmp//z2JQtMMnngqAK4SY/coV6OXytsAoKb51M7/6vaAWb2EOt
mD7LKXz6P8l1NUirXU6E35K+FAfl7B0NrTb6R/5IvxRQ8j8fQYOyZA6TlCEk/eJ/p/g2mEosRIBC
f41HoYdq43NgFUhBd/bI+cThxxadUcBnRlgBlqReva4oBcJflOrP0TKohYeQ2co4NbsH+yj1UR1b
UR8s8sxO22i1bonLtYGA5Kl7UuRvd/YwshhJtVr0wykBQpJ+BYKcr27sRvdWkOHPnkUlCHG66ELP
+uDiJ/owOH3vPxowoC/s3niQFT5uMrSFxSwubWu9QPgbT9vWGmoh9VukbBenizASeA+3vyazd//j
X8GTcVe8bEB+VCNaX7D3/K4rTDqlvHBP5I9a3RWYiI9LWlP02+SZ0fnOv5d7AbYkqawkjW7Gu8rZ
TPF0Wgx+kcH1p+hSU64OtrcCuXzthRHuSpDwcWNiHQMBm1VBwSAvRaQ8i3F+tvysAqWg7AuFFctX
fypUa96UpN/wBiGMA8KQj1QjsKS25rD7k6+wVt+yz9z4F4KHghbKD7QheFqaO09eJcwIHpD4v1gz
XVFhzEbCh2D2h8eAFBacKnMqyGnxOwMOcUBhlxfWL433uJBvgwiodckM6rPj6japz7izcKomdJDR
TsZTA8jzMocRMORHyCFfkbLl+VnA+3b7ou/xu+P2PMgj3B4B1cGWF80FfQlk7QQX/NkrviKZoTqQ
Qp2HLuN7/d2hXul/yshJhi1aI+6S/qhytjWBQjpug434urdl0UUUrNQ2TrFlOlpJMoSdD6ZSh496
QfJnPa6i5EKtKSNcfOM0mJWoGic5LGV+sEaIEexINcRlUHz3ibU6qPOSMICh5h9mzE30q6EKyxMl
nFbpkfqhx7cxaLm0ptjePag0lTt5Y7EvaLUbNAhvRJ/PapCpmX5AIK/1evDW99oFFaOve0ANTwqL
Ei2j0PJWQ61IUKSAcT0T8OyEAvrf23cXP0679GwbrPEVqVLVKgTXoak0xjhnflkSv8MnicVDBJf0
7APezgBScz5wo2ucuTI2gxEwvdjBNBCfQ/M10yIKmAEmXTN2MUBPb8gvHqMCkYdlp2W77KsWpe8o
d3BLQWsfHhHv9XgyH4febelRivWfWzL3XqJSctlhyWlOmvYCPoA1QO1mSQVK698hSJDniJwOvMLm
t7azoGfLtB/GtWZ27Rr/SZkcGpNMSPKM7A9aLhsao09nfM74NnFqXjj5j6aWrXMai6IFUKIJkepk
DDZ3h1/eXVwkBmZK8HOlP2nmzG9pXlRWopxuiAxdeUGGMjf8MGyAlcHSmZLkTmF6LYXbV20ki9pC
ZCqkKlEu7CnPCkm9aTk0g3bfZ4H0Hrw5fRuOPb342Osj+fOv6/+szipudKmAfGkMkifj35fU4iIc
MNptxKhGPek90Uf7t4KvRZ1Hhpm40gci4EuBuHMh/m8tczmLVZEaS/vBFV52dNCfu3SnJXGUxpUn
MUOk4IQ4OnJnZuasQx1L61GS30X18dsGgsVjzfO0EXjQLoXo+AbxCOQOSI3r1XcUusJXiRLbTaag
+8ZF69VTTPeZsWMlH2Ah9N35BP6ahPb4efsMMs9+rX8/B0XGN1U6UXAjxBkEr+sCR7RkxnqdpsiR
PlnPIXDdwPSMGCslvHPwHNuvRRIeRCCZ+TGtPeuwHH0qykSEcFtINzA/mKVcvWlKpBYQtDjSu2UY
93nOma/KU7aEQy0OihI7o8McNoBdtM9L5vcHad0XcCYFSs39qV6vMPI800UuySerZHhxpZFZLTwt
kgOCMo6Ra1UHTNY8DX5X/OFLUuBB2A4GTWG2zobM3nzgF+mZw/qcSwOc1D+09SeVjcZPhYoXJO2v
K2//03d57UE3yHh5jVpCmXgFezKhjzHldi3DggzFuhcClVtNVkCBebzG8k7RKZIf1u74iiwWHXAy
UtxHKjTqNgaD7/8vpup5gn+X2lJg2rUWM5wEeLEdgR77H7XL5SfNK0w1fuew8eZ04d6WOylZ9IJx
h61X5PPqp/MMGyjBfP2NxG5LzE1FIF/EL0AcABZsTXMynUWNmlW9sCZAoOXk+0/sbh3PMyF/gMNM
UP1YA9q0VAh4/UWlCKAzB5AzHJAz1WSEVgZCZPkOg78c0IbHyzJB+1qEVXX5hRZ8sArF1hHEbc5+
BrpqMt+F6TUSpexmi7+UxC1Fq3HDhC/KjEG50ManBMQlG5OtljyIrPIWViy3JAgrgrDAy2pF3GGl
kGnr2y7JkBad5s81ggmvRi7Utr2K0Ub7Lq8jyXDc0C6obo8gEYqEfr9gPeP3K9IIUB7VgLEWb3Km
10p817EXqbdfXtz4BEMYyI9uMwYQ5on2IepgWcCodifkNrBm9vYvgsS3RBIFKPMdEVYB98EtiqYc
rWzxv9zkDh5m3pS5zzK1yWKs85ANkQyKROcAJE7apiFkvvnsfOqDiyOQTJhDjW0vkXVh/kLH/bYd
vRaVDnQaW+FteaI10GTNiOSvdiDneQ3HdVHfhZc1Wjq8qEciPo0l9B1UZzUX0k4jKCW6ujBUOCeJ
ucRF5tRfhKUhP9dmLD/z3T6mK3sg/6aVqquJV0vAjX3ArfqL0mH65wSX79hwgmISgpa0vnZGVa6d
A5Pr9B1Y14fCOSyogkWHdVYJWQI+KyQWzg1Kb13qTJexKXR7fchXxODbEGEQLqTm8kao6nBG7kYX
v+LEy23QdVDhc5KdYNV+MRhwdNMnG8AYKaDK5MCBuoZDLeHQOtMdNm9ltyQS4V4U56+O3Xf+wLfX
7UGrf/yJqhdlshg2UiQpDG1v1pH6zSGtX37s6eTEO+keTpI6/bHXO/Wh9xAKIZYMRkp/gI3J6DEc
h/lOjGQHe742orHVH2kHr8KRyCabriV8ECE+V1HVJGTrxcivqYpR4dnwemM6oImv08pQ2vz6hj8a
eVlX2BYzgUtYC0q7k7JSFWzUCYrLNe/9VSZSrExFSSt4pEZPbH3cuyNQx81iVtL6fk3vK//kq1SA
CVe2QYba/a+psIpIrkfLEPts7EZpDh0zl2vI39tMSfFjj5qv7LNcheowffcW1QJJiXGH445IZNju
f2+f75Jw01G3kammR8NaCk4reLgMf7ihxaHNRfFXFuecRFaHYQmOSj8GIz0bCR9U72TGUJtenQQn
AWVkS9Tv7HyHfZePEhE6kSoHRrpCdaJSOXafOvQbxFMbItHPa1wBKaG7aaImGvl06lwv5kpdUcX+
jRxBNjSkyawNG3YC9d301pc8JYkvJwIMFeCzr5I+/HtivG47pTSRIbgeHDZU1VwuP22dZw7V4ItV
1iFH+ncpRe8m8rt78i0VYTEmmxaKDMpTaWeW7J1bUGrj2I90TSuiG3ux6VwqAc/P3xApVdwjBUwy
5SfAtvtThRVD9q4y80UZm30LIE+LabaUwR+gE098f4CFaiJNuRQRujgUZ+E273D/2G3MTc2TpPgQ
clR0DC7kyUbkWIXjhUhkGiizFL50u5VOEw5SGxeHjYrFVmcTrdu1+ODKM4zlRjDWG31v4zuYA62u
C7dvXKrOdyMNWqf7H+XFgDD0YkAA9tie6evRNnZzGqteUcvkhN2bfir1I59gI4vLcWpeGyU+WidO
TmyvIdYYTGSXixfsF0xxcGKUEmNVhtFU4eDy0eBZGyH/gZm/6L6gdnMvy0jemYqbgk/AVtfQS7mz
ooKoMu/AGY8aRX9xvdgLQZGwQzK8hNyS2UNq8EMX+a49YgwyeblmwfKon2q0YTdeww/1KnW0xoBc
0xK5dHQ7CGA/SNagWplmV0mBGg2SHnSenE3UzsEklVt1n5O29OfJR1u5AVrYdnqV4AzWV0HQWM2g
dpbFH+MP8Ec7hdb4wEehwD6ib0PQ6ig/uUXMgQ8pHjQ2O0xWoNatAPOP5MmkxDVjYBpFAIBJH4yd
+wfyd5nQjnAPVilhN0+8arbq5GipWYBcRi5f9M9sjar9UygVgC9oHUhCjq4aVGzLMVj5SETwWz58
j7Kbk+QYWk4kKp9vFtpMQUQwkwDNnmW5syJ5ll3PGGkLwVmlw1nnimCXS87R1ezMTF9bXo2f2w8H
2iKQCMfeSmx0jmljBpNJuuuaN8XrbrCpjKyPOZfAlVgy1vlkXLedt63ohC2OVqNl+HE9P8PgHRTG
M/9ONxzIGfyfwGU+AsypiOz4npEpNNd3DLOK6SCs455MMBt97Ggp0TarYPGO19bWXP1TzgRLY/Lt
2dK+KQCxLzxTG0S7ZXOXBmCyY45q4n++ToQjDHZ7Nf9qwxSPM6AqLt/jKDRnBx8Kxhi53eo85/PA
pafu9FrXEKHrP0HCwt4hUnlFgEt2gDXTWCs7CnFEmgACT7La0B9daATj/PMmYGmYrGQNw3S43YAF
yBnz1DTX3lXcfhbMswhQ9TtGi65o9RH7UbexPLombuqRMXOqtIIELF63M6RazgrbTJp8Q+AqiYaZ
OeSg2qYuL5Wj5Gy4KwumZdP2hpSlNUOkXfeC9Zm8H+z2dERF9OfKFpHpJWKGntlTXSLYMd6AMWNP
NgAk3SdsAVsR+szWEnEhD9nh3Yglz4OcN17bD2HIJkfZZFgiNR9g5WMkQI/CzZ1DI4Oco37R5e2Q
GQtyRBIdxlAijA3Z+xr9l49WetLyTS1TbwjA10U4IoPrc7t5FH2m9Sc0lDEbugjYvq3b9XpqRMni
/dnelLyxjqPFuh491JXYRV1J9i7ioNqINXgQ9abv9xFI4KnGXlTDHiKpWQpFGLCmAGJF4Fij5w8s
pFE+pBGH3J7MlNA+iuoG4t76YXtqN9pVE59Rz7p2y4VVo27aTT41QuRleI3EkC9EnzXhadqw6DCE
2MLA854YkWZtK6j5y5KSOrA0DyrjFNbjtlN5vSROT7wVAvXiIZwQ3z+o9Nq//KZpqJkHsoGtw2h1
SYrez2tSjUnuRxhP4vsY2xQOJ7CMSlbazZeIG0jehiy1lR68TGRP9jxp1+NpRLYjsCMaCggNV1tZ
ITmJqCo3VuxyluHvOHONHcmMcsv3PVzwwyPFPwB7/ajEIGoaL4PjX5f/kHaQqP383CWfbKIkscVS
BiW8z6llbmHVCbI4gBSlZAX8JXyp2vQLx9Ou4SIVmUmSv11eKWyj6mUDkfwcdJVdenNANlgppg1u
HdeMuzj6kZyn6UrLD0ZHRrlZenLwym6Vi5U3/GBbkpd35/BTHkunPYXLg1ShHnRZkE5xU7x+Df6i
4XVKATezLSEdFYU/gL/fQDGKXNll0o3nclwSoLAIFPMi0i1N6NWhAErL5lDP7o5ZvUMubLs8h/Vb
YvIY5qpANmWeuHE3cninN5ex/X1I5VK86DzylZF4Zd0Hk2Y7wAaWnveBUUxj6s2v2pa+KKiyEH8M
pJbBCCCh8gVwqWc3Buo0atIxCd9SaYzqbs5BjQWa8TtmWqa/IdlpsyK/O8dt83S4S7nutOv27OT7
FCJ49y9AdVXY7VTQYtr3LlhExxa0f3FgQIrPyGkW1OIQ2A2rPOv8jPAmRRS4dBRLJIVRkC6yqeu9
7MtW2D8bmA1/6KynhF1YLL863gNOhtdK5RBKX7gpZHmH54oULcvVv6Svi1l64DJ7gnlvYZg0eUHP
h0KZvZzJ/93VJpA4Y1onHC0Tll+qDOhd92dGi1oGIYgz4LMvsFJxJxEQw1+eSpsEVJNaa/kOPgMy
nrsY3eJDj1OP/yRwVhL9Vplceb5FLUp6ZnlEmSGKEy5phj1/tTc8DP2UBxSSdvr+cHRPulQJ5y3o
ddSBMV9u2RDCx94KGheNE6tjgDL+lF12b3xEFgtyoXNAHTcmK+L73Tafxb8YhOBAG5X1N6dMG7AI
0ZubVxs/vVNlosonHuFRyXwKzSHo2vQhscyeHWEOjsz58oHR0fhFSHBadkrjWsz3V89RueMM+R3e
/0Po0iZeJXqCC0Mdgcq8AaLfhH+e6A6SgDBMdAxKZZeebqUBSB4uUWEZLbEu8PJIRxcTHDX2jJw3
5wNX3BhQqGHWi4SxVsUZE8aVbkxvzK4rrmUrqz6kvJDCFYsBZSWaFhqFUbl7g4zSfwXAKwhN50rB
u2V8VD1/ZrF0c+IZRsSi4UAvX4BcVrSw2e0/0l76V1ZXKdGp3pmX8IUuKA4CxMwyEgxQTDWfWdSt
T0nALzfZHMpQNvY+cGO3REc+RcJbVCJNvxC0mi8XUe/tnJRVzkp3ALbpFbYD9S4WX9ZN+bRJF2nB
Gb2+9pyJl8iNt0+9B204ieczDDpbWPy1HgpR8t5oelcDynASwFfYhuYCXnzJ5vUeoZW5Cr0X5Gbo
85uWT9qRZMHcE0E2lHS0HxeunfJx/P5fHT6lz9Y07OWbuptzAZOmpyy6KzDya0ePe8rsPqjLmLA2
Khv55zgc/eckWhP8gn6ysaeIXrGZJfS6fQtksMpbZDztbn9iA4322VfA6k1tAOchvCWvoHetX92U
Z1Q1HW+UPKZo8Q1k55L6Az8YZ6oxZvUqrlnDavdplkDy+xwjrE1Qm06ztwua8hOscAiVxEUzcJ5T
BBj3zInO9BWmAA4tGH35sD/UJCqtEijQYR09tdGqp9Rg+/++OnE4OGSaemCp0z4qp4qPMz+608Gf
168Nk1094ZJOUrOYA5lEmhFmQh2E4fsciB6/4a8++t3BZdLQEmFW46tHqHqYI7gsdlUMH8CA8d/r
Y8E6hAY6hXl8QM2JHP4FmbAHI1h/YLnlaHmaG9MsYbN1leiSpiG3aI0FwUsqInehbdUNsP3fJSHj
0y6irepYZJKzPx4oFeNLzZSz/wvB53fmG9kwJ990NLxJRuEb2sSRgtL0rSpql5RcadeMCR5wwGnL
XhPCoT8pa2a4hz/Ueevd2QQEz1TU37Nb2ydrwF3EShZLVTLsW+5WFKPzcdWqdf+caftLvfCMDh4t
hI9z+UydXMpP6azijZ7iyKrPnY2WTSu6TRrjKrDxNyX9FxoU21HnwqGe7w9eYxo5tHbH7Oqwm2KN
PBagmQ3ZqQv3jLIc04wkPzgYm7byLPAZxRKW7rfpXnQr+yNtMYdq/uT5pJL7tgLR8SNHQjyoQqnB
RNFWb0+l9smzVWKeIh2mpt841XkmS7iwfGUstWm5duOU4/qs+uaA/WNhFLR43Xb/so4WwoGUje9B
NpWenKObTekg+drCxhNfYupaz5AUD+1bOHcit6R1DO4RObepL3cfAsSLPd2MfsE5oJ3RYx2P2Dli
MOEssmI+lMBh8ASKGzeG+wxSNUqhKzJPURaDHxlbtcEGOVdmvJud/LgCIG9ciij74OHgQE5py0fU
LMbVtE2ccOJGSawWl+479Y+/aEH6bb1A4k0E02WZdvvAoWJxmWQ0zNwFbLEVIZmlLx2rE4XBQCJ/
6HJefPUtZd+Svr5PJikF57aRJ0xSTmQ6/upSFkLAMXOmZE/FVM9MRIcBh2otj4NieRYfDP6xlhaW
SOWddwmf0w+cEaz8U4TgArtvbhIXK72b9s/u4tY749XfPpxcqyjgXeIbsXPl0gLCBiMpAz3Pkyfx
3FZtRUqcD7BEsETFw6pPAqSH3/JDyBMZ273bCGrh1S3OorAHGkHjPpGxIyy7xxiRx4HgBy4+D9Oy
FbJKgFdIX66Ciqbj9FYfz0eC/Iz4Yg4MpQH5Fm2eApqEGqOml+tvEBqeZuxjhT/bN7eMTTZj3F6D
7ZdM9P7wnpRW2e+sRFvmzWUuBdI88FYDHPTfWorYmOsC82DrQycEbp59BvE3+yWjVyKrIfdFx8Tn
rkzLNFGxCMtCqqD5SzbGlp05P5KCyoDyvvFohfmGl8vYK+EnP8NxqpIgTELUDW8NXxlMMEsrI92S
BJw+SYk9aJDt/N1QzmevdeXlsS1AvZXAPf/ZG8fD9zPgWhTBx4pu0FFRtgblGsLjeFj1MpzVPlKd
NsEon4e5QiC7A1HODZ2o2VcKF/Q/6e7/WMJovFRH4oN0cWHDrj5oZzSsDkP64avUBelkTUyCQozR
k1Bhixbo79E7w9ympeBYxSrDWhNnXy6iXc4LaKnizbTEg1vWzithePvpu94ckgAFfmdAFGpDW7yQ
9zY+Zm+uhZjxna3S2gM+5sDD3rPRmkZyQv3mjfU1wyrft+kTvyniRZc4emFPWB+YeWNoBNRJt3/H
5aRotKx64DpYs3tYGek8WuA422SRc8vHaV0sv09FGOZ/Wvcpg3PIXX7UOC6pXNvcmf8e+JDhJMMw
Nd02A3Bav1D/22oDJETElw3BhB4/HlyEoojjSA6ugTHzAkpfbHBmvoQxVKxq6Y0v9wuEtqf3aU62
8cv5YqnyDPf35C2Ifepps/JvUn9NGrDXy2xL0GMqd2L/RmN2JeOiqo1vwkeDFOP3lljmWk2GkLof
FvHINYwA38XWtmnM+anTJrO6Q+fPChrJH5HhkgF5d9NkxY4zV1zqf1BPs85lmjJ4wdQek7XlWgzM
ZnIp0CProFhWZArS76XamZErINkhsYQUktkaeLW2YdvWywkorZBf4It/i85+vJCTYv78zJFwcq8L
upLeYRgDHqby+mmRe+5PbErvQTbG37P2GGAvBQ4h5WI7/OkhzmTw0SpI0EcMimyWCQCr/y6bQTRL
U4y2jLe03hWixrmtgYsb4b7SJERPeWcOdrvWywi1McOINZ5F076auvYJQmvN3CNFUpJnQZYN1QgW
Fo1Kyr+8Y3xEJgXZSSmIoKPFCBIt5KhAm1qv5D2GkwcQQjqHs65Hdm34RHkVq5wqg00RstQVew6I
ohY7ycXaoJw/QX1umBnPo2rjoeDhMTKkX9WStOGresCR0Ugt5zcQ1r107LciTwPGw7PmKVDPtImB
tM+lDthHqG7XDmnMfSVSdkc7YkwmakM3ClKsQXydte9w4zi5QZ3XHcaV6OITJZZ4ikJ8/2KczubB
VbbGA6HbkV5MmtVHEivI1lW/UL8YXS25SH71VU5/bnF7DTBzcWagOLoUU0MP5x5nucapVPl3lvFm
b02J4rQnYJlZAeXCqKEyjbN81LsxAKvs4qNAQ4h+KTRrdfLDcWLZkMpND6HFjA/CZOk/h0rjQ86O
xp4Diaz0d47fF1W5+RDr3b3HGkXoAqZ1Q8nU4WY36KRqkcsY1cpI+uH5qxh+ds1MLWhnxbjYhiup
5hv6Dr+TUo5XbUkrajK7YCEMJxCIgp3jatPI3oCavAWZ1ovm9k6h9xGc+n+npuqeQbexSEEiP/gi
GT+FBQAibr1D0pqAvsuhU0baWSN4TrZqSdYZKnTAE6Q2kkuMrneUX4qEMECuXUkvPtFCd8ool+Fr
B3ZYRxhWpEC2Dk703YA6v+PJf4faWETWVGlopRtlk0YMgjydTe2v4NS1sF+jo9i7XrGN0Uegtg2S
ofnU10xcZx6tggCP30jWa6bLkW86aUWzw5qedwdaeK7t9Ez82Ca4BzaPzLpcpqotajJQeVvaDN6L
vZqY5aOaoncR1UMGfhT2r5Knw6SCW3km/ZePx3N4w+dx8rQXb85/bs8p21Ic+lncB32TUQUViPy9
KggRSr+zbfaQ6/CMysoZWQmPmprmlf5UYwZmoDbND3hRTo3DmH/iBsQyU0e96/LionjH2+L4fs17
j/n3SPd1CTF0eMS9JCDFeSVAf0bDZZwxzSzC78jnzzJxQ9F2PJnRN/IC0dfeGwz9XbZUcO0yWHL1
YaHsHyLhFBNDc4g44nFWjO21g2oh/b+uTGeMVzBjarlWZC0WXFM3DN4/ZDHzQV3+NEbPZQpx1PYT
Ln0hFKRVtVwdR1DbtP6IyhvVfHIgcgOeH0QV2Cfc2ubAgh+0epO6pB0B0YJrU4SjsZxZ94RXRBaK
UsGT+h+aKCooQeecAvu1yOo5D9FJ5a9XJ/FW7/Q8RuBIqVbY4YWw7DOQSxr4k3k4dxLS5qtUktqH
M9Uv2rkNlO0DtrXbnaAzUrZoJzFHUZ/RpqiGL9vpMGZKY9E1JEjiv/xkps6KnUoUMIqWxi+nClzM
fwAb+VJC0ygowKkHwryUF+USvn9n+gcBrfhp2+io2rFHpkdYU5O+P7g4wzguXo9VBoanicLufXnu
yE0POSYxPTfqhdDYhFJxEwZgzIFnDfxS1LDakSQxwOrVYYcCps6EukvkNvDl2/YsQke0TYDrEgBn
IPN6CzG+GRzm21JmVhClDhk+uGI/pFXoGZOfo8uzgoCLuwd6TTVYXLCLmrSe4u6IDhyw/iREvi/K
9I8nBpF7Yeb8ue+XtsqHCvfwyW8gS9l0oDSoHUqIl/+JWJvAA5IKcOBY4Y8GEjXGK/Hmte2nE3bt
otEsi+xtuOLvkBeOws6pjVi7HA9WsFmLn8zlqbMxX7O445h+p+QMtX+CyORtOqb4SuISyGnh6Pal
Clx1yz8SYB7FsKSf74Uu//rIn4itFg8k2WVXELC+XgZK1oVF+4Ai72oLkSYbhOVrmWDzRC+zOuEC
OlGk5n91rU3NcFjr1ch9zaep6WzFZto/2aT7saK30OeKh5SOlM4CDh9+tUyKddQBZ47YrdriSHnk
hiGJe8mf2cDLCeIRuIo4Tb+yncfu29fafnP2b+ZKIG60DwHmWBAuJZSaQtI/u7ee5gbvJO6G66Qk
LAoW7zNth2c2nVv95rqYwhV3Mi0a9lPFfd3KmUk5sB+JuJ+8+oURCN8/aspou6sqAZU8ZrK9L2Rp
jzh48/LSCtFloJC58+ugEOSfVioifhRpJGfMk6IsUziV183DsfA1wseUH4uZF/jzVvs6rTWVC3Ri
2AKLx0JAf2lMK24SLyTXZtCMOP9eN416qqtkA9EgLzRKWNjdDpbtRAhbChuG8DFEn7Ke60MTzqaz
1ZB6Mi4v5wmlyIRhWOS4UQaS/ZL/oaMfpi0jf3zuAARWYiRt++4wPUIFORd09Ui0HbCmK8yflKfo
w6L1fg78s1pn6npwyydhD3k0Rsw4qC/EvSuF4+xN4asA9azlJG/x/XqD6HfJEvBrcPoBNWLkhIYp
Em4lzLOZbq9dnOZo/LFUImgkyEOM1+KTsWEDdO17s9ucI1fY9GsZT4qz7aroGg/MYp9zRfiF2Rkx
XM4nEqEjGn3N3/8z2UM22x9vO4e/yqxfUWucIkDPpmA3F+zOducbcIwLFlPLtMJrMdf/qd9Od8dz
Vl8qXPEf/pMyWpSUWvnhVdVJKtV+ePVaU12GMWUitLbn3ixyGmWgzcvq5SYQHb5uVI9adD/3nj8B
f+4l4dZjxA33Ijgl06peV9/BsoKUcjpTCM9wgGYoaJ5GEdzZahHlctmRnWiVcppAgSpmyeoGIsPs
HXwUu2KqJUqyqamtHCiafviirmatWWbe2T2fllKZ/1+GLe7zJwm+gCfGiXJqO+JmIj9BBopt9c+z
LdooiL+mY2n7hJjoOfvmGvk7SnADpk0w9VrNoUi3zfFhMX5cblE1kk0YXtT1WZ4Tn+FxZEiDO5QN
OP55N9pZxiYI+FK2N1hYbrQ4GlB7aouFZyc9dPlQmlCxNOP6OsE1xxq4mD/yqO6FRmv8+QjE1Vt/
INX3uG8zmHnRFbp7gs/96JQA91uJFdpz5Z82IKG3dZpp6cvZK9WPHYjBkEhEKHvF0OxI/09r9TRl
fTc1I8spLEh/C4UQQ3qb9aPf7MalFEPIMdNkBpemHc1yJoU9GuZtewEPn5C67DJNMf9Vd3OGuBrV
cWix6EvD3/eTb8PeOWxQmeuCwJcCToHe4UBdYMGh2UA3D8AtCSn0PUVVww2A2q92r9ycUYartk1m
lQZdvLAuvAPBNdV2hEZGpCqd8UM/OhZoJZNb4Hn3Eu/2jbSUyGzeVuu1HG/ELCi7oXG9ZCgthL6t
T/NcsFzzGvk3cqepTwQG7MxwV8BhP8o8qGfEaIdC/aO59FNX50EQ7Rbacu+MHjCHM3NxC3L2A9eh
F/8CVYz8rQ2kmbDYNevzQo8n8vczZ7iLRF2Y6i1/CA01pGNxEXn3uLxqV5sxONRXZjKplTkYN7h4
ARpcgUkLrXXpeQQFdk1JQlKUMY5m+erVXMrH7eisWfXam64kIT/NlqrHjS8iDGYvXOVR1QQxpySY
IBxIly36snLAd7T/HzpX8wVxE+jouqJHIHeDXsdjgiHqi3S35KSO/CVuDyC98+kTSdb10KB7N9yz
phWDsfSX7IlYxpaDjC04TptP4KNktCjzvFu3eTfP8a/yYJQaLWBHMwwk8O/Ove5iZBezH+wGQD6A
+m6vgD3xrnQMP03w3zEj5C/rNC6xGKfvdXEdVEjJBSGx3JVgnQC+GvSfvElM3qhFqPuroANrPeDF
kLeNbRPpo2vWtMuyDQ/i8Ra4SHS2Jr7GbUo414Xxucg+/GksZpCYD+RuAX3OI3ygF2BEMtZO7D33
FDlIYfVDKYkwQldjqcRyVYZj63XJUVOw0kMccVm3JlOx/Fv9AsnzCzwdbTjnoOuoVyspK+sV2bgr
RgfPK8ZKIOJFSqWhCCxDR3kN8toW56Li6ukJ9eIZC45m/Np673AEqQ28GxcJHIdz2taHlpKDajXZ
CSjH46YyxMcG/Ug0jdgfY2cmHA+mY+LhJoILrqoR0BqmM8nzFsZPaqN9vEln1YN7hFcrDYSpmvUc
K3AX4nnhl7K0Rc0B1Pe4TZZToMaM/k9y4/LhKRNjRdhJvTlD1nL3WJQ+ogedEbk33aOoM0OYRqQ1
mwIrl3KvW0GxlB0nUYpZAGFThqe2q/S/G52qTYFu9pu/M7SHINV9xu29OOLcXgbuLFFCMozxtHd6
jlqmAd0S8092aGOvz4ZuT9T3F/7xcNcIH7V6N7DMXh/0wP0ODunpwAU+KNhswUt/oaobAEHQ1P8A
XZigV6M9FHeefwGBvl9ZgPKvqYEpVdzqQ3gMYuf0KtQEkmDK16xVCTVqW6EQD+qCBIw9XZFIMlGR
U/c7y+SDk96GViYeEcOjIufVAZSe9CxTSOh5xgR43JCw/v5HIVpclqgvwld53heA6pD6M2GLr5xY
B7DNE2kS+5/FkKPROp+FqVla23bUSb4bzazK10NESrOsptO+cur2oDzRaSivy23o7oNJdGkpTAN6
m54jD+NNTJMl74tvrNhCMHHQwn/J0LV1jMUX9XUaRKcfIPuKzxo6m5zpFBlwh5U6B3/IXmjGJaQ6
GUM/Y0LMu4qF37Z9b07Tj1zd6hWn4dnS4iXJ5nubldbbCU+/CY8t56v+upW+NezwwaIu84OO2mdE
BxM0Bn3QyoZmPAHKvkDYGkfa2J50FnCToqGauB12KT0sH9gUXePIpBzJvvJ8MhlgyBFEKi6gASjW
ac6WZj+j3dRpgKgs27+IyTPgXqMdu4OBeYZiYSkX0P+LCqcVnmNLs9gD8sbuWdGJghyWHw/7SO8m
3M9LKBiPq2m4xAg/b/yMdiWiN7tj2JLF142dZcr3JxlX8uAwYkD1kJDczqesPQHVA2/ipdbyG9yK
RZ+MbLWJH8WYzsOr2eD9yE2rtv9AVfK1K3lfbkXVl98hUJbDCHJvNgjiL0Hv6HjftmJi80bFRmO/
kcOWRilF3faCr+lfADKwXNHAqu48JlXrRwnF64P/93BLcQdzX+gouyOm4Ipyiv/VWqf6iDD1Vp10
QIsH068Lx9vJhm/EwcYr0kIxnaflLr6MG/hV15nyEeGSFe2x+1H0pRcuUq10NqiMCcaR6BPBFxqD
do2OlVn4/MSkkvzQK+bQjvL1Ucn8Tgw/Ff2S9nZCHcQv4z3e8djF4jj5RygRDCsHBs3ZwpHNas3n
sXDzmpLz5cU4XumkNIimqWV9wIOs150KIjerZx0jcV5Ipjs5xx2ml/zGVsmYUPshLSi90vgel+Yy
WAQe09sxPYP5r77TDv6c5Pt+62vMV4oFOOfQG61MJzAPPcyMr/9bygXLI5mxmqaEuLGY8HC/5sHv
jbiK3hS8cpzBKhEfmNtnr7ZbFGgdziI0+rnpcjNmKdi4zpPmGSSBTXcDuBu7iqCoXLbxPoFU/+uJ
y6K99AbmDqb/j7sn64Seu8KUi0Ju6+NcBLtTe3iVaQdVVt1DVeSzvWBOg3A0IhzIJw/th5exLkxa
AnQqvoRlgfylZY5+un97ObzxKtK2b0sGqjLc9hjkSPTEnmH3HiSUVJzzQBizHfmhkGiDYYOdK65I
Y3IqgrQy7HxRn2tMjvxzLiNo3Z40e3YIDHXCvmXi0NHPSDe8VZDD6GlhI4p+GuBM9vpG1Eyty4bT
+ujVZ+ZfFHzUNK9wkQWdqJ30x4vexDolh81HNRA3NpvRZyzYRCHyNl45ewxgIHlUGis5OJY4CFiT
l12PMXH2FN5aex93Isvxa1kRRPM9+6WlnnM+NyYG7mw+9KU5+AGjmtrC2RwLgb+9sNmpbx2ody3p
2HMxec7fCEto4ZEe5UQWVx/alrCUII7BdNAOpAQnzvY/2wxPlB+wXSJjUJE0/m+bDDmZ29qge6Fy
zJg6o5ZPb2gflJ4BO5bC/IifMaPrX/Y1tHmC4A6s2/fKKKfGmPjdsyl5EMQDWnX9xJAgRM+EDKyr
zjQgtCoi8NjR6ycymi/SCo9ygIeX3Jlq5bobdhcWjSCIkC1PHigGfHY4wJW7uwN05NL1TdeofqtF
OmRscU/vqisBS6hX3tCHrT9yZzBeBrHp6AziwiNd9icdgJQLHRPTieUym50+BCAY8+RRB77b7N4y
zh2wk/0U1gBRPTCXtBFEiAqeMXszfUvzTQLzDZHvqYkPO90owtyqftcFd+Kigc3sszTqfTceNLKY
/5q5N6I7MizdmPhFSpBKDt/co39FMlZ/gKPWkZ2qgT5+2+d1J50uw+KTl4P9UOziaMeREb0lbtXZ
gBaazHRZOa1+FX9p0gINO+8twsetWF3/koN4ulcTQc46CmZdvpy+2ezkklBCeEFF6WTpmizourNt
DLq85ohHRyd2Xeoh5OlpDIYUb24YbeAbsUjOqO5mB5yMUM61MKPeX4XZ2P2PXjXt34LSyivMHgk+
DjNLh41fUtyl4/WGPMIfZWaxtzY4MlZcNNMw9TgpR98FPeK+G6L5dbW/9bV0CTp/mQit8EXW6ytZ
o3CxvVfaiGG5XipvDMy+0mkqgGw4Vg/m4Gu40VcylRYwxVxY6jgzLNBTZUvPpkA74+WpHnmsDdbk
wAcTopUBQBxtDmIR7CIzS7qU2lFEH1fzcHbQGUFVQ+ni2hOQ66gNg9nxEXxw8g9LsnqzxrIs6Lhl
uyplZPZKcYo6QRk6jI9HhtfVWaj3HNF+GXIg9DNOimlY5k5bVlDodU59XB9Et0hcBUINVhDpV7Ns
9a2UOJZhgfcY5f5okc0kMQ5nC+L8QVDTUAvWQW/emf+0TpRs/xjJT/oxsECTnWLPjUgBaxdOFfLi
KRS9WkbnkIbNaNg4i7xBuZ/XpuGnC1CnO7tiiYt2OUtB/B9nrYs9KEucQ88vfKuE9zndBa+3nWh5
woIn8mmY8qddQpHFtYvyI2fbyV9YGjJMPz9UFc4faWJ5Ge/D0lKF3jzlWcMhLA1Ld6y+4Dh2Dqfc
WNyqBwTAbXoQwG5sJZUpDq9t5ZtBJAdCh4XRB0XLnKH/nynX7b50ee36YaefL8WTVA1RZ50T9hum
kGCEna1Yqph5So9Ucva4XC/fFWtNNPafzO1VKrSJzsaadm6QScPTlgFScPvrqL1Hj03PLO6eWg1C
vcj8M0QOduTxOdK+ZpocUeYFpagnUHKKv9708wipCX31hDi4B4UO4+JQTsicALBRrlPAOzsHpeF0
qS04gM6bijXFZ8TwA+Pt+SwrVN/konzdlSAyU3UFpfYw8qW5H3+hzCI4QQSywrsDJvocJOa10T3A
WRMC98kB4CAXYlAlU4z+JJdSRH0Zr4P9KEu4XcoChPnsM5VDAayiHdaYSEesvj/Y4xF+4uvuXycI
olifaCzlxoOQd5asqhrry6WcbDTtQLWj/QBX9w+khZpIlUaSnPs+CpVs0mqJI/tUQKEBDfnn+7fv
eKVzmSCQmuW7zMelW6QP+IZE+/Ua9RArXrnosz+WCQO6BqzqIHsSbwcmK3qT5p7pbHW/Bm4Sdu7i
K+GYY4hyEi3WKqaLk+GYihSgZr0U/JAg0GTbxL81LQdbaZ+aoF9jasHm2Kw8m8yNK3FcxHoVFhri
XP390bLsZAIqbICGNyqHqVbOPgtv56788FX4+A8ibds+no7tEmAcSSxJftGtY88wB9WHSTYa0x2p
Ga8J7tUpUBIj5dr8Q7NQSeRDSDJLX4B1ndewhCP8sxDFUZcErykTC30yug6+qdoQOg0yFu+WazHo
tdh36ov3QFk4R6o98HailGJOlFhDqjR+zoid8vnniQe8wcICwUI1/R4LgpRLf0iEMeTSthh5D6Ry
NLQ5QzdntAZmiqcrDqpeakx+lylu+LOyxLhTK7fza5GnoWkVRbuDVmGgNTtMwWPAFpG0C8FNFOiN
YsLWTTB0l7epfzHu430Ag8rj7T1W3AP+Rw7JVnIyZBBxBoZrHOA7CHC4xTrS6Re0kWrDupeqjmOa
l2BmMMd1hYhSS687Nm1GKgox9/TF9YRrRa8ztWVozFPJyYfHNOWm7cbdvl7ygK0yChXBpJQO2Ni1
A+f1WuLGr3tgt/WXIWbWsLhYLLqqkWNF18cH/WeVJpd63/vMsHp1P6p7E91se64ZVImveLRJfU7l
Qze+cQxOEkGJdF0GZNRqWmQaBBZxRS66Vb+hARq/VmuEKu50ytxL9MPsfpOvfpcu/ywftJ+EtcHE
pWJo8rSQ0N9COaUI4ey/qOzQWpbRUk4/aHPNCnobzru0F/CoFwafb5IYLX3LZ43w3uMJ9ROkE9BX
pvES63AFAzpBgSdvdG3NOFuzsbpbDvcU45wku848gh2f+4L4Sef8RAGrKhecASb9iwm3ON0Q/S1q
AXF8OhHDSrX7gt8BgA4cQTfTdEoOPxxgGCM/dP6d2uCd2H9XpofmKSmY3osYDLPZu587+7zIGLWQ
pVuOqkbGwUfExL6tpoERdxUdGPJjZSX2cHHmSy8hfwJX6rvoeysiKMa78O2000iQqc4vY4G7F4EZ
Aah61oZJSgyIVJ8hRxovt2ckXk8SPKoLvTcQjr8/2YeLtiH/CH2k3pZM+MZM021JNoH9QCVfEB4Y
tfhVK8k0n7XZFrd21SqDUA8Z1rUL0ESTgb9KCRa+owOlhRigi03dFP0dVCAww0vOU8q8Njt+1qof
ZDLb8/8L97/O2IJ3MFyeBPRCcrwlqCBWZP3i1OD4Ae3dy0jrLBhsk2zTRv6PJ+H+dZiIa6ErlH5O
SYVkcT8No5Bv1e/gFTixcxFgeDP7Z6y2Fljnm9jX6hVFo25p8FmyXR2TaiVJWSwDMBWJ4sOAOOu9
njFwIquwxZwvR1WOG62FWsykHVN0yYlBw2QJLOx00zlb1Od8/GNG08WhmWVt291J4ZsFO+hMwnU3
TR0x/AlihQ1MrT3cuVrnk7jU6koMqO0rOJ5AxwDBMZnRXwdUsTPy615dyjtIG3KrgHnSIQUWTxK5
tcqVlr6FBWRHSO23slkXei3frIdY0YttqUDBkEwgvLF2qst6hShFznpS/Pm1o6LXP1wvbTRE7C1M
hR4frhzICpidNyfeB1B1fup24lkesT5c6YmGRiOHheH7V0uYSbZ+YjMF13QNOmzLJxFylSrsU669
JkX/E4oSn3p2hgVz0vmVqYwWcpwtsuMQTPcoOC6JZuNlkHYnjZyfz+1E6VQho1eBnQZjqEW8Iixt
srYWEOSVXUIq9KYsA2NUWfLJfTKrJptSsGOQL2fH1nE9wzc8Cy01SbmjMgyXXZXjusahZjgc/lnL
vILjQPzCfvv1QDpwMdnkX7ONQdfTFBxBZsSfF+CAaMWEr7kiArASzDif1EjBzNUKdkZMSlO7FZ26
UY91hJ0RyWLETXPx0zIi/2w3pX7z3nG0jtKjM5qVTqmFXswPl0qsWSSQg/aSTNu3o/zihiYqnQgW
/mrqHgJahPuiDMpE3SuerzOjtZxZ+plb0Ux859b7DHELfW6RaRdcaoTwQBxR/pAZZWRg1g3UARvU
ElqRlX8Ef6isPp8VRprX7yGpDhL0ith6m7pvCUpGme7DGJSHhZFBohkh9eE39GJKq2nHtvDjcBzf
x0LdgjI8tqb0V+0gzTsGLOvwtgrMvZtIUnE1KCB3pROyZbKUPgYeWBq7Zkkd4VZxxSbmoa5Ubgy8
4fbVMDyv+RNgnCFvvaeELcQkuIVKVIAmruc+ZvBDo6YeW3OeqZ5tnLjrU6IeAXIVvNE3V1UCdyps
64oG+D2UE9eHkGTqh2kPCGnaPFh/Ji9iFiPsKItlo9vIQ5r7fq9kRk7L4UkQzbMcxxT1WBU3guey
p8oidVGbtcbeF8j0kYhz+FkoiNE/ZS5nwOxvhDCFDabGzApcNvzmOdgKbjUiEBONKN1pXzHdwbSW
CGn8KJSE6pZnv4i1ljqY5X++iC4MrnGIi0FEEB1FqDCfIzCA4X1+gvYV3/wqL90bsJE4yXRreF+/
3JcDz/m+8PAkvuJbFFRmWq5kcNd+jwGluU5M2rEMRf/dgJQmORdlzimpslqhhI/7wKHCZm7MoptC
7cjKhICVVZgZE0+d9z8t1+aZZGwrtssjqZKPDE+nMJr6YQk7RV/fbHue6q6i/rLAa00eB7xWiKaR
D9Htv6bj6rSQcyVgh5hN24PxOR3CMyRMP544gvgonPpTXU3+8uh0cTXH6s5h0nNfm7ZzunPjB3QL
6Soczz4r/8BkcP7ISbGHzu8Jg4oBPGsKmKVKysjmr2S4PuSEJ0WeEGOY+/r6EjenxRMUz+YXIJZ4
Ty9gcQL9lu4VUNjKsL8SzW9Sxr2hE0mtK1GR3VxATZDteAtbgt09Z9K8SfljTFt0XDy/XrVkIE39
A0r/Uac55SqcSuzkMJGER7LB+XeKfc7gy9KnOCUCwE4FgfmG5/NeLTmDPWQPQRrN57Fs0ZIDV4HK
3UfvBCUK0I4EWxUv6rCykSE/0VflWFJyErlo8LLvlXDB9NeHTYfv3kSuTHMDZ+BE8IHJWHuVKUo0
FgFvrq21tT+/YddbfJwnVAlxqP2ihPf3YveiiTSR+BoXBQhpV3QF7YYOAVaCvNKCPIjyknKqP2Fo
ayvvrKoChY1olXNQn/4lhcrRrB4fucI3NUWIhUQeDJJjmYaYfiRQ8HA6+85LP/7NkguOCuN4czFP
mArexYdML5y8+0E1DQmaEkpn/jplthlGuD04wTsRwKERo2vq4bXDNR+iWYibUrhZEzlFU6WsV6Kf
zaMmMLG4aHzUOVW7UsLhMITaI9YhbrMjMSaX4TQzcFd8TT8eG82VnjNInIEPKnsDH21WZQnMGbo5
DxPuxtNEr6MI2EC7x6y1JQcTeHc9EjlxBnkZiGff1EipXudyG9WFTZJn1Pq7rTK77cvkIDqJklgm
MbBntnQ9lf4aZjRYg/IcjQy8LoW1zAdW/20aL9N0ZTmGzQuIO2Qprvj1+6/Qieuz/BeQnj9hTM4w
QqHGAhGWklCvfjMedI5yGpFoculAAX2b4Ka+CH4PXe+m2cH80+7ToFshayuLt9LNaYMfP/27xu6b
DTKmvQHpSYPbPpBj7/xuPtDcTNkZvKlKhfTUcQBTZlEYXGl9W4eQAlQPwR9qbHgFzh7275Jargnu
ZIvpgG2UT+N9npXksU2hny5ACwlhsCFRGmpozpT6QcEF0M/2LvhxIj/Qg6hJjfXQYlEETHcLo7Ig
odR1Mx9yEEWQYg+QATQRQxiRNe/mnWi1kUTNxvYaT+GzW2k4Zm1IJabX8xQUw/H7DeGarSbyC1VT
cg7qtu0e33rBqULWV9/8ln9r+2UOJur06VShdsU03BwnKkt4Mq9Zsb7jUXLOcuIaamtupNiLrh/+
DZWcMZcbdfXSm9Kld93k3UVXCtxRQFgzxsy/BN4a+fQlmL3d9Uaj3MjhNNL/k7Zca0MPy3nhwOtO
CUtXr5+7OrD4vgvbYp5czfewW3rbgd/WgVkDxh778wkzoAbOT0RRsblcuoIUeRU9T/gFFOcyg2Lx
Z88ACsslvOFAlQc92t7fltkfS4WqawQlYhv/8MDmKEvjRyXiBGp8DUhMTN5l7J7DJOnR2i9tt22h
PNeMqprr56Xq2L4Ar3Js1HTWwxHjPZE6C3iYCkKAnDez9IIQ4CI4YiJ4aVCaTfOMJofNofrTixOu
mMSRqmSEzHbRrroQ0qhpuCCAJ49X1Rm2R+Ehm30Ztk0HFSe9Rfdllcq2RIrGFzrm2vmnOwCMPDYA
3LAxTDn/q53rSmk5bZ4f/mxDidPLRfPxb1cJdVeSmD9qyYj9N3Bc7Uhkgawu71B9zGOG5uQgP1I5
KU78AVtlJlShObuhP5b+sPdJpba/f/hN6s6oJjHiYuVrbD46r03h77Re37DFwsNt4TqPe4Ujk7W5
Gs8/X/iOiH6xX8ToGPWurIdQZDY84C60g+z6rZTf99QjTtuvZGWT9VngMO3DkYPA/d58LeY4Pynx
rHtTSKSo1TkDWJl18ys+ZTLZm6QBDSllnENNGGNRK4tpchMEzv096xqMd2J05BStO20Aqwtsj4li
w/OA7LJVI+EoTLHe7iXmyRcwp9PD9zlvNrgAehmhFdg+hfnFuBXpq2rm75NICZS/3BNOzlLRWqev
vcmIo6Jc4/kyECT+L8JN2Ozc89CKPiGVZTSj2LvezK8H+JZHdgRRuqLGJAjtZ0l3O9BmodDP0RlO
JksuGUqjw4zkI3eBIPO6brAYCWM9lmf4RGe1rirDMfglNDgdN8QdIGNh2wikzDi0lDdZP17z4J2X
5AKPkCejcbAeK+4tx9BIMw6K+luRifSdC5TUqICs4F3r3b0KAOub04VNeZYVj0Yk/DvMTwMNrikC
VVX6773rXTbU+Eg4d6tY7sjrX3/u7qoknQkMvQcCSRePPhGu19Nq+owNz0cq80zt/Nc9nC29cLX9
6NL3GFG6y1rViRdy7PUFNL3ZP5pw3tVSWysLSxsq2HcJEAFXLi4f88drq1NJ0SP4+STNPVHHq45Y
M6ci8voPqBMr4kpPJUOS6lMXvupl4xjV+ZtwRF3GGS710Ipbg6W5J5rpzBNZG4sAyQpJDfEly+xp
TlX2rwePp6XnZ/5wMN2o1cZB74YJkHXsHsJnx1AjmipEvG9W7PnK6sOBa42XGgHXH9WGvAQ+g/Bm
G6oeD46EjSqK9eIMSPcpfk7B155yDfojsj+pyfIeQ43u2HtaJ3AUWVMX/Jrg5JSF3FAYU8O8ESBm
eZmZpKnrGsS25egg00+qrmyJd9/6COwFfLO+fPCezUDFZ18PxQQmpZxKzsfqGzydAVJ2bZYwdh2S
GaqNFFz3H2rT1Oik6JZYpMKAiCS6W/+WB8cIHlY83hWPPpoSjbjdMj2un/ntARQmyQ/lHKmANB3m
cwQ5nr8NREubpTGlBN4PMqLQ2fS4vUiLKtOEOMsS8uaEr/0wgLngGPBmxa7sQLOmAyq3TE6p5GIK
Rbk/+SBm3DXYy0inuv5a2W9/mettnHNEO/AqgVrhKRHmKyqUiQW76CshMJYm4WEU+QX1LAABeT1T
ZXI5WUo6flGl9TCpg8X/R0Bt1xOQPsCkRFJ/lC66Gse5XsK8e93djQTO4WGssF6btH1jHx0kfevz
SgGkfX9kZX9CYlqcPqwxRpcJvLUpSKIMEztnqv5zigK5db8y9r0BSYzB7f8IOSvMuRvSU6p+3YGN
tDW/4c2YusrPjfhSMjr0GcRKDw3e0Qv/RqhqIqCSLzfk1/2nGcExVSBOCOB+SHkJAmJ5wSU9iY+H
xrgd8jrhss5/mJjzThisMxYoKw+5l5TtswbaOQFSAv7i4QCTObVy2+e/XhSOw49kE1zmrzGuU5dK
3ZkyQN3FBT57h2Kdqdz/th4ICrEK01gJnHY03101AQa5Uh4Rryw7MFm19+WQij1hUq9yZb5usPHr
mtRPt2Ov4nb+LWWLiWWB8Pye9aIu92FHC/nOnOoUcqBbJShAKVTvS5ydQBDOZCAIUJYWpgeCLpQN
zWqMC16wOzdflE8SMBO7vpMx9wd/EBUCSZNGVxdvCiasc/tFxXaubzyx3Nd0bq+7PpDoJxNAjpxH
gCXRuyGEYDMbEAZyY1gSEiuV+4R3NYTaDtozYMAreRP+zVUrgJuf1w9T6hyk5/1IADRhiYzoEcxQ
lYH0wR1wxM/EERjmB4UPA3SfDqENupgYdtiYTp5TGVJF/L66VKMQdR8WDZgBs3vGvTJkUwteuCiu
NdwapVWFd63D5G40rPx1enqKYmtBxXW3HY4blBRq93uQjZuJaBLUPZWywYX+FMlUtpcNiJIPd90G
bnTAPkxZ1GDU6FjVFTBbMXhHxe+O3tOf/5ctWNiEFCcnDjV6F35JgCxnpZJhRhSzwg9S/4HkYyr2
cLp2SYaMoxDqUPn3FOTbWQJt4KSxefLEUJzv5tY82Dv5CH5pJ9duteJHRVXkow7GdzEmhgUR+OU5
2wqrMfFlDAVMpuLYyILY1mcOZ6YVLihRHkVRf/zr5t+u/LQYARjyDaPxogauvbzFk7WRUHMNcUtR
0xp5KidqMbgbKu7PPZss2I+XWKch8kFWU9qRT8wZc7sVdhBf7pWIXcziaB/uxpIM2y1owq5LuIat
0Dr/KiuwRb4ZXMBT7tW2Obwgdkts2AszNOLr4/ViI3eXlaqsjfxbUKO6PzHOyeT/qfv15JOIBj8R
pe7/LVlERNaxT7zrqd0V2w1fSJqyo2zGej/uShzDobr4DtJs+oU6SEywm3u9YjbRBVc2D7MmmAWN
qQYULQB6POObr57RIPKxrbC3sXYbXRLyBpesiO4hyUOuj/U/wdn8Z+6sv+8BKDORRAz3u1ANcReH
lpZcWQ76jgbMSDIkQUcCxWNVfw3Vo/qrh7encDnh8Kb8YVfpjtQ12aDhOA/lJa9P/q6/sNxZBX7l
judCoBM1GsutrgT0+JSNIJgPgSJkbg4YcaUzpm6gGRJAHAiuP3K3TClTda2FFyuXxeHhlvOTYwGj
UhfLl5KHInWT7cfFc5W/mE/z8POdFj4bPqWKmy4lIT5t/oj2/WgADsUKIRG3X6U8cKrx8t3I3TB8
HrBWdM7XTyzfnRU4AoHgaFJ5QXRJSOY3yQNdumAW9l0bLb341Z9Lbi40aGdMCDXP3ks+Cp1wSZiv
E6sF/EA1EhAhpcC0y0JkbmSK6L0GWsZeW5GH+H3Jkm6K1Jc9LtMdmmZbDYs246erD8llk/HqM4lw
E89MIE08WKkWKUZJJiGgZTbuEzq0Xpsc9PSkZ06i2qulLzf4uRYokM6mTeU3JrGwF8Wx0lGtuVua
n9sDIWhQF5nZizYz8/4mLOF/oZnK7l60IzLkf4euY1tdNWC/gp5GSuQnlAOdwR8KWhb5MLcwbzC9
ka7eLzwn8jhXDdFke2wrDgmAz6IGTe2YW/wRroKLhzNCrrZbTrnIjdwGF07W7CK3vduR63t4DMbL
fKPuAzj8a03jiLpC7FQBBSQE1CGXqjbKc6mulVS+A3ZzXQqZMx0YugswzJoYs26E9ljmBQ1Hv/b9
zZ+JFwEEDt1VTv9BXDtgjhra5CEHTBF9Ek35VWaHQmv16D39zSWAW3XzaplOJjaoy8jZOo5opmhk
5sxPjDIKCMWtQi2rGLeEkD3AmmmoiWaDRIWPIQSUMNcVLd1zpd33SowEvF+hIkPur8pR7ltzkAqE
BppsUu3kXybjS6IsTUE35ik6K2OPBLvW4ksd+rKG6E1HMzZnIZxVZTVDW01nDvm6uNrUq6o4C4p+
9dlEuqqOpiErw+/w3eoqS8KTvc8ZKbUHN9mWhCVQKtCjPPSFQAKvSZVxJUqhpDgA3pGH1EBC8YTd
URVOe4QXpIQg75YZHngalp3TI3Gac+Qfcm7VAJAoOlxT/l7LDEuugDbtIbo6YaxBK/jgMfFk1W/7
HnBfmBXqYE0nc/9L804xqMJL7wI9ztrEfTZ6c16T/gnsfs3gUV0RKanrWaEjOwq5nRI3uRYkuQEh
PyhEGoL6CcNrgCKY6p3YnO0w11KPaTS4/oSo50wZ8DbH4pRzUSGyGWQIPl5KdPXWz3EGWCbUDm6H
RYIfGs2Z2K6XsC3J4xxvOWAeDQWx4L9sBGcBrkxFesnYAAeL0cV/7/YqVgFN8Ws0k91ZSe2T6Efl
YbfGZhCh/imPfMcRAtvbi258cOcPcf15FcOwq2tKpOmki7fvkqOHwSvgzwfJ8lMTv42lsh7uVtVX
O3viyJCvJwcs4Tn4F7tX6852e/CAn0tAd9oimApZSjc512pdgPsE8/PiQBHPVhK4iUzvrfBzn2Ee
JCS4kG+k7c8omk8Vi4su/16ZksHr0BkRF7sZNQLAT1B0BT25pNqCpPvSPwlzUjrJE+RWH8C+2mNv
L0mRJXjwrdfdYMlerymy/eGywR1nXaXaeUzP7+lU5dPkIkDFP4eFpt5F9dZoRcMIzNporPvQjjsi
d0RR0nXuqOu/3RWrJ5NSjzSpXbgqD9QRQFjTb7yEPOIAlA9UksvbBAybEeIgp1QlDA18kiNJ+szV
bH8lG6IaPDTaZXuZdlb4Q+wDMrEfma4u168nALhpUtfxsPPMzt6Zq4H5ewu0QPzAEUmYvMKPpAe0
BsE9Sx491EO6XdAAafK/TtubR9l7hIT1t4MujC1r8+WlSF6sW4uiB+enYfNHnkgN8onnfdNdw8M0
0nh1biMqdUs+0JtUgJ5G364YYdzOSL8U+1BaCaKC7P/LTWG79E76lme1qUfj9WnZceDKSAXQ0kRE
QtcNOBdCV2RVfajMKnKBet+c15b3N0AewuJod8g7QX7EmB2MXvk7r+tZDX4LicLWLhVWZeY0GRlt
M8t1+Fff7ahu3YuxfrmikT8KYG0Z3S9+McnmfB9xU7d9oWp4auPyuKXr7cW33pvOUiqvrAUXr57K
kEp45HbAJ5S7fLHiKsENiNjgMd0WsYdesU9VFf5bn/pqUuBD53Jc8DO7/klPLZvoSfPytMFhJlxE
PGtWUUDGNRiKgC4hM25kcSGGtAxlKwJu1gbT2b2ESHXMJ5OCOG8ic91TeYq/TaoSaLVTY9aeSPWu
iTD49SbBYWak/KHs7//XNnRiFTrcYPaKZVCqE/eN7DDDjCwdo4rnSGVm6ZIC53+USX2UkdbEDmL9
AM4VbwtkN+e4qf9YsD1c151+aLJ+wSeKM3d/ea7yqUiPnJ/jVRkCcxp9prCvGjEiqSElL65noHFP
vTKniIm0l3tEfGKipfAtdAYcT2ZQyLP2ohKBCcIpG8KmnQNmLjcS2hVb+nKwO6ywBW7sxPRkiNLx
b+cnQfwSosCfavcMlOx/11Uy9fzcIj5UBTGaH0JigeLGPCUoW7KXM6Hi0G13Kn4WMNJLsnsl7Z4S
ioW0PbDN10myPBmmOHmspcOj9zHnVn/zpsr4v/dOX5faOwBjaJm3gWTidVMvB+nT/CowjNTSqZrX
dosgtX1FHuHk40TBxrLk2HXQMmTJJwPBxXbQqYBuEaipaAcoiRK2/ExYFL3GuV98ndmPavkUOtoS
UGsV4wO/SsPDnKc9G99SLoMy/uzx7XpmnFsYa2kdGUN7fqeZkiufwtA8oTmlUxcYpqIDGN7fJ8GG
FnYskqG0BMps4qnptyyvutKbW+HwaFdB8yBYrwjpz7uJX/0cAFt3wQfadBuZKTONQhKu2bYMpX+v
R2fyD8jhyk80OviTIT/XnmfE1I7B4EjZ7sU8L18otC45aDoAJP1iEYDN0mVKRQS2Y7EWuDP1gFsl
WKJZAKLnk2+EMMRu32P5tSj9jy8GdpgwbVrmhQqupOZCNoXw/+UIKL6kp7Y0Nvgb+JoQtSV1G9AQ
uDHzs4k/q6n4oQle8Nm/ZdOnHyrm8+SrQLnN9GM6oTAOPm6uA06ksbNwy/zGcS1jzY6du7XibWGi
9KdEqT/Za07zJdUEqTeR5C8OTl41YMovOYADUDsQ92Trv9bghphsEju2qcJ/ZUs+WCt2Ot8aonkF
CjUEVuFLZACVjBmhOrHYY1fRGdOFaZsZPN5za4igFGTf8p3M70o56ABQOysPatIElZoVUWOdCImN
wmhp0SzDqLngGS/bH16tkM6y6To5fnZxWohgwbLM4WXmNX1D32sgqwT3u3lkICBKJtxnio++OOD5
kHleerIwyR/Z2r8dVOgZxHzhcAIo0AefHpxJR23skQfo1daMmgw6pNGmQ1XWGg/ILhJ5xya00N9Z
79lrmAcJoXYfxq54OIx+o8rLQoZDzcFc10yrao4k+qMtxMApM3Y7u+0Rd8JEszG0QmnSVpQKM4Uf
1dguUIGfV36sENiPHmDN52T7KRmuZQeAnsrSCI5xrTBB9MMoCqlk9Up1clEPwaPTLylYjSKItkE1
otrZiRktlf5PFcABfcfDePD1F++V4DHYQOifPGhl3OOflJ1GYp2ceq5VzkA48hq54qPLwOnzXpX6
3T40yCqf/zR+xP08ZEELvIUqdDiA4l8e+fRHylC84Wj9jc0AQogKjlkbRluAdEoOoexVQat/XShH
i6zfpNYG18apQKQrXxFlAfrhcnjaAKd48ojIDA5mz4nxcPad1eIVMjdmQX45Y4FEr49duNXGErS1
JcB8fza5Nj+JD06aMTCipNkfQZfPHp27FPMIF/ZclUsnjmKw+0/40N5UTvckbm+Tux5NP1YbUjQ2
zU0Gl5XrUeTNGkipLpN9jE/YuSVJ21jzU/6w7OLvcPYLAWXUkn18W3XHv81IfycRHbfrUFwS5Gbi
OkbjbD0Z9URHwrNR5e3kiK3tBl8yLc5AMFn/uHGNFnzzL7E558QPzXA8icTNV9PzevVtFYS637HW
QW+QKaili8xQ+q9XtqHMGAdbtuHrojnxy9MDL6AdQy1BToIGXx8kDGLqVBeB9kfXFQ1ib1uoAVNh
77TCZrr5GJvct/uBIlulerjWZV+0ag/ging4zampYqSLfILd3d2TtRmMYqIgurGij+h4wg1Rrae1
19plqj7nnwgozi1d7MI1EfuwUGAVzJ9DmlRYWgW0bPM4uyrkZd+QC0sU0tqztaDwOXVjURL5KGqT
Vw6juxpkpZKIv3VXKStOIFUPXkqDIjKTzFFuUtSSQTZhpdj6mvIz60KEU1ehvFTSYjDctrOrgUsn
kkxWNEgZm63HhyG3BZcI9cr/cfoMtydq0UiEa0amo65u9wMYN4C8OlWPfwjtdSGA+f9bryq8EOEu
FCS0fFZCYqsl39ETBsR0jjFFxkfoLN5vcyU52qjnC83dEw8HAW5aLhcjytU00eBlc7+E69Ov9zy+
zf5IZvfblORAV9UWz7Rzzqv4OGbYL86bZTiGi6veCun+ds4SZZ+4CfVuX3inMweq+Jqz49KtK8hb
8Fgwy9pj7qW2jsrh+UvlP6R8t81Gn8nVtsEDBIOQSKiPgpPzSRffiyvRaI3aO8d0pDL3SVsLjILw
elnw/P6uXcprR+NXZj8SGg1roAIFj+gjPAChV20lR7XlhfnjKNnd1St990EGqh2nqWOpz2JxagVm
qzqlFvVCzx+Xw4goVeaNoduD4LuTCp9CIJSXrCPON+pdZH+Un0RwJ09iWjMuqAs5mfCQug+GOh/H
HM4rhmsrZ9l4rLWGifOyZgV7F6IKlM27ilyqPsuQsgMy1ErKwH2Ub9XGFLSviyC8jXpXtjPcl+C7
UQ+QFr0T89dVyQFogR+XSUC6E5rKPCHrdQ6YhBRanyHJ3WBT+CB+TBY9i2vaYzsMaGfNNbOa0rnB
5p1fYlmqTb1D7RMMg71DOu7LGn0ismGAqsxC/2/WXtMKhpBBYWmfmSC5IJfJFpj7kjHRKLzXTwXM
FDOSPq9Fb2GUweaTz0Q2QObl2S7zsUHRpbccE2mFXCslpkBRg4lOYMjDB1di+f0/wvbKK4vLtjKu
QzSjPLjwFPGI8d4h9/LMenpeE2VOd345UoCTKB7WQWWRUUJUDkaA2MeFZRe1CDilmblXopOwMj/w
i30wsSAT9IsN835wx6FAwW5ff06H704n8Q6vjKCNuTFFHcbOcUIulwoWcCecawjuO8lanMwadabJ
SqrSOHzQhKqaXKfgfPJbj0rzZ7bstvFSdvGQmHDrJ+9wcXYsweXLMn6cBKhDp6BJ10jMOW/E/H9k
aqwqfI4mLL8tnh6zwvDPEw7bHF31jwvre6Sx2LUrGJsLGMRmX2GLDeUM7NH4VE/twBRqcgGGtmsq
7t98pZyeWJ9/LdJs9Vtqp/WHIr8X1pEWDkEkjj8dcalIQlZn+tRzl01LqvJQBfWYK31SyMl3Dy5y
Oi88LPDyccDOBbhzC1/MH+Qk8QF/n3gMxYIMno6ay/BCgaOnvd6mKQNjNpr+QC5L6Z3chz1O6ZU7
HFKNtKygqyBl6ojWIFbaVMOYbZkVyM8XfeGRovbsSUqou6Gqut1CBGnwaGoST25+yZHdtGTdZCll
0YL2OCEA9NbIefxZYOK55qWN4hAEKcifa/xu0bTDOq5CKVsTq4a+tkXmU5a76A/1z+wi0F/0WzLX
B+50QxQO/8DLBpJM93M2jLTYWH9EVQ+KvsEOp7b9gsvNVIAvw0ZzkF3ms1W2hxl7P3E5DEWl/8rv
4vskPTmLiQmxfOvPxcJcoTOEkAg00Cs/TNURaB4rvkJfokDAVcB8xprbjTbC3sEjtoAJmAU2ih3B
x5OWGcHLgCRWJAI4o8moBtPrgnqfnYASnW06xQyCwu5L83f0C52HgJvRb6MBte2Pm4rwO3Dgw1Md
UB3RE1MvzH9/6RUsSYEoFfzU2WMGxcB5s69FT5fn/eSQZtxzIV1EiRJ4ijI0AE0g2RHX28csRYsi
zq6tBWwNMsQzNghKKYfH5fQeB6Z0QPhm0kU06dTIpnLtMmMRBPmQgXAvR5G4nsH55uvZfeuN4JaU
JTC+wZRP46wb7HdBCGVPFcPjWgbtTmk8FBpyIAbY8CDlVNiwPO2GmEKyZqp9jhARvbZ3tFyIPm6q
PWQJ5riyLj5ObXn9HKEBLBJINxQCTxlLY/pbWo5YPAGgPLEEwFAmrdWNkFbsPBbHredBY4zjglz1
Ghb1gawFwCrVjd0X1P1mhCK8MJApdrwBoSorzYAiayUeCb0g+sgcrFouFi5gHrjtvAyd/oisiCzW
LYL/hCHgZ+sIs9buCo0++/mos+FH7b0Xf/LENJqHcRXnDQ7L5Z5/2L9EkrUDMZ0mEO3Y8aaCLinA
w1iUCUR6XdvUQYER+oYezMc6Ln7d7C3fHz+ilujkBUmGtMuZhKAs3FqcyC/YROwGZHxHj6TzaMFv
twZ45O6N9C7lGC2eGLuzuCPJKmzg3oHoAvSmKrLrpRqMyYO3ixI/npF5IzfZWtkPKPF9+AW8msyz
uKLUmniLhW2LRirSPmSFbdZHO5qLXK0FYqtdj4EmocaVlDgEHk2dT5J9O2oL+TO2oazl+NAWTtk2
D6cPZFkKwMGIW0l5ec7BKOPt/JQgIrdb5NffE66tbHnNcQhCoDZvKRsz178gZ+BLcLqSiVEHTO+r
6GZxprHOdXSQro3T4LxZAVhgTEk9vCZ3629WoVWLCHDXHo8JTboOhZysDcI8XH8bi4r0hGcecXUG
HJYkCGu1Z/fMFAU2o+e/k9KH/J2jrp5n9UMAMuDrXsjwUbSxM1Il3AYEVoPRY8XRFDJVVpOCcFNM
cKnSj9B+0q/au3Gj/d5zaXlEc3jak9N5eky+VWbTrBYj2PnRycQMRqdg5I6RpbDgVrvRL3WJu9mS
dl6P6Rruv5Vy7FMYAeq1rZ3fHrMJ6zPHNeG3Xw1DeHOX7W0f8YghUF4h+eDN3JlmRbjFn00nRAgI
SVwYasSxD1++61xEmxkeidjjhQwiEqCgW2C4O5mZJ1STASii0RcmOn/MVG83qVsIJPoFZuA5pQQY
Vn/NaReeyQFfglxA4QasH/YzpkM98DX9tyYDtHaKj/JkKfalitZwk3nT3ldbpHk9mJwR0UIZ1ONc
PDDtWg4kN9bLd40CIeHiWOw+lr9lXJFW+X07YWNwdnbNFrUP77DrKo++uaYWH/26fAe4xmX0gJp4
R01bYzQ336/wlisueU3BaarqgM7iG7glDhwrhCo2LqvGfpab28Y/ROZ1Lq1bcCvHM48HOiSBOXET
tjhrb1CWhT9yJ8HO2891vxSwvvJ425B03qriAlofTcxJgTgLmluFyklgEZC4SBtfsdlSRDZZABHr
eEkTvMXeA6zgn+VacQ8bOaqy+3gIbT+qKRW4YFMUsNuqwUmOz6z4+yWy3GSCJiFMZwmw7B/7+elB
I1jHHLTr3xKBEVyuSkdpuPx2gu/hHyMZl5h/irwpctal/p0jRtU9Hrm+rCl6YuREDCGAL9yby738
RzVMmDGQ5EV9+sOU/nExyCoGUGW91Fu/X9r2trmBy0Lo01wPOmXjGTHYGW50NCRHn80+TzZx+pDG
b7MauUfwTlGJ63xO74Rx9qLKlNAhujyRyu7DuInar98mXkRp0fGe8nhmWppxZy1nKZL9u+ju1exT
rKBiRtp/BXWv0QfXWpS5TG67NIdTsl9Vj/Lnm9JUKstsM5HifMkHJQ9qkyEc8vI3GKH2kqg+XiYy
O1dYw2a70VUkLPaSuSfE77INcVj9dBxmFhL90BJDpgesYv13MmJ3leAV9mOysutgpzV/S3oXK6HW
i1Om/PMimiYvOQqeGX+bp26TJApCr8F6ex6zd2AcpF96ggrgvV0Z2cOkslsvE+uDG+5eIXWyO7Ei
Yvsp80TFe2q2uAx2o2+Vhxy96/q9R8TtxsxF18oUE+FXJCsexs+E7F9y4Yl3XHPLaKD8cCken0bH
/GskoPr64QXUC3utvOokOXO3ZhKlf2YhYaPVEsZ1osQudRDHMeuV7eeIpn3+XSA54GApq3V3Y7g9
arpDljfQEmMYNVlm3mERJg8QPMJBwHA412TeCfkSCeu77qgGB5ytchu+mPX+7ZaGegzpkI53pBpf
O3rzdY3SnP2JP9SvnOJd3yNv9uXdx6BBvjqAr1Zbti6z8eguFTvBXtwibfikuRG3+ZRm+B2zPH1Y
G98PYpUgAsTqbYDLDVf1WABnq1fr14HPdGTLWc3/hcSwpg8opVYA5iI7+LTWdomozWisBip3q+0P
7O/665Pi4iaO7n5w7CcqHl1e0vobCucCKY+AMn6ZJXjoQPzDSFusVXoLfhas8aa2znGXS6hurIZ7
ZVm1mzOJ2zKjsjjBTC+evcR+gafT0ubJdkJS3aC4VckYAc5QWZhZU7et+/nC7X/0n8tEO0/ZGOXc
4bpt9hLMUj07aKB90PTCa0eOaklJRloAhRtg/zcs4nJY+NSL2TrKw510d4SaG23h3o5FAzxY1OCT
aBn7nPiJY3mQvmCyHrnj0TBXUTZQ6QEosyllePWuC2uolxUtt2I20+DtLgdV5DTMm2UxfEhwMSmd
bhJJ35BxW+thoAiF3iA1SXVfou0lZiZ4MBFLmv4HRswdqCgcS2XHo175HkiU9L6BAfg8lvCjBkAQ
zniHHD0gKGVkoA0AoGr81ueoiUcTnaJjJSmwMaPuZLR5JsjG13fO//YhrjNQuzRyyTC3fDWwSPWL
kPawAgSd8B4guDcb3fiR0vZLa8vNHlnCVKB+3HdWf913G1A4Oc/F96JTkCHyFsifwyi2RbcTxgAb
JE0r/Fh/vEi2AFTgoPlH4l7uSf45vb9ozE2YGPQwfVgfHnym93M4Uof9/s2feQGEASbYul7Rim7Z
NmpN4ssGyAvl30vGoJgqWcrQfkTZbHbSLNdcRshINS81GdCbKyLjsSLkH9+9K5ebWaA4CukGocK9
YJXfHqre9pAy18gqvSSC3TsDodrkx94NQSpfPWkJl+mirf76uFnSnMlRsgzCCx9AmboX90Mjimn0
8mqkWWmyBE7EGQ7qkXX8S6yMm+4k0NqNBpS4WJTzhxIRkBcOZLh5bWdxwcMf14kfqnJS/W1r9dFM
zQ/nkpw0f+6hyhilxauh/DsrAtTOdfb/EVMq1s3wbS3myjWXfd7EyP/+RqusmTk/xjZoGqknERwP
9dz0wlNZgVTSqt/rG2AbqBmd3yOGOzKZ4spaMpVcT4POaH93yU5BZHSC60UCRJHshbT//wg9Iy1t
GB0COguGwczooqCl/1wmTYgqhtOsQrFm9fAFr1nEfltNKCfhjwSdEaKcXbWkPmA6+D4KrADw72YM
i5JBs5cQvcOsTScjVU+6U1dfprC3UZFtfl+MROh+VAqDQhvRerJ5N66yUrOAKDx3pT9toh8LEgh6
quk1+NflX12n+r8rbhCQ25oyaf/+3UF4ImicI4AiwoHiJEYpU88kAN5pTO/Gjpcarx9WPGWBREx+
+3JUt6FGKVLQ2yoeygrxwVzOQNFtuEg7JUFegAR+8RDc0N+vl6g1NwKxWrckaaLtqJ637XwLTWGk
Hpmm9Mc7wRMBRCUZY40pync1BDOfAUaHb5sfpErT2wMOBgpaUd4NpogkAHmMznzin1HME0oVz5t/
TTTXDaxs3hM3KwddKZtswYT+c2L1aWhPpU9lSsvgfQzg2CY93x9zoEh2fnVrR3SPgYNH4yZCLkLQ
DBgLraVX8qTxWfYlXqVh2759N/Rv103LKc58EafPi7K/6I9/5UAOxAsOUboxzrBhzV0qpxN+K3MR
zO1vz97eyqE3P6p1jw/IE25wDSr7dNoqE0kbErz1P6CWtkZE3Ub57KjXTh7NvQWtrgx1WCszuoph
ISbZpANYKNQNmYWlw0IRMqIFskup/mC1rbv6UbU2WPX/UMs6ln3yMSPsH4VwVsRppDJVzEOYZ68w
+YZ6/YRRhSWqgGOrXF7twF+ITzwZdzGw+btsmSHkbVyvqoiL+LGzBveCttIKFny4Mj7/puhbQ4ho
r7VQN9sirq25TIl696DRjaTcK5gIzMrUKY/DpKMJW8kRlZoRfStlKE62NYoKBFH4Lpg7sD92LI6d
4uMLcO/csOePFyifTnWOzddHodyG8CzDOTQvzYmFiDrTKUgoNKZGTk2iJuzkFS1W61YiYXW9uCEa
fKOdzYNbmIoKHQm5xom6froXqFK6hOs2wncFgvBwkyLdkg81i5fpHHNm+u3fEW+1Xvva51KoiUbN
9IoljwCOeqtM7DBuCo+jq0OyTxrd5rkbrdXf+SOJoayEV1ZZ6z4vfuxb2O5X+cPeXLZcRcvORbK+
hY7rwagkSdnx+zf4TEeh/Ngvq+uoo/fRTa3aKnXqd2GVG6AVrcb+lUWtqC6CeorKu9J4m1W4B4G8
nAbZd3RdgMRO0itqOvjWf5fU/g7g/S8lEXXU0b9UZ7Hx3bQXoFihgAY5OK2HB0YpKp3K86d9y85x
kJkCb/mGFxwkiAFcVqMF1f/jiZMKEislT4Frq4exWOCoc8+gNExQVSaRjxG0eeELRl6N1pcrQ4la
BmNrLWtwy0uhLId0/l6PvNSdW8uOJ1GXLv7ZSoTkkTB+AOuhefT+6Hvcz+cMHC3bUExRBEUDEDjK
BbVIXqQnlUtiTXnPWelBHwlSQEQkLtygzgJaaAg0WVO4OgxPtbRs2DrCPeFs+Uc4c9TKUrk2oh69
AoTxWfS4FEvRg1U/TaY3PF66mBxkYr9dphGCRS+M7ABdfM2l0TanXru19JJYEPpWb/Hbjd2Djzy1
Lo+mxjwXuK4A8VEN5WjrvWtnizIt4H4oVMcdmxGf8JzbLZ0s5EXZvhF8yC1Fq5VHMs6zY8Gn1ukK
5VpfESZWMTIaoqR9EyJm5ArYnvjokn4PgCzywqpj51m6GdswHIyyZ9lqKrjtDQgMuI3k7D3N9Lhy
qmpSi65MRbKzvbACTlLh4zxsMWJYcF/kXuwCHcUourpzhpnILAqonL5HDKGdVryVurE8Ixu6w3bA
VYPQhGSlwkRzw3aJcyVOQcnyzMupW0M27Au4OIIz3o2ZMedK7khD8lpi8GyCoPTmu2fWxLNJUbyS
/+8xikg0HKQzyl8QW3fsRfbp5WpcEEVkU3zpJP0g2m4aP1F0XtRjTiGKOeRlMtQpRYgcPQzTtOag
WlyHPykoKTU8fW7cCwBk98yfWOJcr8wMyyC9PznwNw23a20n6CGGQB5OXYB26ULW5zFBOQiCpmeL
5tfGGkJW26bSoELGy9hJPVVTGGyly5Q4OUUS+E+tM3ghPSeZ5EY/p9IYl1xEpeLQKRLHjJeO61NH
9V+VGIcGer4pcxb2xP3ngVhHHsnYt18iitHDfg92IACValBIn8fJJOQsMQKrXhWepMCr3l5bqb8V
me1+IuE7uAN5dxXJlq5d17TWo6UeparuEwMOgOaAa7yhUerI5ZKYCjAg+CfrTtAF65lR2UnGglSk
qKkUpoOYJBEosSF5wWgb+H4zk1zG8k7V3NrxjXunzHnYwxD89khiVmV0bXaJNHpgpV1Pgs4Hg3Zt
p8GiaZCdxGWg3z++lHsGDxsYTdnW9RAqF5SQS2drgnqEa3WC5AFCDT+BWmqbgTow67UI6WbG8El5
d2m0kqhJCWLwvNod85jFaUo7vzE/3yRJTIhE+yQlLZ61EqU59qpPFGfXdvYx/0zGhzNFrPwG4mT/
K43GtacrUyQGlq2DZh27x2HQ47eo3CHrWAFbNdFxi9FwTc5n2NmNv+egvI9yUwwiIG2T+eDUSuxd
2gelEn9dqQi7+6XPUDrDPnpJMsnjmBuHGsb/TPL56/AuqGrJ3uxfl1equqccTNU7QHeCmdEnSfFg
+Aap9tWlZiQYrEB1j9LEC9ZVz18Vjx6KaTXdZQ4rLgLOItpt6kj9Si5WRH5PgENtgNqio4cgUcPV
AL9fzoIf3W9s2KEyu2qpk7yMLgDg36NVdvm4uiWf3CJaoM/jF7StdEsJGgBv2g0vPp3lfBmvMhYA
TAJxZNsGjBPO3JNw+pimsPqmz5tXuBVpWy3gT0msMu4oFJSVNh+SR6JvmMsNQS42BxTXMGLp9tK5
jJjEgELdo1yXJZm2XwmFrOMziG4jeqN/PLihQQJUJcn3pDYYQlOnltD2E+haH3SV+hqw0K8r7tGM
LeIjAoHkzgd07h+BPjK0HJ89aWpDbXJAZM3BWjLvUasy8yPY9XT+rXZUaLtRzubOhdjDaJ2EMa3F
9wptt24LGHN58V58F04NFlDWeU1Xh237wlxsZsqMknlIdnYAamS7I/1nqR5Nm22UkHw/NrTUG+K0
Q7YtgTKIOHj2ibNve0axnDKQ4N5CYZR8vBUsNTlKMc/dHY9b9FXJUXtjbXcVZQhRo6MEsNisAPuc
3NEbwrKptk5sGfMDV5964cW2BMqnxQgfnV/DhVvqYlEZrINXWf439W8dlF9etN2ZbiT9DKxXgSyr
BRxRtRFl8Sh1NsFQitikIO2TUgdmYtp8mrir3Bku3EdoyIbYgHfT/Fet7VX9e7oDE6/Nj2G0XHsx
JqznYyRrEWsLfSLLTsQg65ToVUzF9niBBzP2y+YAPLAzqnEfdFqFcmWS5uPMDAl8UasI3FbcMQXw
Ox4Dr4yBgqt/4rVfFCq0TtJREc2hs0bpJaCbLeO4gmkCaZGELlxsEn4LDAAs4kKRtEvNjOShUIEL
sCCk53tayVFRKsmNghvAFlhXUiuv8WgKzC5nRNdrlt/S6VxiX3YRU+TbcXPOR98kmQAjJslJjzE9
9I7OE0Sw/WkWSH+nEM162MV2ZWMV09A4vzTO/QKGEP1WMfKg0mELj6Wr8LoabwU/bJ7QL+CjMgq/
avp0lHcU+tC+Wdy4IDUSFbedvvhsSwn+vOA3tImeqqY83qTBncWUxaytRSOSHb7Js+nRtvNbBWsM
EN9yERB5Vm8L2c0SwZoOwoVF7frqq5wy2661DII0hpUlpSQYhdIRzEWyKd6vQgxikRkyLOcGtxlL
e5GcNsDS2pAhNZXCyO7GZgv7Xuj2cjtlz1pHD5ErPhpEC4EBGkMp/1QgQT9OwWm7IDm8MhdVceSf
W6WIMLiY8iEwbFFqcEcSYq4lMgKVhU8lW+TprMkknlAleP4LoSSYJILj1QBF8pKvR1HqyQZbFXPq
5Q9BdMBAeEFbbmszKUiLurur9VhK7bXCnTRsNovp0J/VRO6Ibgs1qRY+AexVbqxH8lAeILm3OMDV
W8N7zzNErRzh9tm+W10ScWKJcGsZWHdvqiZzZ461VMgQ5EzZxGXwYN+9hlePWRsvLIJIk0ZhN8Su
U8Yju5fr4BljGZb1+m//rI1a/b5z65vs8lYG0XDTaRlUHUOQEWwAZYhU32BYgQOglqKRkeyZVBFx
JFTtnc1lra936WIFs4v73djb9oisb8VLbneINPoFJRFu+3vKpYiqyptoiGFDo7uJaTKINxIf0eEW
6wMnEiLhznTwtbTnuj3Qph6wjN0Haq6Yls135zQcsxBSro49ckh7z4PrwMbcznbgk5y4GTCNoVgp
VcqILbXPc22hvoW7FbO+9nRbV2UB0NO3Azjg4NcKHdOfbWyVEW65d2wanbxkWRrQJhZaEXKQ/nY8
NIIeOAUfZZ1JFky8fYc5dP4ufIOMNy1QXYVCO5ULaw9PLQbps8Jh6adxIed1EPb8gnBjO7eEDgj6
gircC+gBFnHem94dfqsiKxVCd0Rn0Jo3q/EF5Y5xVS1h7gu3Nwu3Uh6ViSlxHNwlWKBkie+ZjcEj
Q4GGKTmxouz1qFdb55jxLe1ormcfBh5ryFufKX+LEjU7EKFaZqCGQsDHXoP9Up7O3zm8a+DWvLbC
KhhIrixw663sAeIpL10UxjOSuyhs42S3QZ+dTu3RneURE4oeM8mlQdoXZerxZ0R/9ygc91FxH9vb
RUjNEREjKSh66UH1XPwQ/dGUXg5heAnv121qU4VKfK6qkmH5nSi+oruOruHQIMbnzfojIJvySVUv
tzpplW+4z9GMay8hmkXylNszm4jB7+ZDGWVMnbZYB+AAf91AucraQM0Q5OnvsnCgu82EBLb3WfR8
fYbTT+ScmgujdaA+asKJNe77QdGV+9+76EURAx5otkaJvDxw37edrqd0KHS/6pkrufhKfh1m7oeQ
3PR5NV6n07F5SK6IqELNW5Ohko7tNoSyeqAvMIORSAbVhzzvwlNBVnbZ9ztCs64Y6hS2058nHYaV
XbMBEBK8RkrPaXwqqybaES6qoj21NwxC0lHHSCHmH6R8NxLHeJUrHlA+t+0T8YgNq3CETo8BjfZQ
cNq+f1AoruNtuwVVBLHXk21X9qfyNJ42ocewOIL3smOoO6wiZ6uIZVSMEsGSk4bFzfWaAz7sibRC
8AZSdRPyytByits4HpfeXvbDSZsqt61kmKp3+agmmCq/K1B71gSCWioSEbOFxLyXa1Ha1qXJZhXD
SfAUdqLa+LQYpLKFbBMCTyMBFYIDqP4bl4Dahv9UkjjViMaUTx2cKzNLaHd+QePjGEhtH0DXBl61
7jCR6im0whVkwGjC+6pvRbpEHFGEvwLgBIZ5IgnjKeaWSqp9IhoyOmA3Lq7n8121e79t8HczDCuX
aX/LWY1ISndNIsE+W4KpiBOCtnN/LS7Q3xIGLdoqWsMoC2esLnav8pSYI4FMdTsmCowfMoDlI0Mg
cdJNHJTMuaoVTV2ei5L81QVbSUNPg///4d0+H6DFhFH1EKD1AZDjJKV7HY2YBguQW74UtwAOUMg+
HRknLJ9040kcYJjgB/rWiZv6mv2+wdL+LStTf/mJXuQcLKmPSI8zlt6mD5z+yiTcHO1ssii/5GQA
q6IrAWSYQ3xfsJc1y8bs1Q5rpsPnL4UYVNj1C1UMXab3tskpNngz6atNcqWPg4eYsGbwo1Avr76j
Z0o7xBHnQlDC8xC+Tkq8qDqJv3T2jn4x/MSX39M+vh1YwqxAtaSKNDUOePJG2rSzWicwCkZmG9s6
VOKPURzF2E4H4Dc4iJ/us84q+ZaiUPs30MM8Uxauvy0at4b6qhCb7WYBDJ3WMU8eDqoSr1Cm8jCJ
IPl8SiwOZdIOtNmZA5U2B8fdIHOxEM0ooddq5RPnfw/VimVabiH/nD9zqpvT665sitQpkZUuKWwV
VO1svyrPMeut1yYYomtRH2S9no5Sm/WQYcEfhbwK3VqhDxq+sWDs+rhX3tN+rsjct9gFzw5eLm+s
30J3jYvPbllDSz44pw0Dznfz7ukhcjhis+qdGmn9jlHKUOwHjmuM8WLM6fjO+c7EAwsQsa5NEsru
HGZAiRXtIIsfXN1p+vnFhZZwqt3QQ5PdvBjlGjdaQ6X7/GPLfEeBoXBeqwOanDuuSkbULmJmDiDe
VuzUvtIJvO7Gz1EiZENudMxhA0vSjcnxoSvrJ+2IbeTWcC0FPLaJ1mdVq31RlyHNgP5vszYO5Am8
cb3pMRNuisUqCBic+GlkV/aJx/64HZeFVViMFzMeYrZftGKQRd3k4mYFjsawUFTSpe71L5td9O87
dZkvgpzlpUZiY7rMPR0JEkCJ3MARF3Jy9KeLjNClAUQHl7C4UTPFVwVmKZgFQx488qzKEVvZFd3E
h2dq31/+TvY2BGS6DEdz3jA6bOLW7pQ0xwwumefsFIlGiZQD+p+nxh3lMZ8jwKy4LsE6apRzORrI
miasJZGOEjojJVceZ/Mu+zHGxeywiqGt4zdO1+vxGEAOj1hihKsQn1dRPARiWccfW6e1fs445KoB
HXVyIqbSmOrUeOXDLTnXvETmr9gVBeva/L1ph0wvYn5t5PvnzjHUSN7PYMJkoUHtBEpYo76Bt3bz
mdKLUDOdLLVpADwslbEJ3bBxVpNO93cmOZg9rfYHb/juN0NHJZ0fo+Web+fe7YR667seM5mjQN8R
MNjmfYfNiRvUXGIfz7/ie6pCTOP51ipvUu/aralXI270WQG7VuLp9A6F4GSsOyKuA0J0+R42qlFN
zZ5TvTNO6DJDmYzKGNQzgmk83xN21LSlrtdLS53AB5r10xxYMExWulj9INzRgcUPA1NrU9ZRqkSp
M9cByPaYW14EmG2ivbEcKsBINh5hqGanqmaeLinCZMFVOwbETKli7DoOyJLVpHuzsthso7xynY5O
rqfX3MNaHmjXJqdKLKRRXhX0ICunQcW97faljgVp0k1b77pAqCzcwQmnrVvmOaLqa2xskJtpGFCy
KDBY7BPujuHC/drowXzLPITmXMRG6i/AzN51RDR5jxuWpW0MuGeqdHkYVJdCxJbEN8vkwJEGBjW7
kg9bOZZ4J+B0QZb7J1PFN0pNnRiRPButZ9JVPzEx7w8qP4JAy/FDARSvc0e2Syr49LyFK5s2WQlp
t+fNIQkHeGN5oD8m/NJd4GKA9EJ0eutuW5+OtBRkKagXIfTBaG6huk6Lgy0A7kh1c22BdDXJfIXJ
Klw+6NjDbKWexBd/4pZj2wJu6FkFXio3ndae2vKhRwaMXocxm8y8vBx70zDLFRZ0jPTx9EsJ0Ch5
yEYxz12E++XMXOje1cxx5cAoaNJnqL8cMxUM7E75eJLnPD7JwNBaIVjDW0VGCCSb0+LGPrxyYL/Z
RUTXFxb6CzNicNEaKCydAGaSkIWnqJ9YHEL7A3ftnznOCoGdkP59kiQWJAbZqIMG8NveBrm8Qqyq
tISjLTpmcYGlDD+nEuRuO/EP9iyTMU50ux0YGvn3fYrb36kWcxo/t1Zp9y/6FZ3AZxLplURMmLbm
/iU3v3+yxXjMsLiD7qQ5UFgmcUjTk09uaacie/rrp5GDXU6ld2X/z2YXzSiOoWnoL+8P4xKIAFnz
IQ2NyUHve59ejM6/cd1f95Ituij9B1IDHH+k3leszY8S1Px3b4WGVBR36wiHIOfSwJrE8iDXS3xD
XAT6RLXVckdkWiM4twLjUAmsQ+2hOQmOACvIQtDTuVIFG4FIS7qLfoa+DttJBNmIX3JeV4mdq7n2
TSef1f/cdioHT1RhCRlUjRdmwSYuBVyeQoQSPiKfCy9YjWxQl44mvuhk4nogH6NS1Pl9aTdzDHQ4
BeX5mOxiv56GmVD5IG/V5P1YQi4hn7uJ3Hq9YzO+SL7zrGggRd4kJ4pntNMTZmDsLXQ/kYlc0PLP
6a0HLF+aYrYV9WIQ7+YSEg+hNtGkeklFNfi8UGbVhOuRZLi0bMCzfJVMJN8SZwwFQ3rBU7nKUt/2
SX0rcxISyWCnh3hg5oSO7X6xpSDeUAuzVJcPcS+wnv04t+rwJpxjWfKPu0JJVdarPrjGqAOoZN67
ymZ+fddhTczq9+4oJjU1yuv88Xc8VbUCLqJThZX5K6pAKrHLVt/bb+xzMIjAAP1iathEjKETCfoK
a3lph6t8buY0D4LwTWlHayrGA46vscWE8ARKQ9+9ypiYjFBnxnXQ6IafQj6H68VPOKNT01u3U5Ex
dTVdj8V+mviFBEqaDt2q7/eiiD7vQnlFwOjdUtZmXq2rsuf37uh7W7apOZHl+hhfkl7FsWv1gGFp
DdVFdZ4XItrCJHkdGT6uFxYQ7hpRRAevDTu/VapO1EfIQDwhnzy2gFtkVtPDreC0aEx1g2x7gUEj
T/W3nOC5iv8kWN+6Nzuw+rOCDtu78CoA8t8OtALHJLl5UDhWnD31ZZGB1p18/xmspDvA6sHPzGvp
9vg6FoHog3v1XA31K1/VAGu+AsaO3SSpxEKJ3gqDDaYKlplzemgzEWxAfOK4DfCPfeA2fBJmTuVP
HojHP9QH60p0oMilSkysUTEvgxOjuS8dYpth7wB7m7cZc6+62RK0fxeAaY2LZo29Qri0bm+3NjIi
NTkiM5PFB1oz9yAw1rynDQAUxZKV/VlX+613tIfEUehHjpuXihXVGgSOzw5e41WGBdsCm58ycrUE
Y7+LmXuZ21/E7UdXKWwUig2a2eWYXpKyY1bin7q1b+d/QsfBddyNXOtfmVWqVIBI9WvzjJf0Fp0k
NwEkbPjeMzlSt6lestTXI3dIf6lgb5T/Hfd301qKaCmL8cjESXk6unKZaaGnTcMVAG2GFqL2j54u
aEHUrfSM0OWxdaPIFkecZ/bsJjTBqFkFDokPEvN2ZIgjqjkey1DCjhjzknIVndajE2psD4Xh+RPt
LKys2+fbxNWckfpcs7GjwIkwmvrJ9ydtZaCFjyFZMB3r51jS0re7bAE3XL7QFU5bLMdCCBV6Cn8E
xCxMfqigRSsGisEq8mPNqteiWMNvoFtS1iOBIuoG8r9OmTpaQXmHzyawYTIIu2MIOkOsXpyxLFi8
DxlCnMJm6RlpwSLJ30nbiOWDiijCqSimIvlqg9gUwFg5Rqe57cP0QMd3dwFUO0//RnvV+34y7iCj
iEmY/fJOxsd8NWT7R0JWr1ggR+p/tuV0wxAWN71SV+A/2AMq28rg8ZQ30n/vZQTIQd/Q1CN4r6aQ
r/23GCgL2KDttxyI4gM/U0ic/q50xzXa5Px5uCSCFtkVqOsG1imGCJS8A2Fmvmr0JNthrcpgAEg4
wV28iqGubTanQfROPF6Q2l/sbNQyVYBDOdjUSMSg/AMe01NXSExq2BcNxR6zt3bmOKiVeAcQi349
IoCjwza1HsgV+X7bggva8VKu3Gn49v8U64VJ8FtJYZ9UeMGOifkokYwU8k6bYNcAkDEOs8az/faf
BF8ddVQHU8O72KHYbL+d9mgy2BhKKlIMDeLeh266Un78y5q5p9F6FKzmSkdlH+aigaUDjVHQmSRS
VcepZRavl2G7zKhOPCnhaQRPFR1v/Mwq/MIaAbIJVNjCDRgrmm18ypd0e3s3bniUinejUerkt6S+
LChTQB3N3BnUe3OCAT6k21XcJokHl69Z+iTCzJfwy81pEpCqaG1Tciai1COUROSDknJYoR9FSbGk
tXL1HMWM5AiTDAtLE1RLQyh0m07lVG1Ikf38pTLAAFIG1gTMmHASabkzlksLTh2GzWXIeBTgsyYp
lVD5Zhr6RhCWQAPAO2TPgavmSBtLiM++9XMaLm4LYDYrmWipTJTIu2THDTNQCJSjQovTsikW+Y4M
yuigsx6JOb57AAL0gyNI0zsyDF344ycSW6UNFdbrQ6BjWRIjEN1xQLV5Ui4nG7bPgUNoHKaBhdt5
JvRC0LjqppW9uj6ByBIGjICXvIqXtR7yK8H+4IRsljrhpo21S1WoSk9urr2c4w9wCyOIG6hmz0ns
CVbbaqL2wWSiRp7ugyxcD7vxrqJKnRaby1Vch/GRx75CTLJKo6xrLWxHmELdH5vewX7rZq1YGerM
Lk4Qh4EKWOf/Py+/8oYgoIFOrD8J4Ip95GF5aec/K+SOe4n1M3KlBVTrTC6YTUHK9s6jOo9N2yLS
6J6I9TzCYUT2Ar9nnIaSKFmWY2wO9tRlZNTQ7A3ouPmS6XliwB5/4U/RJiCGgbpgnQYLSckE7u7v
TWK4oTDJjdphi8THfELtTO3B8ysjMA5PC1DCFpcG5C40IJdoFu+MTWwU6dBbcNaFAyok1YVMttvr
1Dd83KwhJMdvJPFOEzEEjKTxdPy0tdiIcx2iWnTwCmLbZyB84/1cFqGHGHuyV8rpPPTmiafA254P
LM5+6rqF5nH8QzpJKQx86ujxYBCLNDeWni+C585nuhmDEt0tV5wTqURhOg+BwBUQaDnGrqmyyUFm
f/E4USFBtu3wRpPKDpoCF4pVS/ESMkjCMij4+Q6aefGmyvk+lubbpou8mY+AnCtUYg+kD5CmNLco
Ej1xODsSwjEgZpP6EjJoP8OH6d76aL/i9yFzEvtQoYkzIwEXfUbEioldzSrpQXnd/oYKMGr9ZzNH
ilMjgEzGIUDPAjJPGn8UAjKjMnOOaQRRPcIOpKFQGIuV/bpEwHW0zZFtAIkgfRLoQh+Rz6KNRBYd
9yNxlEe4gzSSsR6Xc/Ott0B8rriWsI6T4uSgt4ym1BUXJ55BcnHZz3bNKFGcxU2KuUA46PQyHXgx
gnGtggGWKJrfAMPs9IqEy5evnTamBF0mgxfbmADYbf467QbP2lyzkH2Y05bAHnMaUgGwrMzXqEax
UBmCS3dIk13vFwe0hJDIyjqZj2goxnPlm+I3Ah7FS7ST1v/TpzAkrIsusevnz6Cke/h9dR50TK3C
GwK7n8claW1iZu7dymq6/yF+JY+UhZPvJeBdjbvZqL2oiR/Fqhpkls7bSa7h/y3JwrksXvinK3Ty
s4zpuMERwRoV/wB7blL5O6R+f9zZNbyDUps1z9paU8x5KvadVqW0S3CPj0LuynGEhUGUhv+gIClP
JalP/hZeARx/PkSyxEd84HLPBDauCsd7rG5dNC9FwI5Kxfil1cgXdqDof5/ZWvGZ1/N+nCjcNS+D
9SRO0LBZkudQ2j5pgFqgs/XUq8ZClZfRiSeQbs3uwC+cBlj0mbuULWhNpVuLJun7xYfeJpXGxebZ
Rpba4tjMz8CTIx9pVHD9jgTgvey7Twq4c2Kvo8aRtxKie/FSz6AZbQuxMrVv9QbV2vDH0PonqpTX
5l77oN/LIE3qmav+M9KaIQudf7qAUXrfpprKbGMIzXVOZpLtZ0W/e4dv/dFJXm25YZhGVgHxn1Yk
FLYWepEz/l+CkBSBxE2b4zEngh3c8E8bM7mOvB9+5bUC71Z2gXEne3HzbDY+OZArxJKR0uBw7za6
glGWcfkbzbzN5lJH6Fy9VsTMdL10ihkavYVidaozkvVnJFViyBlQBLI4mxG/SATd2EQZKD279e85
Jr4kCE1dMQp0ILbFeDfA3aW04giA8JXvVvl6ge9pZ6IhNSA3MN1i+jzZmpKcy/IfaHIOymPcq9DY
dPeGrzUq+hqVwktERSQ0ERLjPnyo6fWL2XeuAxBFGAz3MZrlkygP0P3vl6rcCOo+PA6OvnozQEr+
i7ER2r9mfhry7/qgTCpfDNW2nqV2chksT4X7WWFBBz/n9vQGOZzFNCbLb07dBxd8/llBoDlH4mk9
5tvXm+gemXyypY/vZGKxDZHBwSJPax+EbuXTO2bDuqBnpUxg//nggND1kk7Hy2X5AvedWtjCzFAO
5xVcUYKunA1m6zYO2nR94sAo3n7ZpXVcEFCFO3qn5bgZlX2e2ywJm0rbK1UFrrJP0kDv+QKLZhd1
qSrY3W4/fY86io2ttVg24cVZkBUHkquX1BEvW5UWUdB3TIIbqkHgO4RfF5Q2R4c9fi+3M4aTK3Mc
DkYvibCHolif2FC44FQqyNaUvCgXNxoD8335bZGGG7eb7lbKKIQg/cz375meR1bAgvtBlYuEZ/39
olPfewU+KIBAHY85NxAekNbHO870/T88zQkacQfUu2SM963ID/E6N3k9Go00g5RtVT845We6tMh8
cPNG8572spkizjH4KWT/D3uTeimcQkcdLmreeIQpEKy/UI6fC3W1qYqRANjDwOduVFzZrUeYHZ5W
sN0NT8ffKD6XmDbgGifaPPk+bj8t6ziWMQQe5EX5OH1WdT/79/nNxay+/cwSD5nsAGcDInUab+lU
QptyX99HP6455TCYDTJWo2tJDSmwwo0V3rbcsbbor3r+aYwNYw/7XOrbAKqM3/HQFexvXnkBHvJW
Vat4CBAd+D0B7/rpaHwXArij9I0UImuUruF+W0se36b0uQV1Mqc40+zh5cbRAQ/H0QmA3lEDSyJx
i5XFk4RGGyW75w/r4IeWVYFFYmlo1c2WYUqyaNZG3SFAQa8YjMNOg5G8HuRvhfHqrfzjYG6QqZsn
vplnZvG0YYspKBcaHLrZ3VY8khr6k4AwA1uOBu46O0WdDchqdAHLYtGyMIS7GbupTIQfZ/EC7qbA
ZXEPaCOkz8WPS2cVwwEFAOdK1ItateNspp+Hnre80QWjUfaMKCx/n5Gyjig0SdJP7Zdw9EbRjhAO
Fm4if8kzu0ub3BUGwKaIPWQ/NeNXwFx7I6mgrmQVFNoeZWkD/sciQpo9MIL4QS4rE92P1K1PUu3u
yRNmK3cH36rVgvxPIYfqpJ1fPMbJWh0zcCdJ4HetnXGa7Jjf0Qt0qeewHKmYxKSv2UkBVdOp6lbI
oabUj6mE2J6oneq9g8suJqQ4BhysYXmS5dFTUHgXrDYnK1GbXK/Le2wHATe1CoYMrmLEPUwvvAP6
UBlkZOTHL6nrh8YB6WUF9Fw1nPVSuaAGOsnCQFZwuDuCX0cpgcMN/IjZFzpgrPZJRRuatdhY8Q+W
MItBGk2du5kqLkLNLBnk+MR3e5JGE1QyDNyKYRH2UCcBqpTm45fXgTjcD7vhipyejFGkBzaLYzwj
NR+mhK907w0gDZoBqvugvb3UefQQm1VhGrtw+yb2qJ1BDW3NovUnuQ+JTIL5X6+mKAJH+hnaUyjh
gvfkZ3hoWUs2DW5wsanYxp+c5EKSnRjUoHQGE+sX9J2tWiStRTebf02Sr0767IYOtmAYP9Su41jo
KqHRcL0CWExVOYMN0hjfLRacQD/ZwzP2xULcOeWA4MeUmkSqHWVDDPIFDJPVbccm6ZJxLmRRsxAR
nSZxCgdXL/ttEWMQDfQLlJmE/LneTkgvwGS7TpemZYHNXYjA7arIfCy+GWe+LqL6O+BHdjvn8IxQ
Gt0c+PD2G037UNnbr6Ie3lKszVUJ/9/aYK4BBBsNohZptksAhZsuxQ9u2MDeP2RNPlJmCt0UMGzX
xlmBDaHTNKTG7SH2U4bd5l1TVdJ4aJ9qq4BqAj84k6g7Jl7FaKdkR7V0wWP+VRU8PZVWgFKPXZ5V
2aYhdVu974ZAai93z84yn/KFR3nhUAZcENEAmPpb64ZuEIJDdM5TZIdnnFXbYmlk6sP6zUZG9xZl
trGivgU4meHXYsjts0DRUV0lJvfm0dyA5KSK/Z3fCmBqUmUxLNsAGIHipiP3BrIg4uwWo+Fc759h
UGGQwsf4Zw+32rYJVdPSQhpzSPBu9MQEWJ53OjE//LDkvxRS+wtqmISXaxzxk4Dwmwyu5CfkvXHA
SIksDZPq3RvAajkFx5M6lsJGrPuBj+TaaurZ0lLSMHCv3XvyaBRQazJxzjtXzikc3Cf8x2lg3Gkq
XKUxkMp22+ji4IZuwNXYfqAKVGHSD8e9z6B/+5whZLleiW47+b4g0/h/LTZPwioSK42Dp/ODcZFz
PIxfXC+4cc6JPjHP3Ry2x+wF/VlBf9a13dDZ4HrHPEnJBVTPc8MjB2iMlwfsudXVlr2q0tZw7aXF
oUZD7v41RiOoFb+dPTH39oX7ahXRCjYm+2N+pF2ZE2n/LxIlAi9CVOLxcAG8DDTCGfSqmbetAlBL
5A2TUd09nLXegpeh9VfY8uPQr00wxH22I/dOfHOJDFv3KdEk4uig3EZjz0j5Mc1jge7l2gh5S215
d8WLQrKYsJUpp4ubSZz4DLr5DTsqKj9O+CUq9PdpK+N2LFn8MvuAalD8PITKNMbaR3ep1dYA7PYX
QhLfE6Vcxk4S5IjdeiqeOt201tTU4PJLe57A5ZkkVB/atOiIokYLkp7uKJsVuxQq5BnTXV1X9TPj
evfQcW9w8UNEsJ7A9zs+XCiSid3yLAuk4PaffszMk9vcRWZ11ZYtzwrM+WEOtUFIoeJ3I6vQ/cRa
wSFgd7UbpUtF0PMsad3stoWarpNOFfWS3G7Eh2Cip/PKVVEq8g2mruJ0iDRoqxDcoIsU2CKmkvAD
MyraXC+iZzFOoNREC9oZQDSMkBp9bgzzKCtBrghZ6fBZs3M4I9nJIvlCtWSaiaB9UIhUpBb88fpP
H9KjedHfoMxnYMIHGlVOMeQEzAUmDkH4AQ3ukC/9HkJYgjdr5euxVLbRntxjBrPIapaAoZzi0/KU
1azCI67FD+us2xPjEeemLTPxsuQgl5qpFfNdPC+gMR4GUz73gg+7J98Gy0Ns8zTOuqs5NCkphIUD
wS80tCrNMjGqCN5xpiAMCFl+29k8vgwtURybCoL3Vdf8OiNk0/VWWB+0o53JZM+0w3v3WqbIhYi3
A5TOJQtZxtjKW0O+cAdsV/gDwydH3XtVfLuXIMla8xvltSH5ehSVV3cVfJizaNidcw6+p1w6PdCo
D0rL/FYUMLb0q0sYCs4ToUsUSeKDjQ8g4zTXz8ZknKXXTzjwooGHYXHqk6IymBAT/zO/7L1/cBw7
HXH37ki5kRMr3ByaXJipFGT6mUm5WwLntd8R6YtMd1yMKf0U1mQhUN6JMnui+qBL/7qzAjDQ1wHo
LJY+ZMuTvfLRoe2GOW9oQU1O5dhUsUGgBNaFXN7CxI3rvrZ8D3t517Tt72VoT2E2RFuU96rRn6V5
Vp4S06lLL1REosEd+ecJvh/iq4xZBNg8IG0W4cd4gqzHbxUHLUwoiZHc3z373ZSFJEfNknAdbfDz
88gGT4DZRZStP1nmNe76TyIp0eeodbrgNBm7NB0nsNRbrarNs+anyyygWIHeQVN0DRiQQqU6t+4M
LBmAKWOXHpxY9Q2hax7uGZE7qUmODOWzI3RAkdwl/9brxTQshQFDJmK3RWHRA3rFNPbcFwCYuatE
s07ysk7Q8We8TquH8+ry0xSaFSoAXyIrmTJ3/22npHZ3VeICVM/BwbYg2Mu+hDsHMTkWhxCDGf8w
YSn47dCK3hTGyaBmzyOXGlGMmwZ0RwnxDJcTT9pnoU0LHQd0ujsNRozTIp0+OKifX+zqtV1bkY1b
yUgf2jDhIwwyun14NQzlffo5qm20hTZbuk5u+8PjyY2NpuvVHK2Qf6Rmv7asDQ2Wpr4zW3EapcEE
MyWl7RAYY2+hpdWrBFedf5kak5RWv5odZCUpnMsfxB9yH/GoD3aAit00dw+42tvviqvo4loEO+jq
2rcvJuy66+OIOvCy1ciWaVOsgyKXj+VO0ZryJOpF3HwJHTJk6TXk4US8lZrHjmw+T5tLYeS2iU+B
rR+DlHkqWdWPMr+ySKeAkzvl4Ai9NjFH2a9oNlXx0iLBYFzk4YzlzAlmGtia7mX/nfMjN15nfoQi
e8N0/UDE7I3FN4dtXtyF4OiyRtV3I2D4YnUIL08jl6WMW+NeMxts12DD2oFBs5BxRsR+TMRXezYg
gmNTHMquBP3W6UepsQr6UW3RskNMLDoLB0QtYsrcOXTPHyp2KB3ciX0ob4+IeTyHCAja9BECCIy5
PddIKrNbr1jRfu/snClcpeDDkuWhRREbCySLHe0IBpyaZ4deSS/HYQdO3vqN7RebwvGtD7EzKOp8
4Wk2AWOf6JAitNhzULbPHatNrMSkDvQVQ8BPdBKN7nuOeniHOPm5xrrRObXB0N6J2Pbp8hpUpIXH
188ZHhnNjV/v18pN61Ovpi+zXndhkaUYgJ1HnHptiPg9hsiDVCK43PzD3TrkBhLN5YPb+VpeExog
ZLZkyinHk1XQA3mSMN9yHKzxzMpBe/ThEJV01BIzoS7ebCQCrugE/bSr/mINpgZiX05RhMy0k+Xm
XxDRmUSvuqsSnzsUY14wHfnNegAjDLXi6Em1yoKZMaY0gudKWVtfmWfKi93FWqDMv5Tr1xR+sDVb
bRYknsYbr8DP8T5JxfhexABjhDDn8WVxNWwT+RXIkCzFIVGOF+whorbK3kg65+ouOuLIMDsfRgTl
L4BrTp8zUpCksOEKNDGf4K9p5OHy2DMhU9tLxlsL5qABMzs3a5jUxVGBXGO4Q00QzOU5OJozWaAc
Yn0CIVyJzlspEGcpSbW7A0pkuzh7sKVLUT4sul55oFA2OaxhTQa7Qim2iSFWPmbgn4iQo/FWBuva
+NzFCocgAO2FzXd0p3CBkWgX3opz45XnLNW/MMwm/YJB6SgIng+WWSFgLrQIZTpH9zeM7RKZVUfj
ItHw2UTKH7/0q/9F3ap/pdPGshzLd8s2dbAIS0fnyaly4Fwel+3yiilD5F4WZNN+Rk9XThx+/IDi
jwbd/JW4kqXRgqz65xsEnizRkSueIblBwu+eY1xqjSr4QKc0lR+I2bsjtNbX4gdoy4GRP/fDUUvH
S9CT9DbBu04VBUrcGytcxkqoyJgs1vg271pjgM2LnNnxDcU7JnPsItBlCJSh5mLZBTCAQFUOfKUE
67GEtUg8McwXCyaI1UDaN4DX9to6t9WwF2cJYk+FfO3o2JKy1XgwTcFvijEjGwYhtLeFRCo+KcXF
Bl8rutt2ksKD4RRadEIU3iaTZOrhC00NfvT96BoiOblF0II+NCOfz2cR+5y2EX1TvIgtm5gBwjLJ
cxA5Z40AgzIrUOxa7RSg8SJ9nY/HaLmhCRSg24MGENUm1IgMHsQbOmkqvxwcfgyeTjHC+5/kfRea
1he89WNuTEs9zrVVpUEHlskUBjU/f/aMNnJ0D9Pw9y8pCiy6I+HdCDEPnq6Z7pUNNi7mIB/4H7O8
zuA2n3XEx071iLps1RdoYA2/UXdR4ZKwIKKgA1ch/truKckOOIwtjxUBapNqHdxnaB10FZlhd7cJ
gigz518Y3ucVoOe9Z+WsEBDLR25k4NvYl2J7G8lhRh1lS5zJQT+4CVvPFqmCwlv3sr6kbY6KDQj2
OQbnZgbxqxUWZhaEgy1laLEUAuWKf4avg1+cozbMW4zi0v4pjKy1H1gjU4ZpmGm6Sn8YOEWs4Eya
6PHwO0io4C8ONap55e7R5H9HC3zdeOeJil6oTFYqCBaTpJetn7/d6E24ciVzQWhGZxd6JN4TGTLt
gdsD8wNupoKovoH8SBAcsMlpqvM+qGhJzEjhaomvPjfcLSvXcDRhl23HmN1tAcNUNB9xLedn4OTE
YvDVxOBrjwU0z7eOGR7zUrRo84SVtpJ/yWzLEibBAK7yYafDjcm1idVbv7Hh6xwcvychCs74p99g
O8969pZj5mHa7etbjHTIDBosIpzWoXSf4XEEQH9Nxn1Fd6Y7LtQDgJyzUtwIy5fHOoGT8ux58tZx
22Loe6W5cpnlsmF5tH2vsL7lPFfLy9uxxyuvE6E7U7MM1uBVJUhKEJ3SDimBuNY6VzbWg8a5De/Q
SHiWnIeDKVKqaL61ZvzgLJ7gELwMKsE4Bz9CShB43vZdHGXoIWlBvdsFF0bpGskyrhaqvfr67w8x
s7Mqv1JWABb1Q0iX/jui39cqrtXosClZqBM4rE/J1hjkcyWUEgYu9mIf4uquBBugTiKc7lZD7q/f
SsQvroykft90I3gqUmJpAXRMhQn11F89ehZ/bifgoyVC1nECX8HciOwEqHQwQ007JOeQ36wrkO1e
xMOIV12pkDkLnlzfkE3mvXifdd26RpaCZpHp1w/RpVftPqS/egrUJ5JdaIwrIfovvJVciBu4cma4
J5b6edaR+wHp3tekGGD5pB6GENlTT7O/6Wspm/EI+co7RNbRnn04CVnXTXNgrcj9XFtdWyz4ejD2
Xd22FOMm+XkPI8cFT9H7aKcZeMImbgX34JHWSLrsRUXy+mxz1NXXA8QRcj5TZWZIkEl+0AysuL6Q
s21lbo0sgEMUaRashrkZTF5CToNuaPKj6rMqgflpyM/ARxEYUmfvmaEe/bO7BnERbqjn4XGGGe3g
XMY5EacTJOJT3qNs+loWhuwpfRpoHQYdJj74RZlbIw7vHFOkSpNIDu9mMXbfuLqPGcp8ioxUF1U8
SgkIqtpn6txsE+73CpipX98BDRu8JgJwOoeDio6HoIUySnLQvU46FQtDEqpiT093e3+nR7cOsChD
YhgCse9EdC0+ZT2gDIPRhNb3L7Pvpq9jB39RtX3qhsyCGTOKO4G0p02JamOXg33/LHijZRQw4auO
zka9EUJI79wfCsRJuIHzlBp+BtcIAgn24tK9Jst69Z9Z0joSxAjCLvaywK2BV+tBEHWvbPpsSsbo
t7SFkb2v1rw8TstHm6DlD9HYCucj3rnr81udwmQNVKWWsTUVbyRpwZNON1Us7Ql6uGSB78hwIvRm
QrP34mAVLsetj8IzQZdTz8ro08qZXfCUAe3f/B6igAp5VcmMMVAo9JXcJBXAmmAmi3RySGYlj6bs
cjclnU0qrCI6Pj/JuQLfcRTVmgLXaFyeCMtFJSA8G4jT8I5JzUyqQ+pfTko3nn0ReszmxUDSQvv1
+Dq31acuM5Xnb2Q9OhCqGd9JIcpTJK41n9Jx5Ua/xx5oqN6hUmmyhTcI9gEOgiHxsCL+NQWKLinP
hhat52mSXlGJ/AlJoO8+HeRkgx5ghmxddnGWTZRixZukozzC6dOZ8Q8GpQiFn8/kwbn+SM/EYoFJ
HlkSj2gGCuUlTBUJ5fWvIXR9t6+VLRKz55//eZgui/Gaa+2azhNqUYAOe0FVg9gJ+EYgmahKwscC
I92FD7+htq5apnG9k80DjJUJOIEQMy6BhKYkVdqPpJCL6bLZH07qSjIVYS4WxsorK9nD9cwYg7Kl
GFtw5JxwvgJJskkkzpjkA2F6+Bcb8cQ+4oMFsBZ3sq+xeRZVvsghEXWZPs9Rs+LQ+6LX9Lt/aVS+
exu+OISjsy4F/bkXMlJulvO0x5omhvKhJDErKiA76noGFsgmvCxAYzJ03VJ5IFwb+cyAOYGrDW1Y
qldyXN1YMdF5XiUrDYwO8lEACXMYVxJM8axcveAbXSyHMkdWNe3z/C9K0+Gh6yZ9ANMR/WV16tDB
ete7KX9i1IDUXp+OI8xsrfWSkHGRdX9lsCTZVVeceHtIKmqkVYZ6i9Sp5rNN0s7JLzK7KRB5UY2L
op/bxAfJKS97j735jHLCYyTo37HiSMDOaG383R51sgBPdJ9Fr+Lcjc2QclqxSqPZxaKkYLxrTmFO
J2FtacUwMyRtJBkWnB38f60Km6tOkxw/QCIslzUEQK726I3ypGjKCf3MH9T6v6R4r1qTZiocs1XG
fSAarJ8fkqfcC9qMFiEHQCTH19/Z25K692HkEXmoN9UopmmanUqSQR6h/MnOBSBwJ9qxIC3Ub31I
kyjSAxne34+ZrNVfV5Tg6DD6Z/HivFw3SxHLTh+BB1N+K+oBVw7QJzqi7PEHiOEaao1Abl4qm87i
9mAS5EqD6j4bofQGhBWfyCERrDnhVsp61Y+T8ZMXGvb1zbMevjpH6yxg+Vqs9ilPRZ3yTCTud9ib
UdhsHgN8YMEND4m0A2T7dgGzbcOs6rVn/BI+aQiOONM2kI1KfTFPvy6AgQbtA9Gjl4IK2Qxb5oXq
EIlgVAVZ/q77W3Ky/AQYOmJ+a+LSnf10dCcaHVbZ3lxz9867AEoCg9Wi03wzbKK/4OH/7Mo+Tx8J
gTQmX6MJoCABwSW8BiXLw2DxlxlsvRW43nf5ZxRfh9ReND0bgupDUHG5Dzbu1nJnLlHEIyqMprBy
XNcP8gNLtDCsEm4MoOVOTgu9xkPNr4Ay4ruD4bfuOSScj463n0OZF3HZWBhlcOinwUObTIMDXjy/
5GumcjEFIrpJ6VHFEy9VYUJvG+6TFhzuim5kKFsnXIdnPpv5sngtzXg5ZPCU/77xRoBdB6P2SujA
KmghyEOXGGeuNNrU2gkUDdil85hGE1quXQUHGrWZ7FYRMnUPb39pvt2IHvTlBGA9penlQdt15/Gx
XK8L5sWGwV+15fmb+8nRdbGY158wH+QZB0J31YiNPHJ8NHLhdtAEVBvUiUFjky1xVqKMATjkkjxE
vP/wpj0MffPVEvfma/jSyz+RUjDffYx3NpnI2LNft2zOnZGejnvExcUDmOwZ2HZICjfTkV2yQEej
NISKPTAhIPmVLddvWiLEdZh7cctb8jA2h8iQT+ygGA2UGDN4fAqlTzPHMScmKDId/qsbPbYy4gcw
7uy3UHdBjmXXsNkZoNmLkD7nBrNQFUd/dmrk5OY5uXcE8ArBnBL2/SDjBcAX+mBFV0cjmAtW6JTl
m5q6bBPcy7jvrQXYx3l7eU9L2ewPcnKvxkO/ccGPyxOetfniUhLf98bL6App1/zv2kWulFChYc8s
Ju9uDWNMdBc3cClUjYoDtdxaVUbs9ekPCqOMovOTeyuYdLL/vxpB4xYq+DEs/zsHM+Lz4TRc6p2c
m2u9qpx0bTkQ4AEOtt0l7nJKk4cs9cujXgom+XggJudw+7UTnAgfH9Zuq7N7EdGsirdyJAMB7blL
gYX+SO3gk76zNu6ARAhmbcQCYQGYQlEadHAOroIsLsJ4JiaGVQIvc3dr5D1vRKTI1sSV2hrpIL74
askCkF9Lep9h7TikC8s/HVSdGl9EbsLviTm8Q4Q9P8KRslVDZ0uvjyjSB63STOLXGuzoOLVV1RTq
xLy9cXo5v9YE8A8jqwqrqsm3NAqfCseHalaJ6ZirfxQrCxLV7zUdMKjV9TNPk8HL/Vhnoab+uTTw
kvNytXmcrUWT/JXXvMNjMMkTiqmfXoeqO6xM5ElHWNHbCNflhnNRvWlEUWz979IOokfIIFILKiKw
WQgDRYvNR7GaOcTgBz0ByIzYGOA0M3vfo7GEFoJHsm79mL5YxcF/sVD2WPiWn5lIHDqEmBWWxvBH
+0zxey2hlTrYh90YICmyIGtQayI4fKH3AfeFBhBBcHthoSf/V8svxfuJqVrNWsUM22V67dVbXye2
D0gRxbWyR/+yuJXpxlTPAY4DV6JL/vPkkfF+lZoBBFz35gGpzx3dLwKQutCdpe4HjGChE8t80Z0X
68qn6WZrzdg1i/jSyaa788ZHwIktxFJud5cztv4fq5frjyAzXQNpUixTONt+Z0ppeWF/B96N3v+/
nWd9aYczWG8sRYzK2+sxvbsnYn0rLUDnOwzd6p9UtFI3aJOv5XpEv/q3+0BbLybsbY0b6Jj5DiW2
pjYiork5Ib0P5c8SMoQuXRrd0rrgvxYcNACjAeajVE+x5MJNdibiHOVMY1NQ9lUkTUXUjvLBiWjm
uSmeYMvgNfz0NanCDFDifLxbKyv/Fco0WExDyV+EkpgS2e70iLKATljTCdWQmslI2j3JsRy08Ocx
MYVURoKXfdcta2FIfZ3MOYLot/bwBoH05Wht9DzTHv4aVeOM+aWYXc2Y5ZfiURa//zxDCgezzHkF
GkUHsciBbY9IEtbt2uSxW/2Rsq2KzDhfqxSlZJa6UGIG4j/vP6pB5k/i9ujA2Chu3ISSlIiL6VnD
2zBxmS+BtxQwECzCCVtUa1e/BLbKvLcawzLs/kBBcKNdDcudSZzlnHcUAzdHCpvT/dhr+cV3Iq9x
y9yKwXI2XoMR5sD9Km8WYSKA3MO9KY4bkiC+PDGhpkv/UdoqGvOtS0QTUFNQHbEcrf5E0qVunOJz
t/fiza20hWfBGcWiImckufH8zpkWEQsobMS0yRLvgd5rWLRhYjNvB/w49xTzCRBIdBjOG6TbXb13
Kcv58kNtLE2vvyE0dLXcPkm17U1kHq1RleVV1OYsNHlPGd/Ui1H7LGLQ9n980q3rI2fe4LrjB/Oa
Et3Xu80MGNYYX9tQdb5paqDK4ZxSsdM0gkn/9OD/TOueSA3LYrE2zIyvYH1tYaAX1iHgqH1DD4we
WL5dTaDLY09eVJck8SXpBBgRD2RKZ6HxDrA3l/Xekma1lEttCbQxWIju9+qcSYHQTBU1G0Shg01G
wEiSCDP9xqVN9cYmZz7bRahn/5BtlnfZ4gtSNDJAx0jG468fc8kgUAKU6xnUxDJdh18jnjLlM8sJ
uwADhVseAsMnMaGPv6bvFz4EAhm0OAWQ2B5LIgRewiNw5qjDXhW8hSkMeHkV7dv+d0wXxIW3uYe8
7UrjjV7JDWZAEnh2gVDaI8sI4YEI5MuDdg4YhBJs70Ln6XmmUwjK94ijD9M6OJOC3UQDSXW52Cdb
X+YDze1Y5mCZjvqELQrBXovsDHO3VjPtyLxAYQ6Vhi/ViPNW1TW9vLcu3g0yeKY+MMKVEJGSwR4R
Qz8zIleJvXlW1hXvOGrT1JAZoS2I+UPtHN8A1uCyvuWrj0I+4QsyX41WttjZ0hKby4Bpnkh1rMCN
V+zIgfRhfuJyc3jYHnbAb8ZXGkB7H11vMMH7ZO+yVS5ceWP3pEgFOHdiewe2A7NrPznoE2+Aojj8
oZYGhqoPRmyuGTg4o1PfJKdk5Qc/LdjUDcx/utn5ohGbhwtxLS7NkY8eh9BDaPCJPisa/EbqCTSX
ZaB83z07yL1KOs1GEI5RgTmvqBObCZsCYfx5SrWVMC2dPmgEhLakzN5TDfifU5ViWorwU+NVvUz6
4Ay7WVeVNO5CgNiZmBL5LvCZy144NMeZIOHsIqEM7uy1Bktji9KLfodqmnC/cMJKkjbwTWU6Gs1b
j3WyuRzRrHa9uYsWRMDtAhtFGVz19TysJjTvF+fUXUkCe5nKvpSvwrxDZv/DV97X2OPgk5Vayeai
ZuQlMjjYLtOBfjjL9M451EOLALRKfC3L/t2rfqWN97MGJxq5O/n3YWpXKY5VplOSgerDaXileQKe
hYotbMB4xveobQdSCLwdiKTFjdQyI1/e3FfmaZL7L0diXieTN7Q8S1JhPU6K3zFSpkm9pbvTpjN3
HIzBP9fTQxKv7TCecpvlFMQHdNvXHiYF/EJO+fmbogNWUAVSQZSQ6sZdjCPPXZ8uC0EY22W4eCyN
k/wz9rB+cCsvMVAHQjf/weEZDWKrfZdlYxbRsQkutD7ZYMcaO1mDV4neDzF+yyg0K52b2H9JMlVI
xcF2jLUbjwqH2hf+K0VgtcDmuUxAH6LJEzDxMk7ZjhCzkmiNIXelAzrdRAt/ierhgJsU9tiKi/ig
AkxV3DSAi2v4gu5bDEb28ZIsJJj46/+X6+SeLJoElLO5rqH5TEbsYMOzm6LwW8zWnDsljCskmC1R
5XOzmRgt5MFWIL5XkzBa/l/Llo8iiOnNrqLUWGPZRMvSAHo0ThW569+G22EharWiyYwTNn9xBnhh
10mzQgsUW/miFZ0aibL/GN+1tug8i/4OUR0cT0hYWFtul96K6ILyDWcoeiY6t9o/5S7+mY70dxge
fC4XYP0ByTBEWAgnvaJmXA7sXj4rkbf+cGCUt8NwIvgvUjilkJcGVapJU+7wRfmdekVOH81dJlW/
CHbEgzpAvJBRw+MJIyPlMYt+aieEPrGuGBvnI8r7EzFh52kMzwJ7tRLhXXzUzJqG8w/dRW4xPMSV
lysAkFPdyT1dYF6BE66LaQCyOMQ+/9CBs39E8quuN9T6/+jTPl2EvbGz0IOAo91z7nBZTPAeV3S7
w7HFxMt+MCL5mZhyR0AMtjki8jSmxn77IRkOYiL5oz1XETZDfyqp6lJtWBxKM8KyaxC0TSrS2y2Z
PChZq4TJrcUgMPCiNTgowZmHFiMVazjy6EmMtcQV8R2e1+MWui3vYvLUsqzpFqcXrrWO1tTsFwW5
tI1ppZJdWkW/YIAIoqhy+pkDiTDzPeMRYz5Q03dfMH5iyITzGJwaONBJT/B7djQ8vQZu1qAIEwK3
aaCgyedBq6DqY4pVlJmQMarEul2SNwpE/pLrJI24PoiCGF/s+iFu1xTGp/LIV2yaySFTKn8JdiKJ
/4vjBHvAShGT0ACp0o9QdEYxF3tOQkQh8ehoSevDpj0nJ1GmgqTONpwhrFMc/TGQPQQBTkjVZU24
kOHiE/+XQ3xrDvh0tlTZjFPubVlOgUyIIXfz1toH2ab3BmM14k6/uRQISGCP9O/B08royWaJtV3D
XgA44jbgppom/l+JVfdqSVij3gG9gfz+AON+WPFT5i+GQ6sbnfR2Y1AVs1PDkN/MrVD1p7Zng274
J5w7zSnnExT9CJkZ5MBLytW/ic01Zmf3h8A9m97rRRVSCFOTHewcOePdMKIY4GWc/Xlc2GBKx7Ii
SyuKjiPhfFqhwlV47N/q0MMiBiWJ/aH1U2oXejbpS0O1SlLOXcMeCnTddpkZhiiRDjvxEICXZhTN
IwwJO4t/y2twN6sl/suNlEiZQMZmaini9w4xZY0j0KpIXo8SXskPS1LjZVWN6pz3QhqlXOB/cSxF
DjUorzls7I+cQ82lMGCq81KhVHsC1ccBtdfGg1UFWuTIW1uQiJOOQGOp8MzLVCzP0Fqxid0YdxLB
E77iSKz6U4Xr6xWtY8Ly/wWI0nLChcpRcggDpx5SyAiFrXlCUqXJSJ096kHjm2HwDFA6jWUx+K+w
LXk9XeQa9zXeMOqs8TWbrbdaRbz/7kicHjA6uuKBk9Pw1krGiXaleETqkI+U59GUkjFFuQHieV1H
YSjJu0sh/ru2wpJh9tzvNKz1nj6sOzf+LouGuVufE6ZUzRtz/KXz78RxWiLXNR6dmMDlFgxBFzYY
RURS7PsF+OFRY5/jT9fJi/0rIqyQN7E6tQhnfbTU+T5i4nGxYOoswL1LaojiBD6TIV6JM4QULTuD
7yaeH2tj9EioA+dl4ah/AvvDfnonTbyIk07PLgtDOAUCtoug5U1kjDJ+NG+wiFzxJKD+2wxF2K+2
8u8GCssBHd01K75hTkVu7Z+3jAqzQN33kz080xmqcsPxkNVk+f4B5Xh0WRTIXIFaRJsC2dQ+zEqn
RQ0Ih7clB9iSohqic7F3X4THGN/FdoXSvnMmuGnmoVT3TgvC55Dp5EiYwQLtqM+E8kGKVQnNJ+GD
nEyYsOnhRIHYRe0Qa6NTR/BRhp5camadH6FiGfoP1yyTO40igJpW+5h1PqIqYb8Dt/tQ0+3ftnoU
q5KP8/Vu5FlUy6jWZ+dB87ju4eKdAFLt5v4bJ8LYGg53LRCFu5ZIsoFwD0kahVtP+LeR1OeXwywQ
TGeA/ItLfu7IUZrx707KAagKrm3JsP/9GSoa7m0xaL3GkbLQva+dxfJSS2bOxIjZjeuPoqGkSJzT
WgR97yyDDE+Vk3CSSUM6jVK06zMKA8LSvVwG90/Uz+hm2LC9RCIsOOB+ZvwpQ4OMm4ZDhIIzmQGq
OIjeV0C7ubG+WSNgZ76vwn2aWI/KenJqUtHjOU/dTnx9ve5CJZkqco92NMqvuvTykEQj5NzL/LXH
YminWndnLXuod2b0j04UODnH9yKJj9EUqW/tGMmCZph/LsOFo9F3jn83ovjxEga7sUgNLNzGazEg
bc79fmQCX+N/BPfe0+1k+LAWx6fAsligl0ctfhZTvfjWNoXBPoMm0KocZyZa3tXkdj1QT6sEBAV4
Rb0gFULn4VpzpRyEvGIJYVXX5dyQASxKTYxn8X+WbQ8vr0EQBgIGXXpwlJPdHpis6MHRsXureCQv
nYmgkNwYOhwembZNlmoAecsb1mOWJqraA7qRQol0ThV4o7YJz/c05VHTL3GbfQbabm+whzZMzNkS
N0x2+yLzu/8RwCiDL4Fh+9w4mBKPolx9RWgC/C1+H4AKJawxqLDapESAp3vtiQF4RkR92W64Im+a
OfScocJAuciqHXxo0+TTc0oCf+FN1mw88agofWLSxz6xjhWxQ9yiuzU2cHzhNMkJxIUuLfnO3N2R
X8pQIbV0pBoRRbQN78hO8kEzcOK62IWevMUxzD8P3rfECEr2xxTptPq0UO4B33fj+Lv5pQ2CvlDn
jMlWMqiF9f6GV7rK75by0FtskilDEhMcGPmp8H6goT6K/s+r0iqH3lNGck9bnRP9d6FF6sRskqCh
5hZUxKMy2GAv54zxFCgM600z4VLk4mwD89wrJsqDImycAlbonx0e4zVzn1ZfVHy1iIEB7bLe/5h/
cKW4NzqK5qX4KR90b+eijOnwcn0HLshhBXQbMMPbHZC4rGWdg3P5v6S+B48LCLACUhNjYWrXF/8O
PdKiupsvOPpa2ZFE8rwf+04JptfgkGf3wpVIHdfVLDyOtJCRHwAoQ2nNHRV1oWOX/RThvPiSE8wQ
cxmB325PXtaOeMN6P9CMx59fcrw/5KqLWq30M0+pV8vdFaNIAfWuX5dlpERr6Y2S5f5z1ROw8GBm
BtuU/HyhVdewPiNmoppiSXL/bCsUEqYuMkHzcANhgMY2HBFz7yrgpBGhfa9T9+QNO+tlTMb8IPPr
TFAXchh2ETGALsxiWfppOXOb85ev12HX6Dr+1iShYywqfZtaJ9rL8EhHFDh4CNTs0uHKqo2MgnlW
2N04lRzq4ESld+Huv5aQvXexyfAXw0TekLrbZ/rAi8+Ft05fVhTiZLOYbu497Rr3BGzqPp+L27ef
OCP2bPqpwUnbUgCIjXFUsQbGJ0ui5il78E3H6jwWk2LwObTv8YePqJjR5HHfncFK0l9VuXsN72oa
jaylmIgEHnWLtMyk/HjJivxeE78HH9pF2l7QTTsZ6OdDH6nJn/BF8WDydpf/ygvtnLK+3svGOVB6
h7ghA+70GI+6kSC6GMZ1U+2ND07yTcWRO/eGFJlXThiJxKvavXjvM2D1cPVK1faZ1urDA41flAKZ
pSxJBjtBJfjlZTLuYiDyrRDQIc5hqWAtYQGZpzZZtDMQnnW74UYhy2tVq/T0UnPGU/okXb7oaTmi
AWOvFbBi8l7G+NlhgkjO4HpHmDXEPy//wLbWRYCkWJbCCSOFH+bQGycITGOZ8sr68IoI58GiLvO7
04ZyJNxc4GswhW8fvMvhqvXPKoZvLik34sygiT5MbcmbLHkj2Rs1gfVTg35DAR8sivG9IJ91e2Fj
bUERheEhIyDbHdtb2ABp5GMGgPxvQ1hqBIUV3drmdBpypBk09zq6lMLgb8QcZL5cLNrtc5J8kHVu
6Zn94RgRh/h7+i1KgEvk0okHRQusutyrqG9/14w1oGYyaH8pNJIwWrhDxdjBzGyYRihwASVWtUmz
cysDsLhvFPub8DdvK0bqrcKssx8Lw2X7Y8UoZhcEEHsBUS+QeNZYzzpP/C+sZ/3DAEhxAf4r+S8x
ZVskee1IV5AHkzD7H5N8lLN8JNmoGPCUceLuwZXGGKflBInHNknddEbtQRVCCgN0TADvdUS0zugr
uO/II8FyGO67J/03GIUt2jQyRdl70GqUJV4BdO6ALOs6anWKXOBhJg4ebM48z5+comunahIOL+mn
cQ+6Fk2iVQaCzfFEjc+xiID7uNPvUccgttZqFpiVgQ+3VSX/VOIfatkTIlnI59KAQLlfQGoC6aiC
NBEa7VTbxipTDHVyr9SO8sWzNKvGVW0RN73tgoUBtPi2t/r/tPIXUMJ44HKqgoltddWXs1kNtrly
xq2jAvKRB/RIuf+5cKfti8uxopHYQRrUqbXlvJX+28uL8WQ/5ybK2MgZR4PRS3VZ+v8ehN9LSgRR
UYj8YK/fibaI5GAufkZ6uFpI5gVOVP4x+tCiPkfQ2f9Hjvv1d+S0GCEJNUkjy/lfoIkARktB+X/J
NYWHkdjktiDVRxgjgFNY7OdFA1eYPkdTXG1Lwh+JSUg99DxsnnZLkRguKecpWfrGBGvsPbYskpsr
0S+w2dFP0IGM7CBGjIZFNpl6ai2Xq7l3uLocx5nbrZSUF29mhquXVGVdpmBOQ3UK3zNkeiImYfvL
UZS7/AkCiOfwDlZ1dPbftvBSKbB2eEeb9NCNRWHxmpRPg5VMuy8rTKZEoP7qihq3rOZZFHuVPP5O
IhJPQ7c1vTIAJNpmZ7+b1cPa7O6LPWf/ttuQueGp+EACBFtkkohAOLS40aL8R/eInYRSvyWU808h
X8sdU3C2Hzjk/XneovUf2VrFoU5kAW1SDTXwUc5XKmHDvSOd5sdmRlhP3Yqdn8YRCzySzp5vLqKR
mD0nw8d4g3LD8ttIDlSuYVseqBy4uffNE+Z+zRSY5ZFOXfxfzHjoZgsuN5+p5KcQJqZAYOV/77Hn
PZuJ24SPXK6oqQ0PBnVvGw3LbiB8dFMwlJ/hncf8rHyMb4i/cwOPCefnh3XZ1KutspSKF7RIzFOR
g5QiHcO0RFmpkkyYhNymJlfTUdz+GFuqHeuhr+0fm2dC23rJbxnpwwSa7DLgrre9v2WxgK3NZUBD
S/px9UU3oQI9s2XxJrKZVR8ahffVskghvjxKbVHOng8UOA6PciCTG6fBwmrvpoOqUMOtCJ4Yngn8
ERCQ6Xy0NX9TtmzOW1DMzqhb7JwM0PFp8vLmP7+JJUOv7c4DbTTILCAZI5P34BZo3gKm9izKy0px
sA9CsDd+rJAZFic/Fr50M4VViCUSMYDYvHlOCxyIJofZSoVEBN+LLCr+aZsZZsIEjv8vOEDdI24a
ttZTnmMQldlKrWLlC8EUeHNceaUbM/9Ucef61h9j97OaQylPnwPf4B7BCAscutq0VVqrdVIx42lx
FP6LynO0O5lOsyowpnxFHZnYObk1FbT9SRA0AeyTMuufsOmUGWN1XARqMUW11wzMMhtTbR8ppzGi
33XNYmwxC83eYVp6WEqZAIwoU8fDVsUM1pQjQkRAsV4etzo/Jmv3VMRjxwlL/kdTiW1ZGjMDgQ31
rnCiUdUz3wM1JM97xYosM1+vfV64lQDOxkkmvovLI3Hwz2c2WG25b+g5InbKax5XV+RDCGfayk4S
mQp2EvemLlmN8aNSXxl8wnxkh5qjySAnCuPK+NuUN2toYLQkhBetTKZ+9iOQKASPG/5z6PF7LsVz
TvwLKhHCQxqNufcZUQ7GqBEuw/lNUsEncClFfCW7L/TV4smld9MTg9I8O23r2AgXimpx58blpFN2
HaTUw26H4L77TQpixjJw//3ChkdkKRZLHJBdd9ppDoK7vi+uDKtIyeT8l9mbTZ86GyyzHsgq4nsZ
cxNSLtw7EqzwBnKGYRYzm6oNwZ/j4wzw+60F5aQB5k92S4OIjHxB7S4/gRJltOGXQ7jbHWU0j1L+
Mm+SyCjCu+a0InOMnIEuXoTMrQgfgxY4wXn7lCIph94L4UVhmczM63VCSVj/pJosr7H9WM6jNV5s
lLuYg+I04CaSIQNgEAC99m+68pIR/1DZcxiAyDnuVHRmsnwel0JolFNTc1M+iVtEk1XxM6KNYVYA
8xy4XOk1iDr1ptIZ7oLNPVrYOSOkxGhOMmuwWodGxW5xCeJ8gTuxzYaONXtOe/ZSQo+3f86fiqCY
i+RspVQuUhabmScWim5gWnbokLHAckp4LAPFzyWzIcsz/XjU/U0KonTR9gnxj6A1+Jf+P4Pm6e+U
rLx9Fv5Ox2zgd5dA8zvEPO1COWsxS1sev4d7sEbV/+0PqU+4MlbGvKHMqfBvBlNDfoQbxdD3YQFZ
URa8uDhbBt6c0DSQikFugXJk+MUMoOv0dy+TN09NJT+JL4t88P2EJHCO2hdqUt1BiHtyd9CK0yR9
JibfPng60Yrl/rWkO/XGRXr8w3XJKhvwyOWG8bJvW8OsicXSp+dN5GZ0uTOIwn13Fj8AUvdYgB5I
5rvbg1/WvgoKBKJ2eJ6UWyZH0O7arJ+v7LLTzhzBWj8LiyvoJEsXWSag3e/oGACd1yQUdwueDl6V
BKwidN3Nf+oO3r8k3Imwj6alTbqJLfEmc51yFc4vkuu1/DoB5KqrexZGg4TPZzCTsiNzn+vUcVgJ
Hax+RncQP/tjIy0M0w+Rvl8xho+gAC8SsB6QSx3T9MESN392jRmXk9qJuOB6utprMqsuT9c92OZS
BJvDH8o8fsjlKFUoHwS0IP0l2BjUBgFQoIaUDPXkBoAal+0SE/Z/5+Q0wInoQg3hCVzU0K7V2dJ2
2kOK/o3zt4eXLhKrQ7t1aFLELyzLiCKKl6JkQcYrcmXnxxXh4GpUiDsnoKXzsqmuEzxlQkaoJkCe
pcpYipMaCj0Zw3sQyPhYeuC/wyOtCdqAa+OAEfxgtxj7/o10EL176pre2NrZZ3arIvx7xjjATAyE
L67FMSwNTsiZ94ZYwXaTFZ1vqVuVJd/J3tilRFlcfNA2D2ib1GaCwalwMT/p4uCOjp45mor1mFlk
QJIK9rxO5LzJmdCrsK44k20BKryqPd0JEbXUBlFYS6izUrVVBCqTX/d/GX+8ubJ705PLciH8cDUU
/8CLpahIHTp+Irf4QBrtLDHb3pqYCTumgwZtlU2BW/0lSWYjzx8QvyYXyXMcMmGImJ2PgS3eAapM
jnZglsFougZgeKmUrLOukM90anBs28nKFXMhS7MjfN4isEwvVZbgRa/pTwPKB2LUauIu5KfH3JNS
Fs/6SI07wAYoBbJ43D4HG/Xz3/DMQFP9A3biQ4qxwcOnQBBaeQQl1c/7o1sb/LM5q2JBY3WXj6bo
yFs/PX73SChMxlwFQl6ftUN/tbKAUJsTbWFQDqX0JeYQbS+qSWV3ppyKh/282aVYwP39SE0DY9yK
y50Oh739rMQ0kTH3yNXiximdqr6rLH+CnpiiUiIkQhoOcF0j4a93+vCqn9SR0i2Fikho9wUtswMz
ekcjvuf0YWVVWXTQ4TRlL9ZWHf+Ah7mAymr17OVZouc/iHsAriMUtMQb5/OlOpw1V3wg5rX42pJ8
I5At+h6F7F3VGxa6bryz1BRnPLCkvEYaqwK67WVw0+42T8QlDEQFClqJ69L+jhesCSimQH+wI4AC
454SV+QJrzNyZgo7T3lz0Ha/Drj7n6yBpKy8INUUrs03DIjThnr2FW8zfK0RjK/7oq3Sy6K/J7H0
BFkEAkkdQTkEnCb28jmRcw0HpHEz8zJtQQlXVmv+D28Pzgt6BQRI0UyQfXcNEFEWa/N0MeppKW2L
7WbMGIjeJEMFC8+jWuSAzmaUX2XxF6/tU23eWsEKFfX8lDXKjscMIEbC6cLUY0Pium4/3vITKAxJ
MctB8wveQQUBT8bkv4rvHvIQ48JEWum0PuitvtfwJi8pU1rXoFfoEs5BdhzUMiQVv3+73he353QE
ebtzr5wxd3GFW78fJV+lQGCCNvS+lL+pIvO8D0dDcX5JY0SUVWwSVNsZkLTjNjfMIlnVfkmvvRAU
Ab6GjaBpsGn9khumHj72+oefAHZ1tmDshD8L4FS8recwsTYHNO9aIH0dATYV//s9gB6FHfwckGuj
d4Pt84Eb546VZ2M9dpbKWqgqoPzdhzIW5FynfL3aY/iHTPsyI+Hw/xx/RUJHp8D3cburfs0AGHZ/
peC4HvIZSXK/TnEVTKhcjVQfKxGvBHIlvIoojQJCMBCarbFHV3BtCx3AhXLOykTBrQeyQu4tqO/A
AFFbj0wMhvJUt2NdRFQ1PRNh4AdysKgAf97rg6PUGN/14NUSf2DWccJ8tvc5Z6AMzdhur35aTyvW
dHcCzXH93JFcimrrXcitEI6MLfzABPReHCJp9On+cNdaIWrAf86eINUQdjDUx4VCo3tZ/cnfwP++
xIkee0OAhQ+0edAuAcRJUyoNIWLhx+MYXpzke1ogcvTrU8CFmoiV3jZvvvAtWpI8vqapaTOncsv4
IMzmvaPHNQZ7MuTsBaYi8IVag2tHF0xlk6lnEM8UMJMM+IgHk+tgvWv7ls2ECQMMwQJtiqk3+hLZ
W/hn9UiyDhsKYLV0dHLUptZFAhd1IdCnBLfEgYfXxjkpaKHkyGjrHqped4xZZAsCKQDGCyvPhyFF
Eu06pEg8/YW+IA/qY+4TPAb7h2cZkClKCo9NBAQIGsI6FG+nRx8VMocaezzf1Je5/L9HOnOwE1JC
FUpoqFEKzLCKvET/hiZMlhet0liuBTR3NBnqwDooIT1qnPjgbszHcFfclFFdnvqRbv3kmdu5rT6G
gky/WtivLAaC9JPF3r51gQnJrMQs409R9X2LTGrxHn7NHA2smP02997SxpfNiMH5IwHaWMzvEHoB
8EbyyTlbt0BOkhr8bUDbxxKZYkq3g9ZHC0e6vlmx0KoiEeEjT1JpIwpQkv8DRYI1gtWKfPyXeTIb
yVTB4VWfqpEeJ/vf7pkFos569OZUSIs4rdzAerS2vSeUtxxXVxRSe5eFm1vY1kHA5cAldPRr31Zc
NVKivfYuygTQLdRpT1DuPJ8/pSVEB1NpeSU75w+Xdzi6UvD7y4X+OWu4l3/RLMg4N5LdFo18kBmg
8Y8GSadusMg9B5ljSBnqI2oiu9uk1p5i3B6fOkQ040qWJGwXh54COtmgks675QIckz+hyWC8Kv5O
LQbPDjDBhJR61yWS3Cm81N4RAj1EtOhL8Hkr0cYN4rQ0R06OBrzmsMllwjmhRF2gFQTYnj7vdna8
tAxMcnKRRfez06B0KAARDZVSsbuJw9uJNn1TUBVBK3xZCCsbucMQZoK3oHwzhttBgPD07DHTbBeI
V6YEkSMT8Vf3ys8HyIu28wJspPld+9YvKrMg6jaEHwoXprWMzR6d+s1fST1Esl1A+Ifrj/FX2EKo
V5wh36ABoZC8uesDsGdUisFqTExAMYZeAz9FnAJghyPx8GahCtc31gCfOUVZ3i6y3xMExvgPUrmY
ViM+aNIV14SjMo2GpzNRPON9NM+5gWFWd5jHybSeNUAt/dkMJR46cMpZhd3qqXSlvcdxMTWpc6Re
hfIBsVedRd9YnVlHQOX/YRhiYO9fUA+87kRKNul4KGukfJbkVWOLFXmuXtd5w7eQHXISKyScrIz0
88P6CU5rjqGfbPqAjV6rJ7hnMtH/OFP3t6swrJxZNkhoA8QmB+loPI1i0qJaMmTH8z2gGRCu36rx
D6wVgWUm5XaUgDAYpBk/zMTaOh76pRAHyYmWQW3PimoYtN0asCMsc7Dusakk7d3YKxpFpElecnZ6
+L8kGIR5W1wiin3qrjf+NRgy2pdOCbra9EJTSHSEYLpS5b3W/b1OFAZwb1QYxS+ZZPIl6G0p3bx+
P0QtxDam8zfRd9Sqv78MZ3p+zpdStY8rIylO3ko1EI3PV8Pqun7fJfbYTNymQmSCLufnDLeAWYvL
i1bdRk9fpcgIj+KwNxd5HbzXfF+KNrXNjT//QKFxZTAzze2tTjqeJtCCbte9JGyXPv24jM0uBE9j
TlhHNMBCvWQayzVA9Y7W8gyNnEQ1/5DteGVp7LgWn2vc1bfkBgACVau53ETb4uG9wpSvgYAMB7Xy
UadrSnuBise8cxwf/aNPr7t0ugJtnGEsMFRSXy9J3G83JQeDjxm8IASc62XhBmEsK0cM6dnmKCH5
9Wmmgb0Z4NK2bVykQ1aRrV39oQ+h7hCrT2UVmgryNkiCGZbqD9mZkXW+OXaz20QJ3zeypIDfP1d/
UWxsrkOJNLra4434FRFoBk66VmT296xMXXkEVD/AVK8FzV8J1DHzidwQtvxxWFLIqH+NbqEYiove
94BuBQkIxa8WEuCWOcI2u6otg0oArYm5MFgq5J4rKNTnFKymxb1gieEgc/azndbRJiZaKUMOia3W
C3MlR90bMMcOmuK6sZvTZPH+b+1tOIndIyoxtxUOUWaX2db9BoL+7dj4oCtZchOqZftktn97hh+4
Q0Z7R3UhZSper93IctSHt6g5azFGzbl5fRlC490FIzM1Y0mDgH3k66HogswIHloMmyQT3KJSzbrE
uS6CH4vFhH/7EzKKHILYWFow6r80sJjVt95TKzgq4+9BYdy3Kq6/thA8X6ngLmdlOsKQGOhiJMqm
DRE8+x09IsDfJcn61h+zo04FN8O9sjjSUuEbleTKVA579mDzECc9Aax0nxiAaVWALjxsWfuLSGaD
JLD1MODDtO0Dz5H8QNQ5vzGOwfqOPW4NPDwRv85MqPdSPDJNBoo29rJUMqm/92AnTaqJ5GhUMpp4
idK/TcG2FlMJIx2Kh+u1dFotr9Mi11u17zj2GxnPmCLgDIv7EZdHUcHL9NRoMP0VXzrBU6DbKSjQ
2sKxqQxSoyEwmZS3/MRguefH9QDIgh4d3BdDh+JymvT9bCZwDt4e/e8c57L36WOElrCK389VPB0+
sTsCmtd9vawYcGLkSwKFJj0l78kGXNsQgrm7m/SfWFR/UxYrj98BgQskkZO4LNis57BLdq1SYONE
+6bwGrGxAUQqK6CItfgPK2oTGmOAKzDxazgiSBLCW8sh3ABvRB/o9upn1/4BAJx3yy9DYP2wva8E
6vf59zWY61Y/IMvlJ5m6Qf/zLK+YkTp+4ND2pKomYuaCkX4DQqMWvQehi0ECYYc1H0t1mRgnzcyP
jQZQiR4juWifM55lpeVZcG/zDoNr97irD2rppbDQWT7fqkcrRaadiUGr6y/f8aUchNTnMQ3sf6hC
N+eR/MVAXieaTT5meortVxj9b8MGuWwFlNm/uNjh2/8XZo+LqqzyWcqNDCR2IN1NHv4iWWLa0epM
eq7hi7duGmSXUoK4URZaeKm9oMELBE4VhnSFlZyo9VDgn2+a849ZKByapNGl7VdOYpLiW80BNC0E
8eyXd3b1WpNZGLvIMDn9MCprFolbpzbOFbuqpwIm6b1XI0/IhHJZ03sEtTaBn2ZyIrS3HhL41a4z
vjOvzBlCWVSll44FRAFQLGxOs4hyDthv9RfcifFOPI7hBAAGDK088A7/pCk1KLBcZH+89zEwyTt+
hQTJVUdyPJBPqfhgckCHGA58hlfryWPkOiT0XylSw3mXwGTZpNq8+QWROinnA/FBHa5/a7/u8nxf
bZegtTd9h3dghgZby/qiHQN59F0c0+CTj2hBIKEaiIwTq3S3E1p2GTjoGbqrE1DXRnZETqaM5Rrv
GDRmjojJ2TNPYIkOZhzrXjAS0Qyv3jBXhKD9Mt5BUngTHeH9PgCvNUZ1FaLGiGKJ3VkTAlvYPSff
J2iueh0EvVDtmDf1BgkIzm/Tijonrf4lvXD4Q1ZkX/Kh0j8uYjOaAagZjjesehGkOKSIfU9Ike5n
u8Zbc8xnFOmEDExQxU5akfeJf4UxoB+9DR+3f8FVZIc/XhJBn5HA0h93C4KO6Ay/gnkvRUORIAyX
jGL2h5pbW7TTkuyshcGP0l56AGWYgr5oNvzRtf5IqtAVlWpaC1EGxnDNUP5Kh+EURbHKAKjrWBBQ
zj1fuX++5INEArNAlRTEAqh1dbDyVzeEZ9Xri7s/ClCVOp/wCzf00okHy+LaAjzSwm5NyKtsiiGs
hXVQJF9JFiD74CgcvLc4f5Punmfh66nGuEOaYHA5koKQAGfpkB+Etn4dAsa5oynM/y+XJdMbji2t
PSGQPUoPYlJKbZdoY9nU6Off5i/Mm3gCszIBkg6EnN+QkKT/L6b0zcjBG9pURZZ8/mJvocRg10pg
CeEaGysaCKG5kt7rba1Rj2CFK2lkKVpRtz8ylaOvTBkhTnerVcADOuzxQxUxldL7M15Cl5rglYnG
wPi+7eCx65bCslQb9ydvDOfvY77m8JFAMMzZSDBrDaW9dHTt2Oo41ZrdpUH874LyFf3LZHOGRyn9
vDovmAFq6ZrIR96fGhCe3oRfiakgTaKuxz+3KzVujYJ778J2svrYZzBQnrhgs5sVaAwekl9U42jn
N8OGC0JxVCcaTv31/n8ZV2OoqDQsgycbMqmpbnzKbEDyPAcisBgyutpr7nDLcRlZ8jIY6pUeJp4D
/Tpom8PUOMfN8twP27fv59W/m25CmRahDBIqqK+My+pddODeWwQdgNKwLohYdQoQi+9ZqHxqhd5J
kIWCxchZBcet+DGNJ2A1sb8HqvbmJFrFWsQb6FiGtrw7gmZik7KV/ER1Ktt3lzDQNwqanI55l/KH
XUN50R3s8+TwiZyz92yPoSRGQaBhrUNfDHeoVShf4GaAv5XjQny/EIyWSiffJOUjmRSpZ3tGLX9A
N4qD6lsZl84rVo8UA615cMRXg0I+dxyMQA3Tt8y1P09Pa/z/IiVlwMTAO/0OViM7hwpRLlcQ3Ltm
Pos5DbKW5qJnH5rAAOQz6sZDi0sjGhnZz6OhyIPwYSI7UI2JfDjThz9w3FWU3X3meKzBAhgt402r
p0REXWu40zFGduDM0aH8rqyBflcCSi+n4iFkczH4mKItJc+UiKtys8mQ+ehR5bRY1MpD7eEbPkSZ
fVyhKoXUyYcVkpWutDNhEMsYfqie0lS3H+OXPFWM2hydX3Qh9Im0u2xIynUmq2s4sPHHZLtua24k
VG11nTe6DC0TahZ96oYwLUBRqmX+NTNeEWEcRyFdcsG1kPx8j1b2C9CaIwl1BsL05tWD/3JADfSQ
pns85TPPF3eHJUOozRa1s4pqWbgMx8paBsCiHhgr0zaxoQKAARCUbTexj7oRc/YQaaqTEaeyO2V0
Nd4SSijgJff4gvLuvvCCUUeyGvKr8S6PuKV+UCgNUaHcmPqWgYLoYn2Gx+fxuBUTj+j1l0e7Q5CQ
XHD/cP52YyNIi9HGaIZkkBw62a/BLX4HMPsjNFyv2ipj/L1Z3Iq9XM9AWsL0rLpbpgYiO3XDnuhu
+IrEQ4TEMbvKymc33LU0BFsWUlf8qvG7lgDA8ddr0V0Qs6fSeh0EJ55Sdhl/XgsOy6FSujZ/yeJX
sb9PT3A3ABtYiH7R6Ims6GgeeuBj1rPddx2tU4DOHUkbCoRIe45RnwpniywExUUgfpdG/Ij3eWme
0QPgwFZ1Cb+R833BJggeyb4prAatkfliyie4W5wYIkwLG9JUafVHAtnjYQ08UDoTtxwKBQqoXBO1
8eFC7CdMlXYlAzVMOBSLXb/GagySpBKWlpQCaqbUk5I+c1KbWAkhNQBCAXbEi8uBpiIM4gINDDuK
JXOzYdjenQY7amucsYsCrdGVKLAELsAW+FcXw9dLVsiJsp27Ttj4tmSdOs4bCfiDaUWjJQH8w6qD
ctCtEQaEmi8J8YPurIo8/GloXLEob643xuSsxDq+RIBUvQPmVhLto+dOOApZPjC9TBtPiIOi1Eag
zbV0RmSNTlMg+NJt4xqs4dU7KWqaXBK4EvGu2eCdZS6qrDjZsb/0iWATFhuwvW+5fdpHuBhJqFkY
GkU3cQTAF9e+bqjPHiV24GY2RhoFVnwMCkiOTP5Xb6HIhku/dvl8up1yy9euUXGAl8zpIhv5yYbV
My/caJ6//UXRhFJJT63OL7kx8rxevs6I5hiq0XgGulZGm/bzkHTWlfZwzfAG3XjoNexRpUwQcl/f
rEtUwt+Cf6c5QpPu6ecJ+RjqL6ZZPwO3JcJgTAXctilmuNx6VIIfYtv3CprKM/9w7lQIRr882uqW
lEktH1sjk4QIPR7DoAg3g2iFS2VE2G5l5hATJZyXTJDkZQfJM7RJL2/iszZmfTdy4P8Bt19A4KXi
bTRjAg747V5+pBWvcEsq8YZTUpEojwtJs9bN3Qpjw2U+cfnMEO6hGl2wQY1BGkH0OxeBqwhFanLp
phrpD0n6vd8DpAO2TbZLcHYN2PTaYzeshmJ6y+se/ylhkb/fT0FQQdu0Z1a/xMhIHmzwVdwoQ68f
4Ec+wkZ0RZFAiznMKHKbkXH3fIZ0Cv48L3ty6bgt9gkcdh11iY5A1cZzyiimQg34gufAS+l9dHH8
i/NjAxCQNcjmpCRTcBqK22eGjbEp4cuUcUVDMQPtsKjhHaTqY83vjl7+68kvEde5ZEqfwarQi20x
aFWBhlf1d5apqlq++eia2qgM0hJHO3DG+ZHNK5rsvTwDEQowIIKN3DRCBmem/tbSHJA49Wqp/GvT
ryrvkNvJ6SJkyqOfoyA3rCjf0wMkO+9+r8Q+/wNNmLFBf/bLeyqgudGOjcfa5QwxlBinhTpUjbYA
llX1vRmcU8Ag1dscnNhXrzwe13wnDHO4A7E30gQm2kjUXoPj4mvCjPes7ZQlc5LygOzv19HVyw8C
Bs4ByXpCXcaaSDf1kvPSqjnHtopBt8cspEVFnB9cLF2re7ZFs2GjpTytAZ62RWaZU0k5OL7ENWJk
pwpWzsRIq21i5kzyqfA6oM3CyOhDMnWdY8rSy+GUV5XPMA7LjRhfpKdvtJPOWuXDZb5pSGEbXv40
4LB5OP2l6ol5o8SKxjM7U0zIxZFA3lJ1C0pQywLBkbIXhs3Rz4fLbVr06v9B0bPhyS98DpJ8gDj1
sD4fqm1tXncyvmaBSIQdFfHgO5QWfD9jqb5dZw10K7UPrSWoErIBtuw4SmrKpPrSQjeq6nIUgNXG
+P8azQ486clIcpqxE8rzzizSIIieziTxjTEk0UGkcvVhnBzzRWJzjRbD6CAXlu0plFnjS3+3IBYH
jLgE3qKSN+gWBDizFXiCBj9KU1ru4m96uO7AtD1pU33buA1NABmHAapJysArZP7+mOtOF/kD552c
0mbcjDOWMl632xsp7CPiqE9c4LxVjlEtizh4Dr7gwuOz2gZBvY/uV/642ABL4j4H+C5twmPjbaKn
gxzlDasnTyQ9FSgC5H4zLDmFQNscHQ7oGyv1F5JcJpV3ENe9PzGCCFHArIChoeYay7FXZCKfGQXz
5udsq1y1mPKLGMBToGqc/1OxZyjYytX9t8Rq6WsB4nr+x9Yo8XFmdBqo6QSWMZXm5EkzhiBtX95k
b2aeOoGZy9V9hwE2/ckhBAye22C8oyiGvtiKNbyIl3RMCSpz/oqhnkz5z4OU+U13YLxXt0j9p7lQ
4Pg7YSv5GRPPrzQ8J5TOUiOG+eEVDtCVSP+ZmNB0nxa2NG2sbUuNiB28JeJfw5TIoL6tJOEtlMAW
9G2IPbvEZeLllk1wqdABl3EszQJsTrBQ7jRab4ZvQ6xCLTtJC4pyJW2T5yn4GAugkN8CS3AVyYp0
lSv2YRr/rHduorXiO8GydlA7TAKOHq5WAze0rhCVaTpLRceU5AbYHtWL3m2KBeuqsju0x7SA+mwu
08y24v6YoIg4E1tRXVFGK/X6NIxvAqH2bl7M5SITiRPCw1w6mZN3sU4YLqRMcQDxhP/HQihojUy3
xi/vuwjigam4qtq9FPrkTI93fWXUDLHMerDwPbfETKiEsuh5zU+kRC1v10TYWWbjW9ADP9Xv+wkZ
t8JV+fU/kfkwzGHxf/xn/f0I/Fd6/WrizUJi7T2mQ4/RkKyDnhLnMrWzFzV2fB28tE2/t4Dw/v5V
ybL6tozzSUvvzQEdyt6OHHgPQJQnrwIQ32YfsRoMuYjWZZrnBOS2At4IlNaPGnurlHVw5kqRNOiZ
Si1eZo8cRMQY2mQLgtLU0cbDI06v5bYSqJNWGUqMGuY2MYfm4rJsoj7m0X/LRORe4lL8Ra2qUKsJ
uwGDcOt5pHm14+Jny0DEZpKp+5qRkfkmvZb4ssCCAo4Cr5HGcLPyuASodYhFcUGVa1Hvg0+1LWaJ
uqayq29tf3rMe3DBm4qDVBxWDme5uSWfLj+vYB7AchOAb8sx9yQc+GVJTgv+hTdXJ0ze7xXGpCQt
spDRBO8AHUSbN4w5BUf+K/4Tj8qbQryQLpKZ5G8RuIZxaF79LUdynFzki5yvIOy70F7Gr+GrOiIT
q1n31YTH5MhS6f5wBLiVvcdLDTunAX4o9JreCDTRaECQlLgtVQRi7NO49p8fwD6eWoexmga3WlUe
hKuiqQMrZZdbmvqBcoLUTEaJEk1UxWkQVIh/himGze9TuM10ViksLHtPF0lFtD6SKe/4ktEE2xrm
QNLjm9MwVLSHxOm6BTNhkf0+hTow93IQfzQZZw1DFSXomkg19rRwVQd4ayOT0fa2uhFIdoKlkkeV
JktrMaIDscuw8rTabKYVJybtRtEV7BPm4HwEuQbJHXAcP5ccIMMKt0YlAZXJSi6TfQR0dfRNX9aR
Kj4lKJi9cHZi0Czk9hlnzk3RU8y5U9NquHCXntVAXymp85eOHfyz6HFKUtBeLeI2cBw7eOJ8jtAT
eeEO9ern1Lfa+aD5gp1GNwl2N7mOcCzvcUhPPElqcdIybuB7HOVwKR9MTi9ZCyruYq3WYVZQ3+6C
r30ms18/ShrSCn4qDDT7rpFGoUBG0qGva8U85kKihkjtqPNMI1yzqbSQj2m3CzfV/+2dezaAiugq
CjsOhc1mYWs8trN3anls7id1FwiZLDyScZLgQHBlL4s4ZMYNCXcM/T5ZcPeDZPaLATIBErFCeDEq
vpNyWAJcoVW6a1CX6TDb3wz4Ys02Qvm2pNUAjqzG3zLcGEreY0bys92HaTUwkjgp/kKCbkO19iDP
w8/fr+QmK6E9e8IUomk2CDzsljtS6V410xVNOM5bnTYu52vICCxYk3LX3xI1rTuNEFeiYt9+qoFd
DO35BthivPQt4/UfqvkXoaP4UxXMZpFzpdePZJk/NGgOAmEgOT+69u6ppzacSyMMpbCUpBHiVeMi
xR7d2GciImuk6o1VagdoRWWdOr4eChCwuAeYyyoyaPgIbiHEh8cHInfHMYR23tS5EsF5K0uIGIlF
2lyvPSAOZyhdRcyt5oLAuS7OMKyk4BPAgB5M8I7JH7D1J85LvLCS32JQ0JDoeqM4ZLofaQ7Gg1c+
F4TbOKTAHLjmqXsbMWawsoK3Sg3ZTmJNCUvWajJP7vypdOp7ZfYeoRriNQxgM78ssAR29GfoAlRa
NUQECwj+ird8Co459juUqGe+4e39p0eIsuV6EateyiYGf9KW/i8hivPWrlY/Q76TyIyL40DAG4/H
JsZ3DMUlzwPDn6xq8a0MMmuaTbt757IKI1ujpAGodgS/VvtuO7D2KE0J+7E/6KBoroPXD2te5tDE
i60BXt8DireQLpbp/e8Xt2D7DPuWNw8+YPlqZpj6ShDtShb9RQM0V+0SzWxjC/GNAl1GWD/ar+pY
iodYeVMuBTljHNoBTSMP73AmjW9OqLUUiIeO3cDVU458b1yKmM5LLfMRNomINWLF80m/Vir3n/dn
g+qc/NMUIDin/TlRYyKz6uXAyosaTzIgf2WWFnCuXJ0GPyCE2h05X1qe1eTD6jmtYt1qXHmZlLTK
f/7fPk+ycLt7kPudyf5kLBXFSwW0MN3i73H0gD8GqYpmJ6lpTpcp+p5QWXQOoG6a2dd3+Yjsuutb
Jm1gcy6k7h1Jr7+CHX1ei8cJlMo5ZPSEY1bILl1XOEC4p41I8KNE1pbk0ITBmQqO+mj4EWoaccPb
pwaXaxv6+bPUCfaiKCl9iDWBpvh16yj+vnyh/odvB8vr/z7aaYLza2eEY9iiKuKg7YM22L1oqZzs
t2rVW8Xd3w23/dxFbJwM6LQ8qn1ayutxponZrhK5Q0jHA71+URPtAU6BRErkdTkyXGsqLG1SLKRa
QBTNgzQHIqFBEiQs1sT5cOTh+Y+CRNljz2llAbNRi6eFyZbteRA9cI5JC0LlUQFYFReXHcLGwlYI
kHP+BD6RVT3Y+GiUxyzER/OoBhubvBF37l26lpHUuUdXP4nvt8oJcbYiL5scfkFgt890eP5/Lvva
TSrx+VlAuUZ8sLrRy1HAAVGo7XmRCvmI0ktrdbbdgKsRGti+chQ1oc1U+NlGN/9mHkM80+H05xUk
azLpIRGfP8PQbJddnX481xgxoNW+cCK7JEWWTWCuhQczSmMig6d2/yEFcN/rhF81tsRhfcjo4Dl1
tHxawe5Jt4coJes615sqA3oAbJ+SzpdEZcCJkOGU2EObu4w36AaFP5krtS+WRh7K2E6B/yPlZ8xM
ecY0Ta9eqqed0m9rTGPsWLQirVKyjnrzVnCvVpfmXy9pmuCy+4jJd98tg3xKLAVPHtoOhNfmK6HT
96uF+N7P0y5YTeZP2ZQ2oHcoTamKXZufkRdGVqPSXg2YN2eemosRzhNp9y3TOiFx+pSENbtba791
QZ04y3Kju5IfSsJw1xJQmZs9Z8DQBLb1N/J4s0xN5WE440kCj76YzANFeIu7cUEMMH7dgpqYt/ff
qeBJiEuyh53S5HZZMJkppZh5kxJKXvhb9G+vX27kYPfZMeIpziVHWcmOShclPZnbGkYjqhmhF7N/
5qLgFt3uOMrOo+TtpKMx3rSDS9rD9eiS2qaVpe430Ki8q0f0c4ILye4PPMlNm3ujGybezwYNpi8q
ns+TdKgemJlX8xSBHCo+pWZ3GTrp8dtb/mRUXoJT1SRUbbwswNcHWdIV4YLKGzPn2fuXkWYB2e6V
z519UdZ2TX40eLFXGXlvycnc231qAsWtvOgiooycmvmgLgqLSIIEtLjJ5lg9daBLkCfkEr3afyIr
sJq1eWrlVnhCPeSMdNEU2Th6zoxL6lBfgB21Y1Xg/1ad23IB6NKAbKXL0GobHgo63GoWdrOq2BcT
jh8nLYhXgx2pIc9tNuanB2Uivy6gILVFNa5giESpO+qluHubPxoaNhsB6tgoPOqIlO5EGD7Uxb/b
2aLApA9FFUyhLjOFummaZzaK4sxfppmJjY5QexI/e/M/iPY3kgJ0f7OoV0UZfr9b6m/4BHihZOTt
4Ssc7izTCWUT3TDY0a/gr8QhE9viJfhugeEk1OuEkL/FQuLTCnX4vo2fIi29nLccWnhiKvL3gbC3
bR6gpW37jNDUO+83Z2jcMWnByGU3BZud+G9/9nI5qcJmoN6R1rJTiJwFefEXUnQQZYsUI9zCG3YA
WAWTGTdaHLl+UTtPbyb/tUmmI0MnZL/aJr3hR5J/mGI5drzX6SIMlllwww3rMqb87zsIwCkxHVl7
V+jgbSe8ZnLWbleRgTprSWa6zenr0wjf8shW6ewPeDW4TWf+M5abMzqowy5XHfecm0BChudfTwLx
v50Qs/UC9HbwGOgzv7Lk8F1FOLaDOZv3gSWKlgCHEv4n8y4Yk+Tpj/p9DiRiw1xxByQqbZ/bh0cH
7/mWgWpibhv0JSJmWZJz3MctQeh1ZJ0G7vv117spL7QGqY09yMKCCbIgpZ9IvD0Tns2Oqse3IbJG
yleIZAX/K5LJGh11C8NNjAZW4v6V43DGUhlxSK8t17aP6WNQCk6URnw4vF4epzGacMRwGpLe+MeC
WxeHO3bPaFblQq2W/o3ZrGlzbb9pnmxWndqvwZ9HDFLatIIiXTZxk8Da8TDVg5pyINKEssE/H+NI
zphOzSyq6C5tqFfCqPqrQTmMcHHqm4O19si3Sp2kn67cmzxg5+5kSuJWZvVopjRGhNu74lAxHVaI
NKAv/ibp5Lma++JK2PNBJ0b/HnA7B5z4nuwj0PrFGOvWobuYKWjGtMsJnCMeSj1lhsVKAfl3tuAE
7vn81aJuh0soRMwckzm3wWkcO4i5HnbTQmDE6+H2Yn2As31V1tk+B/K4JggNowflW+IkYm/5kTpg
ca2Awl6ITdXaJTBM1w43tu+cpBn39TqYGHRVBt6x+kVFcYwO49pj1P9jfU47Dy+6L5Xl9JFmE0ix
3er1N+NpJW05L8d9vlDLf2NoQvCMdhFq2lkZt9bxtC2zBl3ggr+zw7UwENLicXTxoi1NWKUSB/uB
b/6nnbT0fUcNw5Ya06K2E49AnG5q8/XZvVFame+mQ9aaqeDzpsQVFi6P50QfwA/QbzrPfb/b/wPK
AguD5bwHVNsmPGxyyhcLX1FdyJbdKMChXYvk6HAViP4zw2N88exsxhvZgLa0vkRVcHHbdcwVG9Pm
LSymX84zeCL6qX9VCnAI3flxYAOSB8/GmmASDE2hr12qaevRHI5itc3Jf+d2jJNNjwraWjCSZjjX
XmS2Aegs7kuQycaipgHOXP4ns6PB2BRLTIjaasd1p6cPAnCh3nUlXMdrdu4P71YUBnDgUv5/MZv6
tJGjeefWfpRUFxWfdW149p8SobyAKGZwlfKUqGhs9JkVm4wFPmEUgMkLZREIEcfVRO8FDiX3eM9+
ESm+cmCxUIUl0Ft8CSSYwAbNtYKccCMhmA1KmSaHW+Qntn5s0IGa+7sDaumrwjU5UX/xRTdDuptQ
L0TmVayGwObdBZL6L7ghXkhYkxHZuk1j/t3YeGUvmT7hr6XUC18vXjaYt7HzUIsqUtD48oolSz4J
0TEf8/HVVJ9L1AHV0O8DKCkCUp18OQi9sizWNvfizGlnSTd4GB9R1EZ0NSDfnjCUhSTH7Nb+ir/d
VlAbRvDQNlvjARaca6eu1a1oE17YixkPtERZ7lSpAgizYBK7+Hb1S7C9f+XhVRTJohf3K2olvv51
f9W6QmJH6lhxrs7shB5BFa53sH8LXOFUHSBd4Ee6ufMj33QVjw7xSnXc6fpn30GW2P5fxv94Wc6S
9cXs4oQCdsijxKtcBXVsnf80OApkUXxzWB0obRIxeURlsmi362bDMizp4fW550Pcw2sMskVaPoam
f+9BR4wiP6UeMT5aC997CWb3gznmgJt9x1NYm5dM3n3G8Mz2nuFVS1G/w8GOlDFBQOP2ShApf/Bh
vI8KbPCNcfADRpBIdMSkcj382tteHVW3CBnwQNo93yJfJc3bkPcn69ESRdDPikxmpNXUYINA0Bec
Bl9cZtYuzWWVGQYMH7utGt/gepDPfZ0VRFps2e/1EGo/XpF79rbaHcn06/LoRibbrZOubvv4tkRw
9mAQ2mbX1/IsjqZJIGCIBLpzivXk7G5t5P2B4n1UACDOmr9QwKck723r8SC76br41rKOQPwH9yUr
641lAfr1ZTJA8uE/ReWfVhk0xCKp5XdEFUarx2RBjQmplhhDW9gdA2+PNZ4Mfbgl4f4kcUzWR//9
3vMpYhW21WvIfWy3400pmZSsDruaXtZtWt1rs84a7EcurrbmW17trDjd1noA4qakxJ+IdzCs4DLg
yynYD6c5sm24zkW5ol/XIP2r1moLWb5Yf0et2/oSzbgm/MI/+qOdXnL5zVJwYS4T99toFbOTX7GQ
mrVJSiYoz1iEkfg6JwUnqjHSGm/GGEFitg2lJ1jb4oTlkWARUUN21SzHwLQc3D7sw2oUXq3BjsyQ
8LlVlxMSjCvtzf/t+i7Kh+bE1I+SmispiiFgf7uL5gGMVnXU6psQywqSM62wm0gTkbh4FYO+Err/
wjahAFGoq5uYexLjpF29+8Qzll8R8mjfHAXHcI4WNdLWy3cd1Kubb15YZeO8Kl24niDalH6HBNGx
prhRhNWcVBlhrIAfLUbI577mcTb1t+ikRFd45k+GVqaW82kvK/HbpdtKJu1y8ZPUUf6aaAXmoiM9
lxPhfNDNQJrIKsEZHtIcGpec2lXg2VvwbhCaoe48e3KCSYpbgDFwyevhvfEgjDhK1kl4VQIcOwDv
bZDSDe6dIRj0h1PqzKY2pXxOxxBw+Ak2C+XdpY7SzfdqpvE8bWbfNQHevBxAAHJqF59oAUId1qum
Sxr8O29i0CeqPerYNCQGgul1he8mN5b2wW+/v+wrCAdcqr0shFszS2scuwQtjjv9+tOiAPFgNbjk
IeQCCxiyrSV0zw0d8eWQPz+7RyjLqZjbIGyWRnL9N95q2QU5NwNGwZYp8VYh5zhV0Rk1P9/BfNsf
5Z6O0i8OxLATfeYAmDCDUe2INw8TJhXcWGAaqPyx6nQaRf977jkw66G4qAFlvY9Y43Q+dtsAzs0U
aZv1WipDpM1u/OKXIu+81zKOUzaqIkYnLhUTfzxCLOdUBjEpMNWFEF/u3Bmi5CT4urA1pPS0GrgN
5mc1RgoGekU3dbu7FJjsb+Mjt4lrajEbk502np1FIBEVA8S0OzWwxkDAL7DsxaQSHIdAgWAR3u7K
kKx0I2hou0cdJjzE9uOAXkQcIstfOagJuiubcaJPdvhGWf3JYi3TECqjbab5oArIW7K72Zf1iYUD
jUcQWrU+FSJUHHeP/67ebScPuHozJxRPe4OwD3AhGbly/82E8s0L2Fa0L6xkBNYWc/pUp73Drpx4
C/oOcovPel8aAvrfKUEAHO6ry/KZIfuBXgMF14c6iDvxmN+AvVQCb4ngQ77MaI9tDhXPUprcV6O+
oHneDbMWFTjUtUUoS5CsS3Rm6Dn6vOwAumAxztlwoILFe/QlFly4nFlu/7HowJ2q9uv/8MaUp7E9
in/oEESWQ/D5h+1xv9UXoWx4q6nIlm+0u++e9c+t/NHSrFxxPt2bzBUBa5ODpjoQYy6dZfjsG3yt
4vm+RKnAwlP7SwXP3jq/P2tl4Qd3BSY299gQs3ogFSgtggBDyspGBOFUu3sXA7Me6nhu5L4Q/aYn
Iu7FvaSKVlJpZbHjG71fVIBurw/bcwqJuWM2cQB2VtIrfF1d2MD3Iel636IVL7yAcvUJ+WhK4TzZ
snseM+iVgZtIWPQJzBIWdu3Taw2NNU9mtP0bEil3QKXVjjtYMv4hFrMnhF+XrcbVBp8oaHiI9o/i
+/vFRtflExFI4ri6GAapZcHgT4bIzn35rsGijQ8lvs89+JoBOpYBwviWQl5CZZDhqYwgjJXmOi9t
/PvaPA5NMuCvpA+oGzbx3oEm/Fo27kCp0M/AxlzN3gIUiISe+KvKYhbYSIhOLhA+v/0/SHFkl0Km
BXZip3UA/Cm9F+HBlg4NmRf4NAH5pMn/+4JBeaR9TO+E8OHwvvBhJoINStYs5EfzFrwdjRi2EsJ+
8pBQvCU9rHF2tarudFY6lQgGxP1VQ9ghnr8wt6MT/CwYyhREnSLALEQImdnZ1mw05QHml3FqQvWo
vmEboTTsIE6c2A50Z5yt3/FkGnzZ2aN/hrSd5/M66NbXQYUwhAIxZs6izEqjyheLiCKAw4HGPK1j
dJDntBNQLktdBIxVk/lUbhxkl/0Vrdk2lZzG+LnWqTKBSmq7cW9U1x8xEVA+dD9R+MKyy6c01ZkP
foSMU/+KMp9LSTcjI4TzwABjMlKpoh8vMZce6EVB+XWgeJDVERhErB9wSQNNTmB2CM95TliPjU95
bCFEoprgclYiNQNDA9gJHuNVMSG4Z8hi0DNqcNE9ZZXYvL1VGJfHP53KuOA2f648P/H/ViFkSpuy
DxwZvC5EZJiCNMF36qjLl8LjOzlGmLF+0Qr+vdwL5iW1ePF0BURtiqTrZ6Qx3g5FAnpbhpzXePmU
gu0plVjT4d7gFMfAPmoM786roAqIu1+MX65/piSegLfMkb++11V8zk/tGUh8POp9Zr33X+5WClqr
PwbdGzk0VhXg51VwPVaZV1+LzP9xS+ITU3HQ5uMhqX0105it7sgUyhPIwuxYx9vQlqAQUq8EZ5fj
n0QplYPrU7z9X81bfqxhCO/Kyg9i71o2OK7eOVUTdpB+8SFkww10QWv7l9D+XtT5TJ2zQypKcohd
eTYxLQG65PdN63kDA+04msqzwx0V7WDBtARW1DQVIWNE8V7KNNUfP4Xfq6gZ9YdN26/QHyD4/wCp
u9AuRxQSF14NZZSuIck5NQ0bqwZaMugPMW0zu8EnU2rbp3CiuSGJrdDLMZgrk+xLnwudA0tdTA2G
r86as3XEnmCfcHXtGo+TW5ZZHzfDLIFTssdZcFW47DBUGZAtXmWwCWVJpPYe511UqW5q2rTEuQWg
295rHPxZO+PLHGUqUSr2xnaC2PKXkMeY46OYcrkF/R7G5Y9cvF9ITgFjOGidOghbp0+NPmjsdc+m
yaI3/IfmSCoYDlxbdHtQqnBhAR6e08A3uYyd5tny7rRagaOYOkLDQJt1WB6gMbJnUXiPW3XVhjri
gjbC5o1pvWub3t1saAVrWqSACwepLDVFDyECC4iNf1TPVOCvl8XrsvT5YhxlpLEO634u0K8C+8eV
p+ChsD8VrUGV9BYi2upkNdY+wBslhfJdZD7EgeimYpkCuQNA1SuKvSy39gsLOOchPLx4QaveNNvG
shURXMiplPuLSPBPmJJpI/5gNBGntjl2m3tBrjdcsaxqpq0dJ6ME5VOSw1ivEDkFbYmtJxIWjYE9
sEU7TrN1qLJK6xMJaYPNW32YT+VDdnmVfQWvoyFvj/smrfJBFjrB09BpVmfpgG+X6y/EIJMM8zu5
Gpd7nYNYJzBu039tVUrr726oB3Zm8lwrmdJLXLPjtVCcyEWo3uuwgPGTCGkMjghgjZ2zsV1UjqjZ
JH2IJ4LJEsw2+qLrufL6Ym6Js0OlMnONK9E5to6t6iQb6CES1WSi+hkv7j8qxg7EQI6nfKxxz/1c
zndjMbQgux/1wCEBAxnc9kjXvda9BgraF7et5Z1t1EqTIddjfawAK34I1EEJf29VLBtPBnD2mQyy
ZhIgp6NjPBjTUmjMx41MRbWwFttaoKaMUenH+lnPtGpG+76A1TE3D+Qos+7zfPy5NlISE9gIcwjc
GmdS4m35Spm41EGFUpyEQVn/A7OoeXKf4vUybhD7fGWoNhhyyPNumn282F0GbGPbkhpyZr+lusFL
xJtWfZS0grMbrOdcpcIvJ9tRrnoI8IPr7y+fMTAAHsHLt6IZwct/57l1Xpmh/OQRdItu85XWH+tk
lr4mGdIPCR+i+XQLJkpL0V8V0/h7xZDm0rGVAvu2fNSsYuyDwn8zb1Ot03LorMcEEZLHQcyUttp9
Rqe4g22XOtME2ARb5v3eyzsvAQC4hb7DQjGs9cICEi5u58qdJvs4VMA+xL24HooheZeklCupw7dT
io4uK14ntzwuRQpypGQ+rV1HhfT3zAUILhruJWsz+M6fsNIzN/nWroT6DE+y7YmvD3+e5GvXRVvN
P8oC0GzxJBk2bp4rk7Nq5qemg3m5DBAYfMWB1cf/hqjKkuDs5n9FN6Wdl7NOkdcvQ2dk013cejr9
ne4rG5oPt0Dq2jlm56bVuQRiXdutC9dRnSM7y2+xC24MgGqRl25sF4fRQ1M2m5cXiXQyQWOtWGSU
6gw6W8jXX2LwgtsAOV/q1wGGXbq7vMj1u0ZQquRTdcV6SRpK3BSlgUg5Nuioib8RYt/fb2ZAlJQj
9hLwchB0MX5ns1P4FImUH72FJYvmftsAGEoQ7FWwOlLjxATqDX8TazXIMrDWnBmanCLWlAhPdkvu
S+M6xunqCgXyEvU5+U+/rIsQfzalUsZ9/bO3wcCmSva7O2UMFJMPSb6/ZCv5gMH04hL4Fj4Mvson
GN2jBiWEMf93Zf/OOmDXyzpHxHK/nYDNWG9Z48KvI/tWDe8BQJoefGZl4uAEuJTvXYBQSXz84NeI
JYlYNnta0U8TLCqhG8MjZ2Ey72dOJ0iApby1DtFeK09qzfXZqgLnQx6T77DAYlKonICsfJLylS2D
Vp2yjQsvAh2eWvHynhxymxW2cXNGVFvJrKLp7fkkL2x0sSzSLOjtmLL2bMZNs2+jspJNVsbcrKjQ
OBbq+Wl5bCcI2iCfHrrtoLUproBszpcR4457QfJQk8ncFyzIN1a+8Nb7ZFxbZ6Pn6Lfr1FXWWbPG
v1tKqXzZK3vSS2y/u22wgli3VS6N85Sr7zzUZqkTXaV87F4wN/9tw9oCeE1k0MGqxcyNHgta8I8M
NsJMGYpuqrJdcrAGDoXITzoATnI22KcyD8zwAIVkt6g1eRQyvbXE8BV8CxV0KbS4/auwVSsR+FFw
tg7NdSFUsY/LBiN5hj3fXu6w3sHoxcjDeqSXBapzEDWL+mhML1Si18DcuCiQi5Nh8ZQFHbNDSs80
WYu8v0LefT7JouMRIa/4DFDEJG24VdUFy8YD3wuQ5187LwWFmWb4GY2aLsV3KpYcszGPZRvAO9pu
6Zl/yfQdlboqf2JP8b6YBoT1hoj68R2qYrSeowSKxVY5eK+i+LqGVE1keaoc28iY9oc0gGRdDgbw
k39XHwAKcdr9RL9l732sZXkFKcmaIDSzNaqioNhwif+wWYPi/4c7K76KKWTMZnsObW4zdLtR9tYf
ZC103C0P7QPIUQ2bWwk7/GMpFIeLucTqa39dWJyGq+jpoNd5j4oI4AY3LYakUnLRr1MkAFyxGlYJ
RiqzTkDl+CrQwGIgYrgDVkd1WsJXpltIqaQsa7QoGpVB75hdReBr5iYiVNEgDTEejSKvoSywZVc9
MzsNdYPKNXwNFQEnqqzzedkPQBQdB842NRO0jkZQ+oefAMU/QvjCxzowUW6LqVijJDybFdoZsK8p
PRj/1hTJ5S8GcOtgHz+B+b5IonE87kQ+GB10ZyShPMrwoNe/xlhLp8rtZ/kfNwOGBsTi9bV6UxRt
/P6xiFtxiDOnGM2XK0v4y15qN+x62BJllJL6yOBK/PSg06dlpyy2XnVqcjq+ds2N+DjGzpg85lS3
jouJ1RLwAz1wnMpbWBu9bLIdjIjcfufWsVAmZGaFd1TLACW6ZkbCHtHM4DfAPVEbbPBStoO/kR4N
uS+CejSrWrnaQIjwQdydhSm1KEdoNxxMQgXWkcu/7RomSbFKOgJQXCO6aPkLx1BDU34NnGUhyky1
0iZeVqkH1V/oiaW3AO93cP2BgskYH32jN9NToAysYAItAM9D1sfpdNTyGv1DEHNMa/hAzZWSu+up
Ff9Gz5oMBEATv47BsMCzXBzbqYmCFsO8FcpW490qO5tTTd4ernC6YRMwofpsPoF/MpnBb7ZG0s2W
Ob0rKJehLca0Xwg23veEC29aHiH4igIM9JnfF0nSpt5qLaLLstFnv3JROksWRmn9uUPE73ruSWyN
vSMDSV7bBSmK+XG+/j6t/Ma7qm0WG0725aZJ+Z96Ws3h6MFmRaI6SHmb6dIf0uAWgwwMYX7BNJ7x
qKAzO6AlbR2OVIgDgbMJsRlN63vKoS5ijF/4XL86nNxJ/Q5Paus1aUpSOdH31rOZKcFQBf15C8HM
RPRsmrHCAGryJEAOAp6/3NB23PZG5tAeQkU3KhjlAidlv/iYxEVsn6QaMfZaqF4pE2nJ9w9l2eIG
rWEZInchclvbm+zVMcbVOP9XGcsROpex80eHY0GaEISloNCoUc1IfsRHdPswrVbv8BKR1+clSgEO
d0ED3vaZPEIh47JMDLS8UNGiCBm3qCpHGYDLkXK3eHjZG73GntcZN4s9XM8LrfDJRC9AEyV1fWy7
jFuctE/XhpZP5dObUV0XmQSx64WaKFVbyPfHZ75v5UDHuu9m83/2UKo6tYWX8oPlC7cNxZQzrbBZ
z0AsexKDdDgG7/CtiksrTfPDOtk8gFjzQ+tlJq1EfzeKM1ukKgcT8DeiJASEQt3RLiUHQ1/5AotR
13liR47CgkzzRsOq5kH8Zg8KcT1Wfsmr7Ty+98CD2Ohwr8ZwfGeCqob5uoZQLkol7Q1O0I8SE2T9
DiIGGMJkBF1dMcyC7J+f0F6fhsG7WMibT/po5d0SoT0cAln+/Xf+h9W5SBEGW1W8LS69DCLem9X0
h2VOaCkeG9brrytAQ5VIZdk+1pE+Wyymkkc3lvCz0YNwfpPXxnpuPIwtYFT11gwXf4gF1/LMMbae
68VksrrJLQx7yD228SHX6aB2NeOGgvgcRDGSsLDw8mSDP2lyGzHootPqapUAbb/pwVW7KgesN5UG
O07slPLbvIHnqmlUE8ttb9/M6i9KIh+Kxz/VWwL7jRtwEj68cVK9NsCWKeLj57IxyPLZCxq1ShpF
hJXWxpj22W9bDqCEmn+8kcZISzQHyDN6azjoRxcbPlu/+eQ0ekY5vW/tfTMdPg1zfilNn/+rUG6K
qZMzRTUQztnUbQtejTQyxqTT3o25daQVKuq/ufF24CMVVexAW6/z2KQc3Kkc9T7seN+oORdElQ0J
GnqZ7ieOkikIEkZ0UadomNV72YoMaIhM/GDd3M6uMVvcU4EUU7jxiFQpgOKE+MsbtcmgA27b/z4N
ECXbGdrxv6p87MJ3Wg+Dn+WBuHC+NahrOBe6jAkENr4YMjIiEu+6KRob7M3W5e5ZfzJjmUTvJYPU
rhpqoF6IeF+TOd/EecPyPpQNmWJ/dW7RbPFcL49H51cn7gXBpVps4WlAaz0thuJLkM6EBVLAQnnb
MIPacs463YuQyotUYe2EqQGGxaEraCZNUlvcz5g8R8ddksFvdMNlETuZBQTfH/SDZyyiAiMptDpz
JPrPK5NqTFBMKIr0jfgLJv65grxreeHyvQkEPMOlrTG9ThwPiYtiqqkYHZXRf5HcCToUg8+opGKw
NepgwEKLyEp+sUektObCuYtOcchMYngSSJnsGo0scLznAoa1afUHJvuvT1cDKty0f2Ht2SmMNPy3
4sRWTaT6293dUD9t/yHczG5ha470dNeaktPLWFtDFQxAwucr4BxaKMTVva6oylnfqlzmLHAT++Iv
9cYczRytTJ1ZP3Ok+2Z0YBBiYIowkbxxI7kcRuOgCgNum2VA/R9VfpaHoRghPqDdCMZg4OPIoH7f
SKSTTqcSscKQqAjqboDvpoj70P/n2JPgejtLoAqsDjWsfD0qxWyyHZ4q3O3WXwbir5R60Y7cpy3y
7QDVagsmIV0KNvGairJT7pFmS92e63AnwSdDSE2nLvXQPa5W0Asb3ocVUxoA6mRoIkrEr8I6oS8x
GHS+aUWEeVZ6W8R8Q/zZ4PdJrncY9vb/UmRQgv/WPaSW72TsXJ21256iLprsKJSNlQtAHHyBakqE
BqcjAF299dS9eceqTfYqDwyj+K/RCGx+uvdLiyOJqAdoXv52nszUBzhKvWh4MVrqOCphWnsBy0Xw
fbLwXcoeUntRDHMwhyxTjLlIo/YJyUW5pEu4DlpQ2KQmdMP/jRNbWPPHluAzSFpzawIKA1rFjFF5
dZT3kp/c6mUTvZVqG/BjaTT5EhW9OMhFBuzKDtgmFlFFYg3IRBED3D8Vm65XQ1Bsr+xlI0JviWYw
i7fXlG8HKcvdGnbqOxT73LutdT6n/va+XDYaao5wFDRsiocFwoC4r1Qu/llkmTcCNjF/cQ6SrexJ
JLbl2ub3hGWRoFZUQr2v8t65Kx0emSWdMeNJ0STkIFdFkeJZS7maUZqwPvAsCBIWYtwyLZZu4WtE
neVbOq8FOI9DOdiOFEoyMjmNBXB4uSi5R+nEvBJ17vpRZVW+Yz1pPvhlde+0bEO/Jy23HvK71RLo
oxfyaiDgmCru874rO0Euc2CCec0xMQHRxZ1NsDNSWJOwTvOqxjNc54Uggk3VZiurR8dyxAW0wL9Z
z4SXPPFXLS0umTPaWVNoizdoK099y0+sMEgzHABfkiOrDcbjPSik8KbbzA5am8lH7sTAjgycHd/W
+9+1/18+bXwB9Zcd1QbfiYncuAugHS8zZQxNbauSjuGr6+g964zMmjS0isrgFiBT5YAlk2UlEgg6
dMCAoDlfW7t/S54uuNXg4xhyCJd/hdQ8oZUtFyVUZ2jK7nXWMcdVBxOze0No4UxQgNG89TUes1vI
5adC1+eR/m1MUdziDZHvzG0m/V+o8MbEl8gssP330LuPkwGjdFddgE9eDmSnv8s0m6g90Bn0rvZx
0EFm0w0rK4zGch2wzXhvVqyMTRVq7i92ZnrOFz6w6Cyr5UxUJ8ohtPXoIen32YLAsAefeBc7V+yS
zJ/8LelPq515VpT03yShHmtqCVRqnbEF37qTx2RctNdjnR7xEffFSxAYgoNTYJrwDCUET5jtWnLt
iWabvCulTRmRoSyoOMDL5E0KrYYDaXp+PlJ3QvM7aoBXbRVWJ+IWBeE0Rpao28JAprWEBWrRUkuL
Nh5z6pAvWJXVkJKVmGNWFuKfxSlvzsypnQE19JItWntjQg1IxhVTy3P9/Cc0naIhgtJwkCvG1egr
xN0OTaZjf/lzeFAfGReBlw2mqeJNJwpq5XzLXwHF6Jm1qc7oI18ITt4DaqwW5pnRhBFGmO2BZRBE
jjjjMJP2BjQrc9yQeoMDfUtzH8FqQSwkp9ORdZYLCReViD5ebMfdl/QtbB1vLIKgywTaz3leFnVG
OOqi9bGnVgxh2tTcecxQfFKQkyvkth5YrNBpdi5wOwNwzNwv1dly5aLp9cM31j/mpxiCfkfPwsLM
KivIUq4fL3z4kinMIWZS7QcLyWM+SEySefcRKpBTVsOdmQNGMP6hcOHGRFQQOf75766AEUAf5EFo
6BqD14xPk+1XUXoiRPGT3BPXa9jDxBeo6aEEyVBhSXsCR26JVuJOfcEILhXjnxt36C0zFwa46ZLS
8CtueQ2390HEZUqsMYwXgr2Mcbb/iDt/bqlJ/sM/y+9wCX1wiAQ+mcWmwHGkgC8BOU1Mb+qn52Sw
Is1GrksUjkmLmkxFlX6miYocBy+/JWMTJM99EXs3+g9iUH8Y0oMiACse8ddsHoczdgi3fEH7Ocsy
KVsEbSxC9ta3Ocbe2J5qdp/F5R8H4aojlVoLlmKAQ4x/tzAIlavOxj3zBvI4TZDoj/TslXM5ngke
rFi7LG5LWEpq3an4cRF/XYYWJMqZNS1q4T4srv+CADVCkqm2E6Caac891+2exB6NBN7oasx/f/bo
UJ5yEW+UwqkOryzrySUQJNxt8TEk+xqQlwCK5B4ANes9zm/OvCzFestoHSIG+ib2SvYxFCTHzwyK
HHmE48cR8WRX6B6WgOFsDb+wh7rWLGHZeUXao7sZCWebP/0ZQUrsZ9HENDREX/ZpxmNXezw8dN+p
mN+j/z2UylOfYnakHqVfOf5R6zYqog1QlEL9Y4GBazWkFVq3V1D4KVBOEB/jjQQPpT0RJImSqCoX
27d0kcO5uf3DOTBXJTMULetBS/dGwXxzaEI+gtup9W3jlzh1wC9cudMYlsLel3j3uqFUMzITX38C
ZGqVVJ+9bLewBxWXX7DsWeMG6aDWQ5QMI7WLqSq52/5vQ2imdfQDNoskOADNKBz2WePEqoRGDnQu
/VxQoTlbIfYvHg4Cc2Ykm2jtPtpxcSPrUJUp62f9D7luhAa84PH0M4bWV03ibIuBiasF5edq9m+m
pqO4dECnwl9qF58FCvXEcDykn4CdCRO3buYf4ZaiWbHnYr7psWi5xAQGdWBLbeWZ5ZrihJ4AWsO3
gPe9VGrcVcu0gCEKyl6V/uV1Zv1Tru4BkEgkVmx/eZ4JGDZn1ve0JebiGMgSGaWJHWOHxnR9mGy0
gQzh7AdZbw04Mo6kJbcyFAb1AWNJVf93miqdis0VzW9blBbK0GNykVLaeGap/KUU36VByjeQuh0l
e33RIbymjzq/OYSGRjp3s2OoJ1VcKm+/ES4eVdwJ7xhsb3mp/2f0vHJG87kQELVxuMJDHKVFnSio
JNOZiJchMMGw/MvXQS1MBNxZBP6HBeHknwJkOQs0P1mt1OglZF/xAbiUgBc2Tbl3ay+FqtP57E2l
QpDtNxjBmtBUgihwk9Ay4rO0ccae0yS4njF9m9zWAcem25bwdHkrAyaAjxvok09nTAp1dOmromdP
/karGXxbq6jROvjoDDpRiGauv74rDBs4QFaGcev7OJH1PO2j14gNXZzIepiB63YCJQqp27HKqokz
OIEsXdRLAfRpn6PSJVjAKRjTrM1C5fnS1ts8Oyu3A9q6rh9SpqyCwQrzFUeNUE/rqLObFRCCdR9f
isW9TosAWnNRHLIdja6i/vWdM/hmckxfdk1Bs+kYG8qEj/nCnrVkeu++bk2lt7JqhfeE8cZztmdC
BnTK0iT7S5RNLTJCbhYKfzBt1xFN8001rIHWlP3X8JwWaMzDM1mw7Sg5d5TkJuCpUd62q7w3BNPV
reOwtCpVypsjUcfop2TXFq0mmkqZkZxg51BY7mup0lnKXVAT0LC+eMeT685Tze+WexfKf2hHn2db
zKZMpcZ3C/ND9n8EM6uIXFQrAO3TOMMRDU7N8OqpQ2nYb9uqvEuNIe6+R5GEtKA/q0oJW2pv9V2D
ChVLT/6evXrv5zaauyh5zS87+RTujIwItFEs0rovjlGbGJEWRV8js3OkNH+ixFvfgO1VZMFK0/A1
KbtVr6D8dDCSdVryO96FHP5NKvodeKh5UCNuLjWPCQEEQj0AM5CpUdKbmZfX7J7FdDXHOdV4t6Uc
5Qspgmw9zUeCIDDraDKT1SMUd3xztI3ZB4ZfIUVJaHtsVNAyppxTax0Z5FN/5GDZEbotOqvz+f45
0W3Goo3+KAJNd5cU4F0MH1rMNZfwsTJcI9Wxr5C12Q7+2d7zEsAnb02Csj3sNWtPlUNFCUFfZZoP
NoUplROHOLwLEOwmFBxGvGWohHEt6tLnCx9Gk3LV2WaNfIdIDcpnmgFpcT6JHBp5Wl+2sughibPx
H5YAnapErrflOVVEbvVF8k+p6dEsQ73c4pQ6hUkaT7+vPrmPOdPCVoTqBec88AS/wIfjKH4XNrDr
uPC45gYuwPEmholpHUFL8iQO1NQXMjayjJtR3z4LIAb2MnKCSlmTOeUWkRYi+Ieifze+s/08PS7m
rwtUUJnKjvWzcUU+YTxraYi/JPFHXDNUkvhSyYQHnBINqYPg3+MFjSlV638afJMUO9VyJjxLSQtl
mqgoAS6Jwpff9XDPXWm2up30JdcNbOqMJgd5xK6gzWwooR3tDbbbDsJA2d9fkDivf1XdiUL94yB8
Bvkww0Bggjq7wLTLzH75hjVyeFEZCCnG8Qw+0XG+JbpEVNOezV0g43tpZjcmi8YWRXbSlaGQXTFY
Vo01D4myL7dYR9Z8+IpSYRXdp92VpW/c0clG/kKbd6DlHXFpx3Vo/ihNk0ByWiZsmiOfoOsVBszG
7xKibvxBYBQXZby0KZ6/cOEuprX0ZpL8NnmHxYBDAFrnfJuNZoz/ztZ9GX6+uZlMrF6r/pe76/ss
oBuifqBXJdNIEI1BkDv3HqhtH/Fx4Y78ldUg7wymuUX/HRKDkyPm+GWUwZpRrPK5vEUv5IWaQa/+
q61/idi8b8tvJR9f+XafESzuTHNFxPZM+Lmv1ozFgG88O0bki7vs5ALIki8roZ5YsYmHxh3tb20M
Im7SU/WqPLGZErQIIHLRZpXIw7FgTUIicWd4UaUkGDMzqz9cXpwijQYWahji0iZFrv0fPe86GV+X
sUXF4uBvXbMBu2/YxBw3kjPP0PshL3YdKW8CL++yzNba/iDcwKXsodm2h+llpRLicLW3sM7C4Ane
6st4SVYsvbto7iGW/4ItPgLnyb27q9BJc6yVMTzbcNO67f4ttYeOh8NfEwmWoHiO6Z7lboFG6qgs
XkUwcFnuMNwRHrgJibuaqi5pAjXBmd/U5V37Zti6ka8+TjVFGDteYTpGjShHqUeQ4hU79vq61eyD
LmNw5zp9gQYSIG1nCumtGyu5/DAM8dAzRsFe7cFM1KjvwTKY/2W4i9osuk8GvA8Kpogzl/ZGmkc0
1MJy7cfWJLsYiPb9zcFX5S/qBAbZquIxGzEcqEJ8kiCUe1RDxeP+578dd2fH3w6SuJxtwnbkEtTv
vfKzE/Q6rEnZDnAd317X7HDFMzRCAPx0hkGO80/8i1d6Ez4SLwiiny0Dfvp8B3zW/2DrGeqhjPXV
mMJDjdRamuHLrJB83d4H81YbKfdY+kX7V7ObUg44So5TdsMu+/8ywRGtEOSfHmazONSHvyRbOzhM
rdkzF3t8dXaXIe+RK3wU/4eDySWDG1IcgfH12UT4RZDHuSETJ56sQEkBR63dQAAjyo7X1tG4QCfL
Vuj7mH6DkTuxKhD8GqO6Cdh1E7pMcMAnIIaGsxf3lTlSYc5WStMaouzh1vBdXLWfMinR4N9pgTIc
rLCYigwLdJLyrp+1KNMtn7dxwguwOEyXFH6iNTzc64AuOYxUDa6RXA0SUX4MDDnojf6ZTDE1qxPO
YZOYCYiSxEXt/J0XbtEP50xf+aF25XqtKqfgq5RUEaRJFkHQJsiI/brrVGnoG9HYzntFW3uCVp3G
AC1Ph+Vz+Pvoh8PHeaVYVEYNVBDUul2BgHsSNgM60htMVbUhximWCILJYpMnLGNTR7El3f8cBkmo
hb+IkCZ1ZfU58LCLKQc5CrKoVRkLLUwfFZNKJmoxIxxfK0YmJM29wP7puPxuCULSE41IJ8hOYuCK
WT6QqK6yk6y4rf9rUkO4OHElY6DgTyKJ0/LAjJwFr5FU+oIwiPj+KdNg+J5l7ypTUEWzVvJT088M
1lgsqVsxKZgYjpOmthl4Q+glVfXmhuxWNgdOhRMzrZNpHVJzpgHGxteuAB/zksp7ZHelUDvvqs4S
j6xXM5W6ScrtSM+npJ4jxuO0uUq2VR5EF6w173p1vdz+0UR8wjM/q2qQvFHNtrmNqaXktTleYqYy
jMxIcc5u3vSLGyI2gGHcX1P8l/hl396SuRkuu8akYfNiMb64CpCXInWaPrBeqr9SKplg3zKUG3Pv
r4S/pTid9ZwbMP3zCamSOR3RmtNCZQH1fOA939qTWjFdDsWQsrr6w9bnd159PYdATn25aweqXpH0
tK804cHxRXdNlsowvdQUfCU0LHbg7XUmUPbs0m3IXLm+Szh3FZwZtxWBQnev4UBGdT+LkY3ViZOL
5M0DMhQ7l9OkSaIT0vKlgakekyPUJWLezm+2XGZ6cxJSsPsjzf32/ENYjSQlRSDJzBlbA7aiNBGF
bkGVZ2LhqeiBJH0zuYYlI/d45l82Wpx9r0fYS9dLIBu85HsIEgG4UdTtuzchfrwboKbMvpZJQEB9
kQa599D4+O0bCHLCCP/2my/9MGcegSOt3DKI9V3Cw9ezoKrKGdNini0a+R3jFWFN0uBFjcpN+7m6
VwNjY8ZeJMO0tmqtKJ9d/CNtHxKMzxVNCxgq2fi17ovtN56JOsLnDrCCks+YYKJbhgzg72xqd1bX
W4vJv3nXEsWVVY6DZzvc3yONWKMW0iKwoNrYy5nE/z/eRev4YmvtVv1utE6gkjA37IJFy0cNgBVV
Y/C5uJWOs7n869tDlfmk4VZrMtc5BgEJyEQFTdp7HiZ4Qdypaf6X8ozy4/yRBwNUQnHitBziXCEl
Oyf/WCrfllshPbPrM3bpzcsklOUvhgxG6lNbdIw2IYxQHvIlWNJ7Nl7ARvpWV3vcBoeG7LAeYf26
1UT0geNBcDQB7F6IFhGE1FgvJbqTMnrfSsUhqH2A8wWQfB4524uvkMrAHWjiuaZkJ91pom2D4PvH
z+xEpb2LVbTbNAzMCGoVErE6R77dJg51LQuMyezuM8Gh1R0yto6rCfN9/Z99MHAQdRvlMyc/NqVJ
BIqVrUCbIeqCJF6sLuonRlHTwb8HTwjg3OVX6NYx5FVM85ITBV/6IP7FgehB7/ZCs/iyGrIRoTqc
5gPSBqmzmNhVwTKgav3HzPNEgm3W56sfRtVZR9d0xV4qNEvt8BGGeqT6HOir0cScD1H/XDWdGimm
TDJLhNl77W5Tk3g+fuc/DRfN4dQek/S7UOGOB58F035/hDgVdgF6VWiwEqEw713TfOsNlVSAx0Wu
yIOJLSaaRanIORYQ0SosqGXyB61/p51njzrBgAQuS9rBGWHC9lWj6QrV6lf1xQBZGb98Q6UvtgCJ
JP65XayDbidyQoJ052sUnqWwEOdR45qmCxqNS8Y0ZM/ZjZlJ9oZWVHbvQF7W16hjEXbqXlpGu83Y
zZWBL2Pl+axtKGqSI5orosF78STRZM+x3zQygzSmFb9jJP1cWIEEOChIl9bu0Vh+fZEdbVPZgSju
v9+PpkrG14Bg8GHXymr8LiX1G+hzppzwcJlNqJJ3B1AardXVVnTcYzk3IPBPrF/YzG7kalW7F4VR
ri03fQWSqTmRpFZmxs0PFvej6lfqHIAFU5uGOBFPMKjs9CBYSy4PJTNs0erGQPRtG7xNwLNJRW77
TEyl6tdp2Z7fx/DmUGq885f3eLWEUsy4C2Dk0RnbhSFRga1f7ybRhzMPOrcqPtKwicInA3+Tnune
UotH3M14ZfZXQYBALMLHjTpdY+sY+WJCiRc3/3Si5+xlIfDL82w/gLvk8oH2wGJ3lrNJTeDrwB8v
jgf5VrW+8RW8RE9bel8HN/3xtD4kFD7DXno0HpUwFslTB1jbfkxY+2VTd+YFqTZnR4jJvwFuPvTl
8VsI1m7+FWuuuLReKF9WSENy0+3QTh9QAqu2O0Lftod5gua+d6p5X8NS7aqP7ke7BvhcO0lO/UXM
Or3bfARJJBQP1n0ac5UB4efKXTrW8YIpP6VfuJXeulWDB3Ox7nMU7FIEKZbl13KCNhfgNmiN4GIY
qXhVS9xlieBMkll9WcZpTo5KRQenfzRzl78NueaQgv5O6sQZ931cJ97GLCuOfco0F+MitMAXJmqq
1LT2zznTbFpyY+x34l7YudulsXrwpHGxh4v+UHCkK4qFftk+HBi4/OKyunX2bob+eMwwgXCO1AJX
p0l8c+yLy4uzXZvivXY/JjMNKto9Y2VylA/5qCtzoaoCStByuPuu6gDEXUWkIILT1zwtfNAR/8/W
KV6YGnw0mrrpikL11dgNQFmR4iMTQJQvXcgfVjEsAHvVdZ6LTq8g2GKr0veo24tJ9CHt4D1skFzt
5ZTjiTG/zc12IehqdDqeBmRrZf49zhyMEfLmzSkywNzB5XtRNIFVVMakOmXXPcT0nsGD2yIAVtBO
cckFDDFKYcNOyo/5NmySac4KVVWgHZ1EqA+FUkl7GZVj+gC3ms1synqwJ2lbMGIB/ts8k4W1Zjg5
yThr4rKe82Gl0TbX2IzitVXzgWBFpdY7hhYANrxVPrP9vqF6gKidzhOljpTszG5RFU0fOHUsJu7Y
ZT4zsuuPH7gBu4MGMV/bwApwvlhl+Ug6PJQgu3I+E/Lb6qmH+/X6tFTLlVnbN7Ncs8k9Q7bu0Cy/
0pbvJ8GAvdywkYF4LLD+QI5Cl3Ef8sFrE9csdML1pqzNtcIjzK2cLA8V17jzchEAKxON/ilPQUPa
ONRe5rSqeTDHfuVs5m33VRIpcfAjbnml6ApSvjPtlLviHqPP6CQbDdu8dh/UazxHKVeGx8c7Eh2R
oPfDqC5lisUspLUrW4inZYXe61oD93yF9RjVqlFcnzeWIhSjq3pKfWfZfI6rePQp62t6cPdFzVom
qyKv728E33I3yGpOWxUUTNBmz1jJCyKGP5yP+nlTdVWED0XniHOSruPawUtPzmLBt+jRY0ZboRrs
zwXAPRwmdJPmb26TvJllgZLOm3x+KL3JuDqiHaxcvujg2Aus2KiBNkh+NUFmPo8NNWUxBXRsivrm
3/ydFOjvsKZL+TLPljfTfFI5ddjy46IN/h0NECkH9qCgEk8Y+yQu37Rg8eex7SQTl9j3BjD0X6g9
eZFYn2MSDLfn02WTBeISN2oEBSpWm4QQDUunaJ8VZOLrMllsu6kPyC7lgQWBsjscO4xd6umrzbtw
LCQe0nuXhpmgUD3EBWsZextX5iQUy50MnnwyL/OiKwaJIiABlglOhmfofl66BtGVPEjCEC/w5/QA
wwo2vu42HT/wuBw5CZUEXRAg5k66OD/IMXPPWETniinkY9WGaP23/vv4fSgMVGpAeb6N8TIguI7w
Jp/aMPjIx6Y6R6Zz/oyec02PUHSefv99isVzimYLrtQXZwXc7k7mMw7/UoGApP317Z2VFXk33Gm5
7EN7pYpr8VTMVUS/y73mXbL1jAdp0GkmuW0VLg5kW/yYSM5Hg16xBOO1H2OT4yrfB7TmXOfA4QHe
wLQxOb8I9CmBZStgYvEOiiUj/dtTtNjT2xAC1NiKEtzplpOBEJ6TKGHcndUK4M7GJDd32OWXz9B8
mKzYKpZMSwrpPMnWTkhrBhdxqG7Svp/eNopXlxpEBxbDD325KqPEgxzIZQeY8hNDVlSMqwwDec9R
PoZtQEbJvfO/cY0ykiOmaaJKOzp4qS+JCevcViUHjF7zSyMsPV+ar+9gqiI8iAV3ifNLFBTniJVI
GhSLxakPRS+1Jy9BapouDqDtHUi2uv7eCT/ispyU7mzK6Ro3Ql5KzYYenq2fAbKW5foAjp4z/4BH
RbwSISifGO0bz+1/zSSuMZGFtNRWVwcGgmUFCxzsFuc+uD7WhTeiPKjbofQfl2pmlaR60Z4ecm11
FfFJ0SqCCjRFhpzZagueiWYF3yffQsoCBhFM7Lly8oznSUr3/x90nQozHvNz/1W1Y/8+9MfLT5HI
25DbrBg/SVmwB/8/sdcYhqH4oEBT+uQZVq5ktk5ZDAH1coggh4kRXN8Sb4l20pNZzz2NoGmobj5L
P5VjQWzp/cpKXIoWZQhz71lWb9Sbfn3pO01cFdPVtGJP2HxZet+5fMIzY5av6oXf1ek2aBhe0li+
5DzkK8onUTAqJrnk1CZ1L0w5uDTCui+l3cUG7MFcvLwKLejbKmdFeUM3ntNzZWeMLjrVJjNqFlPu
qRc6knKCFlawIc/0XtOhYpIfAXB+1IrkcxKKD4gSvEfCP4i7x0e22bRlqs03ef4k+MLVv4925LMd
i6tKVygNHq3ApVirqvovQg7sHfIPmsTieD5K+DBYtWJUsDxU/Jm3xqBerdhyYPg2RSfZAjWKKG+N
r7994VxbPYK1le456qyAjELwZqti4eoRMJ6oQVmPK6VvAN02iAjWeyVN3CG8CTR0FbIOe2glrLtr
uEoO4NTQjXFvMnWStYYfRdf0OgivY5BURfSSGVP/+6j7iDCDtkpifEo95Roo/jB/SHl1pXG85aLt
MQtq7q0oz4xL94wKxKP59IjoZVe5X6g2sU2eBDMXLbb3rqd+meEsQxS+WJjo7+GJ+oWAvzDEyWD7
/qAXXZZGTUhulKx0sxQSEMbITmqhm55/uDYIdIHINjsyTDJ7ies6xYXN+PSXcPq55N6vnVxMFzh/
YYl2gPRfo2RA6vjWZySlZvia+JOaTlWomfFhd9CfBP9UKqauTovxQJaJQLXyF0BKN+DVRtFyLT/m
YEGLhL8TIW3lE5ejrED2ZnEe6n5qfbdpyvZVqKUtpjnXz8eDj2P3Au1SZjn2ZkP1YZJaQB5rz0/c
o8p90+W1XNzGDk0ObalTOrSSEI3C2RGex9C1eTVR6WjhxxSR1Sdk+/zi4vBZchf5aF6xLINtbN5u
8x5DlYGqPkIrRIlxFn9kAnuq5z8YV+FPDiFoQ+PgGRbQX1Nfcavz2c/VytxWlF2hj4RLeIOz+ai8
XnId+tmHS2ppb3EMa4pUytBWSqF872/tzzw4xIYCP951uCY6GbeYjaTIgYlPK1LF2ul6Iwf+LnlJ
RdmXsh5JWMzG6CBlf/l9heBs4Cb6dwOD9Oz8n8ugavG3UjzUk9yt37zVHv9bomv58aYhqEINA0Um
b7f6Oq1rjxIkWO+uvvZI3pAc8Nlb93l3QlcFHkblnoHvVqrKCKNYaN7ACuKQFowWN3qNuKSvJESa
/Z1w5yzuqPVkKGHFwlKulEA66HlCXJWHGyH7iYSAA6qsbsKo+2ZU0/5/0PMxS3aEbYTqprDzuvSz
G/qFN5z4myG63ricF9c2t7FYDELWbFJfVa1C8q42yMv6yBoZZ5FQTWCkZLWUrVbhCt+2upE3ndgU
iRy8KnhWOZESyZ++ebxe5RP4wdc+Cz4YzYt78bxCwgF9Y+KTra+MBVevXmp+rB/H9BAmXsUFNOgC
UgSfgrslu+bDVCt1mVx3NJGI7OnDfRo00cw1OG3jeXPC4S8dkbyi74OjwrmXKF7jNFUib7ZDsSJz
R0HJgnLcGQ4jRb2lmWGdyXVXcqZEPiYa87iQo0HSg5tlfN3smFzm1MsczsBreKZASm5tmWQv5czJ
UlCSf4iIpJaKGGqTiEsfJTYrpkp3yUfac6zWXVbaQImV9TeC/jEVKyBEJvi4tNE0WMzZbtm5Or6N
0BqqTBHleCyoHzgzseyqvMtAJ71TESRhMbKc+c43UMDSnP7zfBi+RZJGMbHKkFqYkn64iDAHYaTs
7xf5NpRmpjL3ix7klqRp+GgXZIHQKDgdSxcSTf2ySYYW/a3nHT/xSVWQvKTg1d+0wki3n9FA2JJq
Y59WOjMYY2ph63NPPWPpEk/hauiboLu5XmIAE3skTipbynmTgxiwgPMcPSig26MrK6QoEgDHZWx4
TFTuCzgIcVq+S3LdjvaQsOKBYMtDAzFW1MXDFuzIPRZMWpw4BOA43N3/9SnSCm87rHbQHVYhsEp3
mVAwEp23dd+JK2knhmZaE0GHuqZiu8yseHVhSdQCHJZiznhu/UO74pUZvpTz8A0t0ebTwdFcll7l
lFGrX5WuJalJf9wWkre+T4Y6uoXHj2lJXAXjPQ50pVR/wJ0NlK9DNeNubSdoqjeGhhpFzAHx4tnE
xZOUlMsCl8Ux83WMzsnW84XbaQfCJXWojN3sPnEBOcijA85NeppMryu1yfs8HzoDa8qYdv10ChHp
XoXov0EduMZMTjrl5Dmx9MYc5l0gMvwjfNqptpBPJoinRvkag6gyMlafGnLakeK03OdHfdJ+t3HB
CUzk392mYD8HgV59OB1yyhp5a6hZsujwk2MYKsO6AjiweaH7r/iqOfpBWy+1I8WFIK4va40//kmg
Z9IFFjVhBzf2goWP+X4J4yglYGofNvYd4sy8ezm36Xii1dWp5+gGmvQIkA1B/eQCifuinGBJS4YH
3vZZZzvpT6prNXIEwuTxDnC9SSCCOTN7M8/A8bdA/GZPwlOatXsKrbpYho5PjbwMVjtS1QqeVH2v
O13r8s86ju9J5seDgDqKsKmYrTT5G/anpBD9IxUmhV+hmBU1Rvf670QvNqZKT0lKwdqUJAMOu7xz
HE4fIWW7xRPNCYnaqxC5uKZHP3veQE1EV90Diisdgu/yqKqICsXhATGdzfce+HzoxqYOrPqfiQuG
22EQbzhcal36iqeygmFvA/LNROnxGsavuRMHqXti8OKN+uZvjI5XSkbxBbjyQhApLgFZGIUExcVf
0kvKp2m949OTb+Rl+6Bvm4RrchtbEfXvogs4QTY8e9Q+Qgma4oj/UXxoo0VJZu8mZKMw73vM6CBu
4FIw25LdG0lnrt3axNWuxOT7utqbhbJyvmvg1NiVxwq3aCq7qF8ZVYcZN2am44prwAFdvf3kJQ8x
72K6otTM5IkIOwwn2YSTJPTjXr4mhE2EdSMxamaVcA7QpQHYDkXnNKTQCntxvJVvcYcv7zFd1t4e
T3W0TvBJnL//JqI3xh4bxFPsW9NPvff35lQMor3/u7lmEWR/zk3f3Mlvn5F7b2NVr3uibr7xobLm
ssP4Qw1ZAuvPpZ6ol4QTw7wvkq3rC5YcivXvaxfcmlH+2DyLyU8u75AijdcmmXfA6tpNmlPGqDzo
xj4ZvnK6oNEG6WqtDcfflcuzyRUIh5gPy8ymuyvJeJ4TZG/cM7hrYSG9Mh4kYvF0Lk9xVv3XB/z2
Xli9WpZQryW9nhKZESfzNS6ZsOPwoqjyF2ttwyVNUlNmIAFatFwMdkFWz50Vsdp0pl1G4eStHHnB
Uj7OjvgO6cdnQjnIZy2Vp3KIdXknUTGia6y1Oa1Sd+PfBan6Ybq1Mue9fO4pw6+Z+2K77Ook0pcb
6S6P2BAg2WVAVDPbxZngz2ZZN3cqXqJPRA2GNA6K7fNE0pN4m6OGJ6q/ECqly1Z7JtdAWzGAtmoP
YNi9i88Bso6golhlYq4izIWRnUCwXt0FG8r9vIcW9zzUTue5xlNJyiYcP6f0KGJFsViJW4EVY3Fi
GppuDVjs+zE2dC2xYMPPxN5tBDOZej8eXsST/lLoT2Qrr0CJcKd2Pt1J5NXub3sQl+t9L8CdFWom
u4nwuxRBiLIUUfyjffVn/sXBdOtLLKVPQS+EWM80VRvTEULc4sHQy7NuGg7RRplvHNnfdjzFHs5s
s0hEe3d5DkXVv81aOnpBHL1lWjYlVjQESf2j8m/s1DcwCjNK4jSA07wvkLkxmYkD6kPBjy7Rijkb
3HUdgOOvP5SkT5pF0Iud0o2nRpmlZnNwE544TeTrWeMFFilMHWcp7sQWx10CPDM3toU5h3gymPEI
eun2Rl/jPPQ6ygAaOZ5j0p0iXWjjnWnuRqfBtwhP5nNnQEXExnqBl2eMYD2Kr1pTVActCg/RD0UP
9TH/foL4vr4DqRVxy7P0lajtnJ6gr534z0BsOv4szkAfwTIM2iPrdbgbuHhW6O/F+dvO0usJ4LrE
x0r8drAguLF0ltpioILDYi7o99Wda+SConQzEwY58ghXDX0DH5RYlXs6nhzzJvEEcukgX+XDQ/rW
se1zkBD+hAa6YqN/qmVAH4rjnNQrhxDt2rHTbz32PRhRY2tVhPRb7N8iKa75cm5ZmSvZOAEmNAju
1gVBf4nCIXP7n0cMyh8jxtb4pJg9+z+4/GB/Bu60/dLLnpn+Y9E4smlYTiuIaaXIyBrqQ8sKcrqo
EEfqekzbCFlV7NS9pXAlz/GeC3Al+AxadYZXwl4oqEFRykMdzZ1pY1fPPo2yheNwuSBYjVf7EYDm
ejJyLQhKQbGdACqpKJMF7z4S/Cu89HvTQEbcKPPrErTD3kSkCnLFoExuNzbRF9BJcCXxBR0Qvp2t
7CeBDtsaYPBG4wKxW37OnyyqFzgoLouysZYY5FTuhdP0YjG5mIZviciqJqd67CujFyENmkZZOlny
sY9YOFJigjh8DLTIgUfaAR5to4fhYJNxiHVGsAq2Fsk1P+TQ1nyWSeVjbaZMnHZVxBqK7gPy1yfx
BBbIY2gKVSpkmjxruWBiyb+1JR0yz9wHXUrEeEOX9xNfoth2WqHgVUi7i+iBvciHWxPuWB1r31Le
lvX/4RIwv6Sb152tYnyMYIllAqTzcQRQiiku8HHWnyjBCAa0d5Aj6m2MSB2qNGwXiPZck7dQK7RO
ZKSvga6gckAZ5Tt64edkF4W0zWSg3NV6FxSCmLOkc+slSlGT7q/IrVA2ir5Q6ypikVqE+knnpSoa
rKnRJ+ADcgCqDbOR66sfXwNnts1OQar1asOA3W7kuFRjUFxxTTaqsh6aZIfu/lAJyuQOkJdZKyBZ
gelRZf5vTqY9nnNq475fzzE0KN23mgN+RRYlC0BlRgtIkkz9PcRn56Jeyx4/KeGdiHnZQXpaz3dy
7JVoNs+ut0/xOdC7ZgikGQUyoOAjjdpYo1z8YDjhywbLO0nJ57iW9LvvIGAxfE/JcXJEcs2QX0qy
YCl+dCdNIbcPB22/xiKxouMZi+j+mvZPAnPnmrYmt1N3au51ZJsWCWqTAU5BWGGRmylWLx2fZYl/
sG2xHZ2ZWl398Vq5KlRz3f9i9XqOztI1EeVIF+RQF3PWwZO2soTDawXaqtTGn8GFRsMEdna4kQBz
Wo1/eSKEymHuOhjXxmQmyxEjk0sCc7B2v5bs9xoJyO8ciTydfvmQbLnJNrNzJJtBbXDuJapOS/74
6ZfCtTc6P/5U/ouOhvcOVYWzUPGxhwbqZaM7HZ2xkdiWN6Qe7+HRwjHtty/FSHJL/DcUjhZypPlU
v3tAtuW9NaAjwq9KrrfsFYWBIGm0zeEjQs0t/1FEJQ5n5MbFEjqpQWuhhlJvIAILuH/Q4754n04b
LNvN/I8ejVhPRMv8K/4NHdS9rZdWO9oyyfyYxH3JPSyFhtQ9D69ctGGZCqHw1YYbqbLla2Bq/bMP
18WUEq6gAGPmR3Tr8kppUk9LQlP4SYMO5xdLZXX6XEbIAYkp0FBQUHkHVaMEoIr8ao1kMKjWCpxf
wx4keIeXA7MUzZH9qWKgk5q76tAxDpxNe19OCgDQDmwXew/zygPIeDVZ/C2iR9xOyPTQMU+mFT0G
71qkZiSv6EPPiZEKmrU0d6IskT6FXwDDunO9EHGJVi8bYCQCuT2YhIcpx6dRKm7y6EzttOQc6gh+
OOSzxOpn8C7zXGKI0I/T/w+Qphyx7EyXRkHRfuGkIIkVCF5Hk3/CzRp6c0OKoHhqxkMPX2gc8aad
vt5DLohZ2XYqu0V+7qVIFflgbiwAaMvQnDntM/AsHDCvL4kRODjEVKFGtsVcJZADTPgAWr3rOQme
ZogwOWK/0HWusruyUpKhfKMqGVi+IZ4/O5xgx9RyzlkZkwtYVJspvCuMyQWTIDrviCn8+umPFShj
WVv2OEx2hwdsuMqNi3PlEuXRlvDTTrhD4E3bqi98TomXcddvp8oPGbWtiONfZwrv2ElhrRS1rvr0
3Johge8La2iZW6j4bto1k0ksh8dl/fs1k9JlSZfKELpkOdCfMQupAzWP0UZjfH5DIbYP1r0PwNWJ
5ZkXHwiMh8D11NlrkX4a4Bhm2dsGimVOvw8Sn1LPVJqJ+DzROpTNID2FU7hxAQm3qKeQ9ftfnxOz
9Jk7Q/CcEhESM4uz2+V5Ez4+DV9Xlx44jrlHRKyY4G3WMrpg1DGSzl/UyCi+FNTyaT2ZPaeVioHk
yHbBJeJVs6sjRCxivjv1ez0stN/CBt4YwAfc+kwZp2R7WTAbqIvJ+G3Js9heWKpeYH7nqJ0lURJI
AxWQ6y3IUQze6MQCX0jKUA49Df2ogEAtRCx1QMfGc+k2Zq+80e4pEDVtazj0Yzor5rvsM+tVFY5l
vtHqXF8L8cgvD1Zog39kBb2SlEqGIn0shG9vqUPhLKalWp9wkGzthUKbWajo8n4b9rqfrHawhb4c
liT+wRsupE6pnPq/n1wDnPO5k2Go7qSzD2AF5fNAN5hFMoBqOvCiEQp3FlybCcil7me1+zFPuL6T
dMuPcx31s8rS1HWWlB28rIeR06m/yd/o+IbVaVxtrcJmlpKOCeeE1+5xwlWFW+hpyRIsdt1kDwfm
qHyANygpEFGYcln7VMOVeFkO2ZjfPgClZPAPJQ9cIm1NYezE6kBqWlIvnsIVS58OJf2Plo5yHiPP
1QyN7Z/ZZkXMQSOvFqdPwEpAYysSFTKo+NRW7aNlABbeJr9ekkydE8EGOgKr9iTqpEQKZT3hO3YX
/PvqgcQn/aSSeFqSahijD2Iq+WbfcPAsqHU4N36HlvbdJMRMtE7LQHQX+mxXbT/abTl+wPWOBHen
PEbuXvTpaNfO+SrPoUQlOngi/D6LziRxO7Ppr9VT07AvGPgUjZeHDan/3kLuIqDjJIK5coK0lEIn
EFb0iMcR5ZpqKOFeWoEwobvne2dmfOPVzEeYM2G3Y7Nq9JXVDxNVwhcYboVqEs0HJlGwfvw5S70D
QeStC2vVkEk9gQY9k/GqHn0q1Yc2gUTwqh5/lreSvpM3sx681JchFhhEnTWe+L/Q/PajuQY8QnoT
8Hpzuax52fLAOQr7akCNPVIwRwGCIO6dSy/MDguU9IVvNPOP1QsxlwfU55YsaurTQT5KfGjN0BgS
8KjfhawKlY5uV3X9B/csNriTtGFNTMQonMsa3o4mDrhEkIwg0x/z9cH0fGMtE2jQ1qAJJLwvHlSA
qc9HQhNb8YCM2M36bbtde/aoc2rsmdnJnGGWD90o+Ueyw0h+7TN4XruSPDSYO4fJeQIs4PTMwSFm
QpX2R7VfwebP5Lc/U1nO3BD4ryLR33WxXNMImDgX5JR7ZVzbipMSi7+/34xyDmDt8A3pNYbZ6qLt
iAvg9PMxCLxrqStUR1eFRHMYKTFImNcyWEIYCSM3GntGRsCkLF5NT6YmJQbL3JeSBZrms9230t04
HsOsZH/6EhTn0a2YVSHEYeME+zxyHOgKfb+1qqfiYGoq+IPVu5Z6mhcP/SNguWMgFHWp/w35EMlQ
5FDW6/EssySfvTeypG/RZlW/jnyyK3QwkIVLIxWihaw1Owny4SUu34/re46JHJ5e+NSzeKI8gtIr
3Flt6L6zAX4u4iEh9hSavoz2FfB5p+8tidWgBJ0LR3/Z/HBsVNDk4DRJdHrtuno1cMq3wfSFC17i
yI4+Vmh4bO6OJ+DKzzoMAgYEb1LwjdLmfmNJja3l3IC/NNSLd7+nV9twObE+XnezPD18PHf0Gxqj
pqnt1/4bKvWQov+G/w6xNAAPEPSaNFtyjrznKnbFNRXE2YPZVTlgoWrfy1fZDs2cPhLQDCV/fUXs
z8EOw7FS61lSCwUILdtZST3z1tB+HPPDOhk3j/70eKIY/B/NnzpgnRo0CgKdcbNQbN2n/mFyyIZH
CFao1rIF1yadXME8m8V5V7TAEg+1spfkKcw9B45XjpIKEXNudnnS+hWAJ6eKlm4SW9fJHD+JQPBe
ynUSD5mflqHgxOzSS91GiWXd3wWEf+xWVmSTh70fd4zSnEIZ0x+wWhL6g1cdx7OERShZKZ6jT/ri
h2RGz5EaeDvrp55QFIRLCfVAaGGp4oAjDvUSNXiyNhPGqmz+uUbXqrbPcqUNrBvRk6j78WO0FRp7
48pV6rv4pMdxssLBscRfNpRanVFUnoVh0lOzruaJM5MNvtbv5j+dyGOKG6bWCwYBdnJNWX1BODhG
I/ZTfTGNT0TfuK8AZytxYRJse0VpJNuNds7FX0XGCTJVphtXmYLZE7HofcgXSqTSfIdefnVWPKJH
EVhbdZm3JwLjk+GmljhEB9gAtzo8jM0I9/3CogsZhoN0zJhPiWFKBMZHpncTNFDY7k25teZWPoUi
oFWjIzhHVrgTl+3V+VOhMy1iHPpEteQoQclbVlGB3s6FuifjelACsbcOsk4nrEX+4/L53DqyZmwh
pZjCSDhspZwvJIJv7v4ZHT/q3alBSMCEWd3VB+9ksyjJbFzZKRzCbgJ3lQdhVtRhn6ZzgqEitds+
+FiXqsL3klwzfeNGc9WkzSkMKr5w9hhW70G71t8nxjp6fZYCv2PIRzKDxPKKA8xIfd71WX9fIznJ
N+kwCUZOmoWeoBDC0T/gvXpGaJmQ3e8uaHV66q+9lYtj9k8U/xqb4cUWWqlbFW0EgtkxlmWg89X0
AQCwCeGXb1/6MyDeHzd/PZc/aZllKljVyw5ChI3gWMT+Nop1X9CN2Bax4X+1B5YS/rjDU6hWloOp
RFkumYlLb9Tjqmix3ejwM9tVDMwolCQYivdYMyEGqk7aWR7adf5Sl1NBbGcVbgs1mgCGcFgNHkFh
iGctsXDg+PYPR88FQXOkwAtqrUNZ7ATQVkDiKgRDbxzs3Ef5Bs/9HIazk+d0f4i+IqcQ9Pw1OdS2
cwPdcQ4hy+mKSEWhWntMMFVwBtbxRm4YVIIdUuh/lVjbxNmZCvC5eiQ/fH8jKnfCZm7PBWK1dT82
p+t7hgx8CcR0I7/krTp9aSPLxY8s4gB6WU13EEryPvdVDtyvhSUUFdJu0ZFs54ZjcuNgmdGKGp5x
3ak587Sjrt5vMv7+f0zjiD9ITHYLk6l6kbM1VG3oM8s8Wof/N3Nqwku0iQX9yyviPou4Y3uPERAq
R/gOng2GzXAJjK60oQCtIHuL+QkQ05BEryPkXv2mHdLtJl7WhP6DErTRmPjGP1jBYvFDQVGMdycp
jCeUuLIYGt+RquC8ubEDiagiBoggON2pZ9SvIW0D87OwD8bauHlI1UVcBpmHR960ZCrig+fQEc/0
KmaJ7ha6KRQMdkj8SqH17FcChaY78RK7KiX4xut7SHEvRiVEtRU9eYYS5GJsCkfrVOyPuHp5NPk9
QiSy5bTk4mvJRzhgLoh3hwSGEfatjZISpWwlggPewylZg3lIhKMXi6CrPTeRTXbQ5yUwxaSkYknR
NmUAzDv14iCoqr55CdlWygWV5ysevXteOBQ2lhS1CfIM0rBUB7TH4sxw/9pQxIIMvCqylJYdkbbj
gg+2w6rDkiT85CG8S0OSTYZc+xdVY9TLwYjtwVkP9OIY2VbeRsKI7PJfUGOLsLdMC2L3sBIIMggk
Nympp8HM0T8DDKToOFNPMJXHGgnZrioKcvuo6HLameppAyxjDBOgvtIgYypQJcLTYebmV3Dh1BgI
q//29QMfebRMMF6GSu1S6rPRN5eKua1b5PojuIAdTEcOIc/K2odf1eSTZ9MkSfcO8dR6SWoTAR+D
tE45rHUmyyrtx5oVlzEVM30sp0GaQ+RRAaBI+pum9tAJ5zeMMyumT5aAeyKX4PJ5GdFPraztHyfT
AeIrqBRlqqacCJFv8MJcqN874jaerDlN7uIxWOgXb0Ia8VWTzL/LlbtFZcyWDtlQf53PPIKuZMBx
CsWWjKIJFz5WByvP1dyyf07dM1PVIRtYx8HAB8rCipS4D6Bi4VaY/UO2zfyKIQKaAewXWzFCI/62
umsqJPTxAnTfyFxd+6AGWu3tIvCxvdjmfxXiasNH8CWTTCgL5RXxWsNK9ZhlcwnSnQHbCpGvTIE7
mw4PU6yKwDZadtnCAfa0StM6xYh0SX8LiXq8wiBG02kYsKWQDpg4e9cADAL+gYwCNo/JB688x7oN
oXiSizGFpIt9KbVJtk0sRjwfwqxch8Qg6UYDuz1ueQ+VKTUO7xFwsMS52bu7b4IhquCIu/YqtyQO
iZxYFHdHem1wTOc+urQF4yfWylxYMG7qQl2k0oJdzwGcFXrj1JZdVqozp3eLN+LQ1WaIEyGM9oeV
PbR+XrGmMhNn5VfPqR+pUkMOlY2+3cGWOCHBkxdjwIupOG3vfG4gQBmFv16ciBi8dbfI8t8FRfgZ
zrcL1h/NqM7qlxEX0LMheFX6+1uBUC/HzLbcbbGfG4NNTrHZI+8F3uOHVJzbOgiY8xAO/rcCTuAV
xhVQ5R7hYPKOdNGoQIMWsYOt+MlwUzRm6LFkH5xtUDSSGuOuxP1Qe008seQfzqRm/XwQHKR+9cp4
0zejBu9SNfcfvDIaamesWz80TqLg+naPSIDB5+qoXzwKAeGhO8TLE7FUZ/dRYYjS6/VsXwInRPD7
TaDt+m3BvtrKa8HLTYHRepOSEsH9b4PQC1250YbFCNad3DDNSm+nce7HxlBtN41hKsWi3V6Av7wC
nAbs0h8TiSaEXCjtfppM/J5w1l1MTN7PeXwcBnlTRHYZlMCEYSuJKlWTJ77Ni95jYSrYyeXsRVGF
XOub3eMxvgGeXgCcZ5+xm3AhKHN/AJCd/V0CZnPxWtZ1zKUsbyUoMbJRM35Ri/tCQB2FkVcJzXTQ
6yT6xcMe08NNvSNOfKaAbjNvfwzbb/fJ5sUkjiQbLzQyRRiYFPpG3v5TJeq9BYjYOUxbQrmI28EL
53XXowBbIqBZPNELozCJAkG6PKKQBXCZYakgfaI68W0iDvYRepiO6JRcIwk0F4MiUzed2KiYAtaM
rZiq5vdXWY+yFiomnLHhIQKtrgJ7A7yNZJqkuxlekiJLBX1gksj7c1TQgKvW7NcJyMFpfT1eZ2Z5
6fBFH5Qd4pEfBZM/UhxMIGPqS4X8yz5nQ0Yb9o22CNpv+ZGEmBzq3rnq0TKNiTb551TZh8Sycq2s
+AFEpWHTHqWQG1RtSEs/XVPvmlTF/0TBxr5pQQ7r2DgJkOU/S4LA2MsBAC24TUPrzTiTyqHdUjED
BhJikTWHAE1eWSt5zIMGIH2Cghun4JVK1J4919BqyMAsg3BcBJZVB24NTU4z2BUve3jyCrMqYr6Y
Jf1ATD9ujF7NMbVBue3fK2IWIB70AuZuKzAudHCcm0PkGxOkG6NF0BJyKXiCorbz6gzaBDnlDvD8
PzIvWtk0yqRAjrj7B62C+7Oytigtt4vVtRSbTfxQmogw5XgNt+5KHs6wQGuYiAarI69+2HytfmV2
Nb99cW0XRSsXafrwX58OOQCKFf7lfkm+V29mOMsVzrDq//qOPfNc5G1rTk6FmP3Y9Ww/XgnSdDEQ
ri+PN3ZKC1BVb0OlpvJU64wfzoRVOFIejidSz5rVsuONZy4jT58je6CMvrCVBWt6zYy5O9dVIwHn
W0Fs0UyZ0D+at1y7jlo0KhVx/gXufg5mA3OUbSMpw7S1PoOPbekVU1Cr4m/QT1E8K3rSKl1XkMJw
g64djNQx2eVtopaf9M0AzvsdDwK6cgDBgjxGGCSjCkkuWn3G4z4B56dAR+HpExKxRxve1cfJuHej
JnDMg3mW5zY0ih6BYdEwHngX5jBMLwTkK5Nfh2D3/qV3nJ0EFhulYHBBPsRf1WlDV8CxCtWp127P
haZ+XHJqAye8qYKl8y1wfasMJPR0LNy6eKClbQQ152ocvmG/SxClpkrJIHxCZWBDwN7Tqtra+Co4
J7xndv4LgYuBkKjOXMoxWm6svF9ytQ3yfdZJ/IGMhanALRbronFVYK1RQb8aE+Mf906o2zmrFbI1
170mJdUw//EDEeecTyR6bf+ymCYsCrL+ovBtXoFzRImuXxp30MY9omBp2OK8nCR/bTUX1LgTD2TX
8TOFIUfVhAqiN4UJiQ84vYTJIhAttEgemnRL8XdEfYolE2U4OR1TXlwF+2VzLkU4lU726leEmfmh
HIiIrbcyXig/RcwwLlBc2kK5i7Kxl/Au4VuOHNAEB1aaPycFS1q0g7L+cXL7YfJ9tBvIIlVfEWik
aP8PlKkPcLFvaAO6pn0B8SAgL7VuC5+y3PwVsb7q8PXKH7XlGhZ8YIEPrJGvvfAvcZkkuJQBkJzN
3Tv77LfLJs33U+a7x+mfv3R5n+53gf6ojxnjH/rZKa74uvakXKhcfPIKZRejKXvmurMDASsZTsMf
kAuLor3M/DWijk5qywdqZa4ms/HnTyRUXjfpGRNwWP4mkDy01BgTriu2AiaXl7A+u+I9ZJjxmpyo
MpS9Wy0Pde9YwS5h5L5JIKYgNEwwNG1Tmzs9+DVfwaN8E6i++Be/+qER7E6yoBYD6LrGmgDdKrjo
ZbeM5cL5ZJHZPNkMFd0AXjPpvPXLd2WRrGcSDAUU0Jbuc0LgPkHm5ErNxjgs10RzgRRyfMHS/his
AqvdYAO440aicVBGK2QvVlsb0H7eeYK4Rm1M8KGv0NVeHV/83CCDwH3lUl/TzRczlRy/kCzkDyFM
9ScE3Aoza3m8I1x/dsZGyCLCYENGRFhUHrw3mpm2Hq4UlY7nEUDiaTRFKjN1lTAGIuPYOSVMQW+g
RBpqRJ5BpcPfrbX+htzsrCS/6uyGhcFaeiRgSuwhokh6tLyYSgcwtIkQsQPCmMZZP2Id4GIK5s8G
sqca2kOt0Tm8FQpLyRGvwJ8gqtH0cixe6M8hidLZQGXtjlSdkY9dU+MiWGFAvnhIX9vOloHCe+Oi
h39UTBxJ8qLayvoRDbpqQaKIPf959yj52odjvREXy7Obzlv6p3uOsysxNmthZ2r5d5u+4ckDqvx7
3TilrSg35kXEj2fXkhAaduNaQuqLB/f1192hg9zCezk1dr5JhnKp1VTIuT/jRg5hstb2+dJ6ELyX
z85YV/XNrMy09qkV0T4tbX7gIOA/XYYy5cJ4s0D6HHhNeijD3PvaEcLGj11VsPyXtGUux6p5XjJB
K4+trt7BwnP1izoauwpuGF+Cg8KinPHNY7Jr3ctijmBVWrno1WNGlUlfAGyhgVetM4xXGapmX53d
dDy7KEcp1cGwSq7QMFWVyTLsY0WEC/G+9uFKE7JOg7FfpF6gmYM0DHi+8tTLseRPKMRLy52Zy9yO
LqEziBGazmQuthYFu8pYDhgNeRkttpcJfOJw9N9+hXdQwikgF1TwveC+K64koTipy/goUseXj9Tb
c9CXfEGXVSA0nUAsruzRxCoDZESUNsjX/i4t1G8ha1/8KYnMVRRb9laUFmlsH89Am2+EB8HSrEkA
WH/G/QUGo9tDFUG2nc5A9esBnfoCscDKditugve4Mqk40cBO8e2ooKwtVVB1M6OouJugdx45hpYo
Jk8I1QJszxTuN1jDU1kz1yehoDJhZDVE8VU9DXhSQNTIcg4mzTR9lpoazj1EoGPOFQ4kJW++aDzA
r1jpjtzrV3qYVr2oGoc/led59g3Di76m4DlV475CEFidtbH34iwIibD7Sh/Upr7MPBFQRxL0OQEE
PYdsjKgqAnnLwYNttO/JZ08X0p93kHbcuoZxj7xplM9Zzagrs4KNLADvLZdt+CPf5proh99ztNl8
av8YngBnS82c2EDDuE0BNa8ZI1MqTvIRePaVp2gaej4oOGZTY5J2G/buQTk5T35kJbRDREYB0cQT
ZeuPJ4lx7wxm7iT5VKXK+liKF156U8sH/i2JK+eXtOyaF73OdaRQWkQVhpqroUznxIcddlbNdy+/
GGiQtRbi0E+UQeOwZvTHoc8i2Tbbtt6dpUYMC6ldE25owSTEr9QlM0vJkQ7XfZRW2M8A6kFf5nzw
hx140edsI9rrWicJcvlr603Eyp1EOslmTaUA/iXa795lUReFNND7knGUkpoU1xiRHop7P2QVQpn2
COIaeYiEW703iqEOqmlL4psTQAEw0OG0t0mOvYf6G0wpy/ULoXLsNa3Cl7GdGzhh8yTsExWs4AJt
znN8GDQoMx9h5GTKqiRH6L8ubn8mchRejDzYfFgf3ETKvqGa6R969SYm+oSw+IIqfOIGUa0N05Af
nQFljiL5lwopw896ogBeeQgnOqmQM2V0mZdUnZvyDo7AqQtHK9Il3QRS4znoYxUCK+dZQAsOYwIn
Tg6sGJQBjiH32PPD9KXHcmIeXoKnG6SiNXJ/BQn4yz0irjdSoBHAV0Ar+5/HKf+w1MUM3BmmXkpH
aojbYxPDLAVP8U0n8AbqKBJySGxuJh6cK+oXZNP322UiJP3d9AcXmYaIqHyaJZJvm7WpD0fOkFA5
9N/PXcqC8o+Z9+AqQYJI3p5b4M6cucE56lN8/UAitwRdj4k3JGSADQpt9jluX/+dBTpiZDvGp0Sc
mfftD0rB+O1GapZC7YXntlzBosgMb0c7ErpnYqRgVxozDl1aDqj9HjpLSN3vj+sgskMrdlQxVv+L
NxHnAKhUQgh6rCecD5cphmjTBUJRHJXdwk3LarAsK7Az5WVyqfVr6Fn+f1L9R5Z4T7pojRXbmS9m
DV3cMtaTWPR7Hop1pdpuvszjUZh6ssQ61DBAymblle3rUu4pMOw2L+HKgn5y/RIpVsRneTytbfyq
/sPcUTSSXlUMZ06Cpo4+Meb9horzKwem2oCq+pT2t7vs49kuacrNBl12m1+/beETktIT+VNfsQuc
jOgyr0/DurEfw/BpLHL/R0c0rHY3eIINqUsl7H4VSjfUdDeQwoECNVbDopCq3K1M5c48iO0ZuhGY
srYL1+/xiV1SkmbzLrMVKkM2tnPOy6/wKrsvsWXJmX1y1517EFP02Z2fCpVXdD39l49pT8uG2FN1
BPZWjd6wo3v6g0StJO59bIlsCC+LfmH4OZ4j5DOnbpw8bRWKESx3+DxMEjo/Q1mWLdQWEsiy6ere
ZCqCovAECulTClKib0Ay49mxPUTVlgP/yDKHUb9GrDD8kY0WuJk1ivFGCKHKCiGqu0s9CywuMg2a
hp5hmjlHbiVl+FRhbqNX/rhHgVKFOiJO3QXrhre0M9iWtR5vNKS13xzf5nAYa24vsViT+ReclIRD
BD1qiwaF2JHlzL+li4pQvgIdrZTGMNgucfIVNLD4n8ORbxuXSpcGxLWZJiE21ME8F8Z4hkFedRVc
/mzM4w7U5YaXZY0upTOjr1SYo9V+GO79RBL4Q5HhFMkdNrnqQR/YcBuicRt6TIqrxuhaphOaYFoz
t5vPMdld/mFbQrz+fsiwWUwZ+a3UUC3bGy2LFuKJrDBit2tglOLG8BikTtw8kGurj558+4mqJRis
oqgQ7fDx1AjHNFvzDvW5hFB8ulipS0hgKLb7keBs3wOi2ni9K35dryosO9qBSQVSOV/YHhls8J4P
bNdu9TApu3Kw5J401uxJ/rCRQwvzV4WkWAH65Fwcsi904KnhSwKrlGHvLDSV0SXlBc1lzxuhnA/8
dX1J9VYA3YqD14Bl1kEoEUCDyrMLBlc9tdrcJOLZySeh7NOhJxmWipivSypdCAqmxDLCqVmPY7qC
PP5CqN3Im4Mm7bSYzOhbI5ouJatJ/HR+myA2M/OLSBC4K9mvY//Luq+Bk6lwyAVjzrJNkGO2wJ1q
BTal/zc/V1QNvwEz4rNFRzqApv5C8WywNDLybF18Ffme/1nOUNtp5LcwBLH+Y9VwYOFbxPk+dn6+
9MYgTSoSViRN0s5n4m/ifUqRQXdybptcpovoaeuD4bE+UKsPDji6qZgjSj2fiAWhGOQeB/Yt/mDv
4oa9wjWi8uM78WbLne+lnTSdbV+e3DUM15JBWPr0wTjAWcVz+Zr0KO5opsb9svBJiUxIKf6t6DxF
0x/i/E/fayxKOYieUhhpjgEMVvwvqIGioCKHl0KcB7xMyIswMDiFAyTiJs26c3kSSbekFYESgMzE
s4tJS2sHCDjJ/QF/U0xBD9lmpsFEoAOVcc3qHBwDVOZZZoC2VGFP4GQKUWz06hR6getin8Kt4bu2
L044+bP4vV2Oz55pqHfQus96GabNN8rAkTL5KRlT8HXaHpph0qfIOA54mdNux6enZJVIKJYXiOpW
eTmdTRVL6trm3xPUdSjIqtrYfdOTRdWOP2ZvJDqtfdbzHbGLTX7wFtPbLnq6zTF8boZdJFJrSMQF
hc+uGQWDuexfYAE0zarMt88GZENZK1FJLCgE3gWfSRG3ziWMKqpwqPeXT6f9tbNXNn6XFv9m2cqi
QoCz9ClKJZwi38puOV3PQPAyeukgOMtZf4nhTxJT+ffUZo5Z1wCmhG8t2T7GqypI/aCFYG5xdiKm
SKrcPcIm2xWqj68h2wrltaKW5X/p+jwWX9sVvxrIj9ehFE60n1T9J2Pl8df5X30zxV8coQGGzXEh
IMJyvSku4fhLTsShcvbQLkrGQIvz7BAztINXmdMeDTbkODUzZvvfhggETHNGd7qAZH+CtyGCgd9b
L1QwupATX+ByWcxW7jUd22zQ6mznd8v83X7Y7YQ0yrAtABXB0F9QBRHLBFPvIVT3zXKnMFbGx20o
bSZuqp82sZ/Rk2wAkYZHPprx+hzs4wQ/9Q5JqzxAGKTXLNKCV6Ds+LLixvkWPSNHNJXlFKd/mFOA
lZg7S6VHd8aiLWYuYH3DmnQJPUyBNSeR3HKY7M390DqJhgY0GyMOO94USeksrUdX2E3E0eWSu+1X
T/vPpsrml+9EsCP/msLvE7tW/HdBblBLsZ6L82QKeBaWiyoFAFTmWMJiFCdRL6TlEWuLDGfK8PeA
Va/T3vRtw81uKApl3rz5Hroe7aLhmSawWnGZyjgiz+oMr2cCoA+pr+AdAEouPnjC/gyp0DYAcgKA
YeXA1D3MMFn/hJFiw3Q1ZryWYq8KJBSbVPavr6fPmv11v6L05DrRmR7l32hh84fmFS2josGyv9r9
4I7DQFpxYsVgLY6V8mHuxZLO0XGOoRaKfhUB80nVGIGCzqGRD1yjI9jUuJddJz7VUCcKHmiYaZKA
QsJfwn3wdATacYWc3r4u/hlSjzGeGJRFVIHZpm54T5NapztY6u/rtRal+1csVuxYXzPu285JOobC
HwSTm/2Fn6xVo4cnD5iCPR/s3Mnbgdvv+8S0Bt+MD723tuzK8Rt5tGn0tdVQ5oOfr0oolEI5wO0H
eOknyZfqwanjhfWGMJ+Ufp1t8KeE3+oxe7pRfQ9B42Z/714Yz2O0P2fn3pSjlCk4wSDntceON06y
FE8PjhjpP+n/WIoNVv1G8/nomeUGxQpnPW54RVY8y43aBuzagV8yxTTRAdhzZXgTKTp5VIok5d21
5UyxlCCYPGe89nOIzAH12J4WrWzJcLewh/vDW1ApKamvHQYOzWytky5pIi52JVcQyBC848gwwGeJ
Y+lm0P3wo6t2H9oqzQLGKDZztirj7OyGgsiR5XHrIaWDRPL9O9fDu1YPByT/hE6SXu+B9c67ZUhK
xz46YMZRIEB5uRWCgWQ3OQckuy/qrKWLXr8R/Ow/8RhxALm/rqVfLaHeTAqOB8jYVfzfQIFcAHTn
NkQd20bIAkQ8NVO4Q1SxgzKL3+B9vwDGCoBZCCn5R/08keGWTP5ZJFFC6Xprx8tVfK2RAzkUKe44
P4CG6RqBIPg98MYmuCJEASzdeEq64stzNGcexwrYslWcZowD0iaczgffnhW5LAo4euXJKHdIEEEC
xjq1O/OjvSRjuMxUjiYsjWwkY32fybWee514isorcTEGWfXIqzesFnvv//ztdspCTwkj5WNDR6gO
bYdbcBvdL884stI49N226SrEaSGTXARhhTUr4OKBb3o9Kimp9yV7x8sTy+3f63DVFsZJkFaEqFvn
iM1l5YryUOSWLWk82Zv7C4CrzRC0Lr7MpG7pBweuENk/J07nFQa2NI3HndRdYcGbP0iPBgTxxFWt
8PQrk9RdqQOk+hjYwsms5DZBK8F65W66TDMhSZRrw6NjEIs0hpG9TDaD40fsuJeh2+6MSX1Fd0mE
clz1wKEtOqrqJkdKMBoyR+oRabxj3Ns/9vo/mVMcQI/S5qtKZ9vC/sDj3rQ1R44F7xuMFZS/4WRA
+l0Sq+Y/b3NaVOonkXEu2M1KYWGnPw+83mlAxRvtOm6/1lRzfQ5B05afluUvIr5+V3Il1MW+Cvd6
zMX0LlzYFHZxU6iq82dCnnPfnFE7ufAff9TeRel1P7HvDQtMKJ+ZK/TCou583ZQv5+ZUoQf+GQBx
+pxiJ+JyUq10a1eM9Rv87PaDT4LNbZH+3P3atwx9WZGBIF5kmb48+81+hNX0tb5pOeD74lSGzcV7
u4PiJn3uDlWj0eFoRf0c8IpE4xmyA4nWQ/JgwicWGuJsnt0Vk7klLXwUnjdyaQdrpfpIN463/xBW
bQd2SP9Pc0MB/elBKd/QjOjQ1/R8+Jx9XxFFf0jeg7nno6ewze0od1VtlC0obe8Wq5A/XGfsNBIN
S4m9kCaWYmRGa3xPdZjrCvd3u53ebhEsaAs7idXV9ukz8llF+sDzI6Jzwowe7t4JlgHKno4YLPQ+
DN1fqbZ143c0HiHv3oAqbSvi7y4xLcxEDGEw7HW9LsJFMJN8yTeZZQP+Q7GgISyZghWukxC1ZmOf
Rxk5udLX66Jq57k/ww+q6enUqx12ZODRnFHsV8M7pz8h00swd4Ac0FnlgnjayHDIDf5Q00uT4m1T
vHwcPT7BNZzRYhK8mvpf/R+0qKMLpTU9ScQ2vN3n06MCUFTjRrTowRWsQsTk35C9fAya/xAB4GSD
YKnztQ/wFiP77uFB4sQMKiZbhsva26A/bOnZwPmXNblDQh4PCuqmZ4q8JRPmJ9OUzIREc4MnHLyQ
sBNS5RLGMs1+BHyeaN3BPpS3Bdb1oqHJffgpuPf0u/gpVnVsA9zNOU1tKH0zDbr9Y6YKj7kOrX0e
ZveZYsLE/Gd7Gr0LKzif2Yh3D8WkeJUkgM87i+DAGhGlOxLYga4JpwscF8qO0ERlsR72uPUV7IOz
dCF6PqfUtQNhjqvTqOi5A2z3GCsteExs+7ODj4XFSWC4RwuHWB0w6iO5nKaZ98qM3G/8CUPMffaJ
Q+NqSEgpzgYrd7H00RzZQBw9PIG88eDA7duaYXPokWImNTqRlhI8jaunnDmiWingsW1M25vCrjIH
V5MRsMJX39rLU8w28dCydPo95dnsFJotm9njJakF4HiJn1Gmrk1j+ikkEiZodVYAKdI7mpThSakW
Fx7UBv2Sm9QZnMswyulZ/OYF65zjDpVpYiJ9ZfpvZNo0xbDkooIOSSkMcCWIQmr/HU9RKFjdPN6f
lUTdEF2yxRuaj74qRzgEToD9E3X4utg56fwi7pNXVE+qgWx4rKi7dyTZ8lhmAmftDP7CajRcBnio
5eRmCk/BqFOqq8o0IAvmJ7waIbiY1cIPCh+lq3rkHQbHJdClJBIs7pcAaP1KEuZyTKr1AHDVfwjp
AvZmeR/LccYlxSZ3jgYavbY+JWDq1CIDOvVvL7hjV8QExwqaC/W0lf+E54Cq8EVNKn16ealHtfDX
yzPSrh5XwoHthw8WilZls1qAps1oUwL7tc9dQkOEZvhuxB/JWft/RN0bJMyOeu4SbsVy9XXH3pYN
PAtJmTM0VzZC1LTa8ghgZVowPpq9M/+Mx7JwD6ytg5WtQkUmVcOoXvE18hSfkLYvB8U8Dfq51Z7q
mSlHVtMJUuVBzplfvyhBoQpypBz2ZXJvTQCc+vh70UOgruV/2aECiFQYF9ZhhEdoPF7Zzf2Q2I6v
nkEqh4or86QfSzT0VQr6cYMU9hiX/TeXq7StggL6rdrpf1XD0rLGvVSAfvSJPRYnKh+29YJ6E8tr
F3tOg4yfQgXZKAg/PStaNet8sGNlSgHn4WLVLaYrTir8Zii7zsQgct8vJkkJ7WMjRGpRucj5E9Kp
/i4FXHMWWn3W4OT+oajPIGc2fhpjxxmIHS8BqE98AAZ1uYu5k+f3qr3u6dPxA1++fQa8gaY7Ho5Q
tX7f4RE0FyWgvcbgw9tKLa1d54xY8IQ8vwgkfjSCvPvnNClnqGMYHMeJk9crXtr6x/yFctcn0OJF
kx+VVWh5ikAVTvpE8T3Y9PiZdCrUi6miLAoD0QklYSZ/OP1eSVH7asZMG56lgp7OOR+nukdb27PM
rFZH7xxWAOIx8mJB43l5vWm0+lXiKC1YBR7tcGbsSjIlc7j8HcLMYAJf04oV4teLXKv9uBClc2bN
6sr5n2d6fb1Dwgiz2ZG2pGjweYG9nNOreX2H7Zc4K2GMPhw4NbH8tX4FFVxNrvCGm7LNdTe6Q9OI
zSo9M+va7KKWj8KuVlICXkUw4sqPr46gbXLK/u6zFvCtPagutYRgMBdg5dy5nTb1aV7HtM5CE7F5
01TwW9bR/ywUQETtK31tqGEdzIuZlT4OWworS8Kr6HtsLH80nPmT0ZIRQCh7dsulzsQDWF0IaFqI
+j90vicww1/A7CQ2YzuoNsHAEkVQaAzcBton3IRLWouDdTpaf7AXvuTZlJSUW7jGX2NB4Qb4zfMw
zP4dWCg6lM9cb1eCx6n7S3CKbtIRLF6cN1m3N58lHWGiRnB70jwMwQ8qwEPD5Nu67mL4VxFvA1og
eXEt6i4H1RDDUHVw4F0IFLyHX4eOF7PwsXMJE+S/IEuBiVatytmDl1282ayRd/c2t6HcjDyk0ShP
RJBJRXqe+lpna4YX0CVHOO8rgkdTS+yA2RRTYvii+IzkOh41E/IQrnws9MiBH9scIOI44vA/OOUB
j7IedKASYYPDNvCqplfFmvuO7AmSBGOcBsRxfXwLkOuCDVd5fYYTW+3A/TNevsOC8SweH314/Hts
zLv7gbZoBRsn2atZEqo0tA23g6A9PUxizmLNL3UGnD7zphB56CpczteKUmqZUaGzmabdmR5a7UAB
eLyEnIrcgj+2JJ9cY0NsBNO3dmQEEJhnTMCbVuRqXNn3D7Sv0WNLQnrWb8RQonLqfvj7HV07aeD0
gms19ZQO77PEAyH+k+vTG0IlVktUGa2YvDfDWbODYMz/Ewjz+di0TZlvZsVz88R0SLwpfX3pfrYo
5FyT597UB/MBiRsizchYQx+m/HD5+WjkMukYuMxAkAZGsKIcETLC+asQcmmB6++mR5AYi+Zde/JO
nXPC9gZSCLYzLXG/YUANdj+2/rY25NUc4xQrTJlxs1lHZDkYRjMDuH+hLR7gW/BJzKLveSB9Tsqy
GwbohosfW+7416S3Wvs/R4xP0aJs3Tfd86yOn39yWUzLhaNM0I+XnWtfOVrcPXN0D6enoEVqgoEz
oET+7Mr3Cb0WV3suF6lOEXd9KejSi+QBheAHkdRmv29os4kfgBePoNwCdEysHTCnLsNCUglN0waZ
OC01R5uTZ6GfeifgZ8njQuJ022fgNUIlgogPz1sc+774R5OAxDeAvZKKOfTrUgsQGGARUIX/m2GG
2ISbPwZxITDqtJz9MnFj4hGO3RehgBLTvCLgJFBDQPLb9bjqxKFACyINH2R+66yRRy8J7v0+T9fJ
AmEdSLT/9CVJvth4lZiVe6+yVtoEdBXj/BK0FyO2BE1CekYD0gbaK6SEVLUBXm69G7wbImkA/xWX
F6d4+KRhqt3GBuuCERYUsXrWycjQ7YmO6QBII14UE93kwnuBv6fLLC7dLOVdVNKyyRtcZX1kUGQ4
nF9XEtmsXUzdpNbDoBisivQbn9ZRiZiLxMQdPTLoCEeL1itHpmLLKAgcLfQgZlhOEFzfqwD0rSwd
uq5r5v7SGFIImfoN6mQ2ms/V/Sy/Ub9xCCEC+uItS582ca9L3xs3McoLpjDeKdtm7yuzeZzIhyNj
2fYlZDTlwhPtZiFIW50Bw6fVyhwchDeaUni8d9938iYQrHekNOPXaQKYJ23N2jnFVUXA5gGdblGi
cczRTTl12d4OlSB95R0vIP6xy4qW1uPGFd6YXU9+xQPcGrOqKRWLSkG7S8hi6gx7SioVOh78uzZh
Q+hxiSV9RGMjvtHawO7n34JRL7XCGmSvjZKjmXSA//tiTbr7NRZE2JBxLbuFc4kCGdceHO8i0lyq
75hI3iuIEwrq4vdm1RSnt21TO2mB3TQLOQvWep39tIK4KxtRdNpBd/fwqz4LIHjI3/Q6iIR2wups
ad816SVjOGRY7p3NHdYDzvom4w8VM1TzAypXJNBJimU4587IDFZU4ry9Jq/TKytcn6SuM6e6ZwED
jpkieJzzz/MYyk9ehsol9sfbIlUAIeZFqKTB0JMquQh0005uDok7W7/oWZvT3zyfQPalBI9WTRPT
9SN41yQ5H0lzcYlTIz63wLsX/lWCYQ9xS1ewsOXWjjxd98awH7hZmi3dFcl9KJvFUyyzxJPQUmI/
3gmLn8/fTLgT++kQs7ItLZA5rOe0GpyNHhKQCwi9VGeCGpK5WA5a2UgE82+Xd880y6onyjlL5A7T
Y/eGeCBtmrVOfkDs6n75IFnulOeepIGLu35UhZeUgFoM1ov6349VR1tj/yfDh+9HXIE22oxBgGjT
d3Lx/ueMyxjtAHkyvIYwf5RBrlh27txTecaAPVabG9ZahGf5B+DqCoVUQ9E1KCe4Zesjh+B4ul/f
AMKWGXRLkOmk8Ostp9dEv1mjRtvO0af7JjzWDSBrJXzz1HkLqsFZijqatSc142IYl7FBXU1QEtt8
3nj/hlc9SXTNs0awj1kLx6PIqbTkU7GjroQE0NeBI2KiviTtxwvUwS+X7H6VtuVJe2mq42+Pt+Yx
+jU/7HrKSZoU1GbF/iC5aIKcygobkDD48c3/ZPX4kQzAiK8kkjaAB7CEPykNwl4kQ96nkw0pYgt4
WpDlVNyXkDkXw7Tx9Y2Is+bpvphZjZZ3myO5CY8hExk8WEdOF8qTwZ9dUp/FnZKrN48wV5kSeczN
ruJPy5oHkk3LN7xWEXLa5y+ds/U06atWXhFgWGpf4eMTP1yVXqO+MsopF2xGYvgzJZjfWUS/Hwrg
sB/xTE9E5HULbhMKyH1fM5ELc6B5OnVXElaPGcWlOb2FEtYDFHfYTdbiZRM/iaO+re281WZWhQmT
OK9ZCHKNc20VyJtv79uWBtSLZ0gcLM5nMOM/sKo138SEZb6P7g8epH6bb9WgVDgxK4442SOmpY/h
QTVIlvUZqrHbggLSYflCypmxIM5jssZC7bVvjzPpGF+72GPQ37Jf118gY2jGLLD9Y9RAgN/BJo2D
JG2eHyLDhtPuL/6VN8z/eDV2bHVidkA+pD+f8zXiN4av/JEq1j2bL5mlhsBiXkEI3Qy+iDu60sfp
bslj2CRh9pRc2Sl4v2I76ZOlbngScNTotqe3XwHXmzspgajjkCOUltGJSyAYIAxJ9W4SFIDNMaEU
7ooX3bUIQYs2ZmWrdxFlRUr2V+zcMdIZkz+c8a7swrgqP0prwHrTdn69YRsFzXCntMoHTEJvJDWj
CajsBk9DfN8KHBDM7aPBSgX/EbLHrjCIZn1/wEHl/wBeS0BPIkzXAXoBkHz/xef376EW4/WZFd+l
1SZoaH+dGOfeVWwJILng8tP8Z79L6DqG7qj0xCmjlStr+qCs5klZWeD7ygGod4nWyvZ1FZla8zXm
E//S+N37eTGhpoINvqJa/XkVEijCjnG8BPMcoWjeUxVH/Uy92yMOVGIKH66/pk0N7Fqh8q5gyPld
uvWdStFr4vFuWvyJ2gNskM3uv7hH/CVW10zb+m8+B5cslQyXcQpt4qTEB7o0gn1nBnVjNMZUNkPH
m2oXtjNa0lX28Fc5KFI2fupUaeBzsX7dMlrXW14H09z2JOxmzdjI4kgqErjo4443GzjH8Q5BFlOn
KNMgTsLjmlIr+lwu0yY0aI8bs0/EUTZGEFER2ZXpU4e5t9KPSUUQL+cL/tol+gNX/N8Xswbl825y
7RTaXsz2HM/HtQJ35MlRSJ3U65x2QG0G7ijtWCT9bGNZQ0s4564/01xC0aE3wcxtBqVjQrWBdVOX
NcKYB6yOtrwLDagYmMRF745mLAYlO7eJD6nLJg3G3DYyt9USV6iaFbJyVzw1HyWUH71TIMS6u622
74y+FfmUCug6D72lLGHScJGkHbppCC3IUL3hh+RePOc0YEFLYsKTRsLB+Qt/iZdiOXhi6yKiT5zm
zHhKo3va3XVl7EMygTCBmMTGTxSETl+ZYhUmArkIz6dKNchBoJ+KeNpfA2OuZytw3OqDhLG0ZPQ9
ISzQgVx60k98kf+LqoE+1j909SIfNqTu8KLcddMXp7iNSk72HXAyN5c4agSX7+cf8unc3G8hx+He
dtrPnMdVdytSfaRkGnOf7x8GCypbHLj6YQH7mHh568TUpKE+TegU+lSqPftUG79GLqNcDDAETiu0
HG3ohhu6IGEEUQ7wNFtwAo8N4nXuj8ZntRURyi2YTFETcD2AKpzUIxZrE+5tAMhnMBvldf+18DQ2
JO0/VYAs7/yMWsE7SvA62PSiEkEXhMd5z0l4IbYwcLITysMhQ+uTPX2yDFjJBmCD/h17VXTWvp30
2cUQfn1/oOrcosTAog3jJ9Yqcl5dovaXRsMuY8XtbJQZMTdb0yEiK9Nkolfst3IeXbx7OeZZJzxL
AaQtHKHe5XrLh+1pVFA1Gl19IlhnuGWx/bmqO+LW6uhpdGQ+BTWBl7tCo8zGmDlfBnhXy8AfKwM+
MFlf1vxtZa8pTZf2ZihaQHEB9dmQn/cvEg+PGb67BdyJtoxc00fTR9hInJKLniMzRQNwBbKqs5CC
dt53YNrV7FUHPnKdHdqUZvOUxU0R9G5RlgdrXS1oF1Pqpr6higFPTjLxZzi85/jUbwD27jb3I2Hq
RJw5V19neU0QCsSZ9DyF5K4rgE9FVXH1OokFBzOmvWWWxPlv+UYHGBCBOdQui6GOHE/obyUyhs1t
JVIifWhGLBTOuoPGWQFAyGjY+eTmeCsETQWU4MqLV92FHD8HCcPvWqyDuybqQxzV1LsE/dyd+BSd
JVJ1SEpcicz56OmcV1qTXT4mgbyoidXj3h42nKWkwqXQN9MmTXW6vxE6KU+nkBSezsNO+xzblnPE
S1C8hZmUYVWGHmRX0y9Ra0jiseZHkGDhjB/X4jiEjUdU6d1St/YBhRjH1UI/VcOINg/WnX8PXj0z
BF5qY2xUvi3kKlOuKpZoRHxBaZ0YN5CXRldS1EUK4E6wi5yB3dr8Bdu2WMFxTwNDFHveJIuGDSj2
jeR29xyEnq5l+WuIR6GmLk7xdlX4DE2tEK+f4+p+f0A8nkmy9ulqiWfIrzxbH4Y+vS7uzQJmqhBh
HakcbVbbPDNePBrIlHboqNVOcunjBXR9b+JiuVQWgFdycoyVQQqNUzCQuQ0Ge/duaUE8mmD2jYJG
NfGS5xfFXCxsXdx9oT++C+OOJNSGgp7g54AlrZFFCUFYKyEG5HckC9SwWFtoQ1PtbCyJ8FhZVudh
++0OMh/Qn7iC9glQ5QfvT0dAzx177xo8EtPOWShhBsifDiltd0CpF7LlrF1DVbPTjxe/NiY6Vfh+
77IXioRDKdHfbF/0IZ9tj4Daxg1fbHrMoCNFo5yZf4L7vbZtxqFxEvwoyjwTVsI+TYWRJUCbmLhh
v/MzJKz+3qnFR75APYsp7zeKzov/RxQC5HIDMVbGvESoNBP0QCx/hmqtdiH90veNsBC32A6r3S8O
J4TNtalYwTU8tKzRUVvdjiHCpte1MXTyrt56G636b3hNXsTk4H6Mf2H1p9xvKLYWJbadZXf1VjAv
rf4RFlHKmQpyFg2ILfex+juwIR9Ii+yTy3CI758LHowk8zVvRoJxmf7WM+w5dR6/CY1hMOB3S/9m
b/FAME9b0O8UkDV+A4RG74spFX5Z8EEYNs8QCOd5eATmmchgWpUPcURSE0vD6opq9n+zRZK/EYQc
1H8jj2zYgW6vd9UBXkJ5o2LRhLxkBudTVFXvbn6IobQlLHCFh7urvQNR/NWFTREoCjMAxbRy6iRN
bTu9xghW4TkUH+u+Ax4y+CIuvKHxVpacyMvO6Eiu1n8zJQTBMbek22V7iDepj0Vp1IVcatU8fSXD
27j9mWROjuY0NlSd3sBdbwqYL0cAeXLdWXeYxczL9M4QSXAANFpp8OcPJ+RuKl5v0AMlbUpdwb88
aFWt2PEZmQ1il4K9Q/q/5nMliZyE9QrJqlw4qi2VH8I8ObiSKqcUzP8DmPZDdVsqajqzC/BkoIUy
IS+EJTlEFpWw5bKUF6PQ9rjmFn0m/8kGKQxzxcjGm49fVX7l/4T82DEWtU8/9pOh4xE7BN/z8l0k
ig+kozhcMo3d8RJAxICai3DpHzwNk6AT+2DAHl4uPnWQvdcYchfjX8aqEl9Y3/WPPHNG/XrLWVgD
tL+ihTqQLvvYL2zUrZ/U+FHxv1uqdnX7nb7Q7rJEo6GhaGDQ2LQXdZbCJyv82UYeSKwW11bVTOjm
m2GeS+C+6unk3hTHQGNjnv7pCSQFsSiy4Z6B38DxF1uRl/qfr78TbP43UbalnTPDobWTRKDfaFwO
dLf2U3o5JdVHM8uvnfO38GMa6Qy5N6Bx3+asUt+fzSUfz9MteW7dwr/ESdzUtrnR+aKQibSMH5gt
m+aGKZuEENzw2plL8jsSlIB2UWEL/ny/NLBNodTRhqdLtpRHMEuNzJDYBS7TXdEQAgOku6b8bE+9
7HpQoN1HFJ8raBG/IOjAEttHQcjChO2WKQW3yewbAtIAzAtGG43yboEgjtBD477OGq8HqgnC6vwz
uia97MUZHwpwO+heZU4BsFd7Qlgkn94Tgw2aD1QKZgyIgWIZWJbWvwny5hj/YNtCfjLglZT0sbFQ
C75DMOmzSq81ivGdFZmdx/Gh+R+Xgv4EN/18j77SU3NLD6jqgzjnjetlNPb9EdtFlVqtW7rUu6Y6
/3unxUC/L0roUfLHnqvO12EfVXjpRNeQJRJqqoFiV1hhO27x+jkDD8ZqjWCev/kzJjLpMh+WHlE1
7FhwFISxmBOuA3UW2O22TCRrW5AfB1XqLdXYQNwdZjRjvH/jLdATflUbQUtLOIhd2ohKsdY+ivLR
go4l4cpZ1dfjcLQakgusYPfU0i9mc1zqAyPED9XIQvAnBJfs1MBTYR0eHnp2sAgOcmca833TAxTA
SMDPjAyC4SUXHvE8SGfiTOJAvr0+0j25vJAo/Tkh2kL2p4daoDuEquoKR3fa61RW5IcXuB6idbkU
9/TAF4e+HswxbDHpiDknsPV1PHTGjYY9UcoZ7lzw3XvZa6MJMxECv4ayNF52ebgy35aApPMGHwiC
7wBMNC7xK47qw55a/St6OfWv5vGftwblx9IXfNwoY/yCW0/mthrrQ7Y2SPPkz14XfcpLAbhwJIiv
j9yn83AU+jPGPqwx5OnflWJLI0yc0e0CoProKhhk6Xa+CuCjWbMO1XT7/W/c5nqtr2EyMvLjqpo8
fwg74mqc/6c6QdyeMHScipfgB2JX3rQ8z3qjwpfqJLDKDdN1Yz8tzBwNHhYAcxMkypL0gDyDrf2I
qEZtDitAXejex0ogPRuSAf5skSuEM3eWX54twETlG4tYsce5Y0+iizEKG1a+I7Dt7oX3E5ZBg/c1
19KiNt2l2V/4dViHf/T0z8dNXSAGzIBWqTl2UZmAQumVEQ12jRMJNDQ7+0cUMsKBRoImhpnsAtEE
Lzk2Vu9SRF18IgR3FkB1ps0B/goCECOx8bJ/9rfyg72vEUXfEEW2F26AO067M8dQXtCVUnILulBT
hgJK0vql1Sy59+cRZnLr3WwYGecvQWVTEGdykmCl5XXAUknQKqaQnTuDGlg/RLcrBv07XwaV818S
75ZO/H8jfjuMjXzUYT3Jf1NKEBHvQmMVA03ntMlNRquetJZRjf0Kqpl84OrV7dyOjIu2172MLoIy
XPurnrBcR1jJK0sBaIE5ZkAzgo1dsC3i9ZdtgWmYJ5NMxZ4EbNY7NgZsuuKN94uEmzE7CaUSejkQ
c2yEgpJgUrRuDfKznUKaqNSGasMgPQh8OAU1aSZ5zSwqeK4IC4Zf/yKwmc4X1FHMVmt13AIUZKj3
cpy2loxBMEFJynnVXDZ3wFW+MpsGdqAcQ7gMgHMqBYCstKAOOhyHXvMvT5fcpxG8qtk60o49DJ+8
VUO3N/QZLChadvTq3K9XMEoHLY/fZcAKuwLAjT82PKiveSbcDyXrusSh6i8xOfZzSNpPjmB32y/s
Okkv2Kv/6QidWaQ5I5rvDH5jznKPPHTJaZV5Rb823+5E1ER4a9jkkNKzaid3KMf8C73UpcXtbrpT
ff2Z3LJC3+1EIgiSoC+nnw7TOFJjH05prhKg+Viuby9QShnR6zcCngJ+MLHI0Cv3xuZQWeqSiqQ+
M9A8POSntPcSB1c4QSKzz+HDQnDGi2nEwtIvjfd1d8BytTp9yIYEcjkYSTggaqgL4aA7ddwpLwXV
SHh7nq8R0RBvK6+7iar0UM6L7F3E9e/20D0FmDGDbfP1LM7CfsrlLu0ldcOeK+XO3Hxo4AddwlMB
yRbpoE+gCORgAJ2yOgYkdojRX6zvH9Ty6nzfrdiMDDSN1KbxoFtj4UKP02A7PDtYQdWe6lb5nnDr
6D7zfVlr+KqITAhkbQFT+AmPTe+85MQTxm/wVOzevUHyeDtRlOZh5UIS1ERqK8BmGFy0WZ5OsQGn
lx5hMkAtFrA+hlyqAM/rCi7yTyfbic9sKvkXsxBrH6bZDDIvl27HusY3/1uoB2gA49GyiOrB5rAP
cif4YGzmlpCKIPmToh2dYpnydW1SP0LNBy4lznBRw/zO9vdAUG7zu5KokI0pThSvEbBvkeBeBVLm
dGmA3TLVOUn/0ENdZA61kiS6T53bLoEj+BSLNmJcOf/sOApeD2eOvI3lVDpN42vtRbPWjyc9H1WH
2sIgHpmWxSpjUAkEqhrQlZzyZcMFqeP+PdHWKBpOVykhIdIHNKR2tzXAUCE2uOM2dg5uxszE/6hf
e8fMl/EhQI+E4hJB4J40hBAYIEtVXNdevCdIvn2n5FDn/Ss3Q24+i6NRs+fpcAoX6iROuTsPItPi
pQzOTmcBectdgAweOOlioADWBMloDzIhJUJkH7w9GLTVopJ2UoH/h9IsNoHk5+z1I51wZbvugxDr
aSl99Lfw6tq34honeEZiNMQXSoX1ii2P9IoFp552u8GjHe0sYB5w10jCLtRAqWm05RRBPjKa+vjY
84Ubwh/lGcPOJJqTMmSR7Wfe+T6SJskpvUGl0JBqh9CLEmhCMHjHh8QNWrxTre+qK2jcvmuehsiI
fLSy4z/1gvy9pchrQTqbXQxCOunuIJVniI4UZxUOzawG0L5hcdGnTlWbqkaLRb9yXYMFzuOepkwE
oXkfdsl8PVRn1GJFCtrV21b9qWgVjyPlzcs5iVJV3pFeVpcFQCP/8MgLH6NKEloY/0IW7wBsLTSr
UN35FO22bCnJKXxCKmcclWMMo60DHYAKE/faUzXZ55bVcsznF5RgEoWw+wbt1gRyvZnk6nDzmBi7
CHLn1nxQJL6FeESt2FQUwlWWOB8dML8cA3JWdau8vQpwbBg9Y/HmzLG1ap5rfpIPdyqhbGCbAQEf
ziaJ3WdYZWN757/JKKhSUfH5bFJTyPlE6t9sADLClCyy5y6TltV/OebKfAC+2/woU2v2+2AWFa6/
l0Z/kMvaVaGUlhtK9tQjnoe4KI1Tz8StZqV0YptlLwKp1yYwzIkdUr6kvjIn5Vu7VtlQizX8y7p4
JThjsFdr0kkP4ieoIK62jZdczdTiDax4pj5GQs6UkOrfNwHh6AgDa35NcT30m/pqcHTP7mD385/z
zSr3ZmLpmhqzcY9BxC4omo09QavXnFGb2hx2RSS8Tto9hI3dAYQKMv/8bUUZ05oa/toKAYPc5qyK
rDmlaf2gkNnp6P79fwKhdsFVRKOyuhILjZPLBxL+iJ1J4rf9EY6J1amfkdtKCLOfBpU5O0o1mISN
TYtUlt+IcrO+NIxbn53OJI6Pt8Xq88Gb0kgrCM+HYr0ro5Mj0MaJKSyz/AtZycZxubHZZ+rcuoDj
7tqaZFO6pGHSQXSRRuv0Mk9ve3JLCDTmBIYSvdDksgncqJT1xbaht+k2K1O3kgB15qnA1u9Qgxmn
7tRsq99OHqlquygnKt2nnT73v8rW1kaMySwTISMAGwf/KcgUIhpqqdK2RRILk1jOOjBKoYH682e/
FWvBHnIpcgeOi0NzEPXeCmXpC3NCJlisRNKZVDOg91zxiAuoT66aoHl7DMVT7YHKVEsczlN8BVUp
1WSBgNXtK8Peu97SDZ07yMxzlv1FosSGfXS0KB5LYDHFbG9ylWLpn57WSIidFyeq0U/cipE7k2yy
sTUb8sa+nN/VZiyr58t3LQj/DuBGjKLO4UipS2k8rAsLadlYY6Q9/ltXKThyuiX7na6N4JkAurhR
1N9MaqAAz3v/gk9kLLQvUwxx5V/Rj0LJ6zWDuA0ugdm+7BkwjIvRLyQPjOMdjQ6zxAvTX5/ZQaUG
GJ7LxIhmAYm+344N+O3Iha3ah/yx2TSPvslbN3oTh7W1WQMqfMIsZuC/810Z8k1AC/eeKSCZtV3P
b2ea2tjDJ1hbG++b31kx8z/tjlcrmc4nUJVMGJnHT2WlSeP51bUcAdKCvkd5yZyiTs6PsXIXioLE
pU3t13tAq29wbEl1nUiLKe+Gtt5X0GSWmKOPJi2+oSq3UZMswA8Ma/zrNO981JUBd5pErVjUn91N
ubUA9u767NeGW1dCpbNph6fsdVLdRnpRl9K57dhMpnmJqx7DIDR9AnycEMKbLMzss0yMYyfX9bhH
kI55KTmYLzBMhSklF7ItkxuucdsInxO75QOuyHXdz35QEchQ83H5FZuF6ig0sx+b+IkZSRe5Io6l
GfyYm/mZNLFfaofHJOaYdGJ+Fv1hZFosKsiQG8+dXGXFZiKZ0AdkUITzoF4Y/E+20HUxI+xffVzA
LYw8LtjPHfSfsoEg7SdAiNXzL/wdV2E8ZIujNFEjo2/d83Eqs9Pr3PFp9+oFIeLt5gQ7W0b3QyD5
BLzZp97nn3CpeoryBGYpdSfzh/DrD+mZdtCeeTGlsMZJ+B1YJnZnDmJHPyFMo1In0IIXeYKBY1bC
lRR0wK0Xdsopa3arGCybukBqxWwM3wiFgYouGw8+URxVzh6WV4ye3DTyTKRpK4ptRhSpYAO40h59
GFXaUVSmZpbWFjS/kw4PIUflCivU438po8SKZ82NnSzvS1mRIvzOZQzbzZ0oQNXVwEGEq0QbjNUi
tnWXPKjfC2kix8upVCQ+3tBm6WQymOTNHj9LUfj+ifzwe5DFALehvcRYsoeo3QZ1/s6ayVmTXVxO
Q8iTST91Qgi8dwPtAwZDIWWpUwgv6+vKUYrVTKPOZ771RA0MzODwYhngngAuAvaPhdQXiF3/cky9
b61EYud3xElWa2reb05gFKRdLa2JqZkpVkVlXmsHMD9Qtr02bum6Wk3gsZa/S/Gt2gQ+LgvtoH6O
6wjGDLMup5O6QD9glMeGSuaLfDM+XqKhnOu9vGM/f6jsGtr5nASSvDBvMuiu0g7KlMllXy2wuART
knyF5x8em+rRaqrYvrmtS+VmWxEKnegqB3MmP1FJDB0obTGswVJHaFA1eaBBgceTxCvNvcmdpmz+
ORgLjL4SFCeNMg6WdQGCfMkFuPHL7AEMLSDVxX8RXf2wyA6+hL8DFsFDfPQ4roLMk1er/MgYmUCi
YnpeSQSK3aw1GqUEs10xNadYdZ71j9Z027TVh0BcYwvd+JroemxRFpGc51Rzm8M51Dd0ovlkj/6W
vKqxfrrAK70qkYZDLubQxQr9JQIcuE+mYeUiaajzdwF6WRDTxpcjBTvKDY1MGTxUNEn1Z1XOpVs5
4paH9HNKDzORzchShT0D+lyalFMbVQhgypVTz8Isyw/YaKiSL6glXhaSqPAimcWmf/mCh6jUSZ21
+79EMrt40JfhOGT7xbGX/Vr1kAgAmuryUoWY5/0M7Q1a9hZ6P9kDJ8eljLneatZd45hwdalZnaT1
I3nqFrVXjeA7gPYWsf0wiHMRicc8QPjVL202EpFOrWROFVk+QX+t/CUPb13x1M5vrziVjGFtBCo3
u1CDfPkAvqRZHvShleUqnr4ZwJZznamHEnmyKAThYmVYHOetx41WIcF6d139zC93KI4maPVYEQew
invYlq/TZ3LmClrzh2D2P+Zk0DHrvbeTNvSb5SdTUnlUrIVk1kHg+sBTo4w+HufryIvdBDnf/cRD
DNA+5aCy81eoLnOOPNWc5jPLahJiEQqRe7b6E1aEn4wN0vSwarjRxormzdg1EjpbXB9tqpIqjqDb
8SKAs2n6JQ2AGs9X3vw+Ufk42YTDCXoH+zVt+7cJ6DJ+PJtCuiDRpd2Xg4leIdu+hfLbQmijaVpx
6kk6klV2yXL0TeK+kJv77Lg18I5n1YVWmFwx2W5WQuiAhNbh18BqmUepbTGZfsAV6koTx/XdfJeK
dcAKd+58w2U8FC7wuhy+ekbOie8i3MtNsPlsgk4KCAcEDtCbHTUBJpbtog1pPksb0+s6P4x2ANa5
g0ovybf1sp7hLelugKe9iryd79jOB0zgFfsNvzpZjV+eveVCOgW3vJPtEsYrCagxbhs0aaoCo8Iv
NSgtbcTTKmmLdDqzLufvcx9vM/RtMbRm2lW3x/x4BKqhL5Hzxsmirh1XC7R6341pDK47sO1BE3/A
DMh1Nm++7jbfx67vYIO27SApWUGu97yrm750VC+BARDI+4slxah96NNTUztWiKF/lAJjz/BR3Msi
ruVgoA4K6ri+ev2riJCrl/mpNzUPurBeruX3jW2kpDhwqR0Z8OaLqc59sfouJxHlgYjJztirecxf
tcnkXw+uQS5/VAw8KQKhZyscjqKC/rcJAbZZS1XY6BZkwEILCRM3CR462XZc9YkE0tTbgz6xFLNR
JvmNv8WOL+5PMc4H3ZX7YGVkx3BTrn+kPmDXQaCyHhYgS4zrJwpNZdHYra7zON7WeXKW1aiia8H2
YKC5pnmbYf0y3nfuNtzgwpM3sXCK+LrbgPHnA/L1CD7Es9I6Cgs+4gbr/74LvXtL/1JxqjVvQtEH
NwUsnCxpV8hE4MYX5IlHClgbDFojLT0FGllJhjLiOjMJm/g8MBAxJl+sInZHxnzMVExcZdV1a0Ww
5LdE6n+QqwsE7q+9i7w3BulevoQElRQP/44hHNLa38/FYHxH6lDLPSALpAOPiULhgsqAY2V7f872
HjXEqLY2Gwn/hcSe3LzgkytbPWD9pjQHbRJchOloiSE4G+Fmtkt9ClhQtHLVI2OfsejbGxbUSxR/
aA1GMAjqgis9NYpO2MHsX2jvFovoXCcPaQ+JhyIV/PgFtMaGX50pFLAdp9OLkqSBsyNU35VEx8as
+u0HBCKNZgS2H6zVfrnB/6EBDaxuqf0N72HuA00HrIMWEh/eVCPAtZJH7xe7SpcvPvPHzAVfbakg
da8li390ct06Pctu+JrSITalD4voubi2yWSaMCRgUJZgZpievMG32eIYgtkIdQHVwPIee3uKk3TG
7Y38cfDlpBi7Acrs4rCdZpcuRm/GOnzjR81N+Dsb7ZcoUv/tkOWT051mWDVK4qDNf1yjWHJT8hLp
Fx6nzwx1VXZrO8w5JyMAI31939bYASt/EWasdyHkLOsrsfPszHO5PC7d89v0BiiccfpBwPR6Kbr6
9avfvg7NPUEYq2l/jWiH/7DK3fb94EDvH/keK5UMUUmIp1h4so2DrPnH3h9XldvLKMqnJFS6aR9V
RInd5hDGk4g1f4bZdny927xAWviC9F9Ofo3kzITD66voEgN58b0UyNiMFpt7ox+RaElRb/XmRFbJ
u4M+AD3O5n5oyzgOhF5TUzNSsQoBQ2WrDG2LwBEl4v2VPq5rtlZA1yM4Wfb7Y5Mbj9+CNnmdm56y
XDLkpWSOhewukD68pvcEHrdwLPbxveSukmFqKelOoLNGJtZYNE5Vd+12pEHgCHU1duINmHVMBr8u
nAYe0zXbhrjgiTQ/fKUQ053R2uvaBBNgu4b54nudPup4A54BPqik6dkpbwzc3QX5MeMf2GHapAYY
JIVwxKqx7DEKEtd9uf9xBF5yKBvS9wgQIFGMvjCbOwdUtinxpitCH+eQcmmRl56qb9nQCYK6mnFr
R5nG/vDjC6TZJlA/Bs4JnHy7gkb8iiGd6HMNGVZTz8cuvjsxyXxiwjbh5yKaBwVIZxV5xFHKC6Zo
b6I8+vEtaxMraREeSwLn+xDMWv7MQuAmr1p+EDT2Cbq6axkRCmm+0L0cCPBLKx1ONe7i60BDEn7q
h1u7A7L2ygZKtYrXSJPP/QOqAd1v6FmD3ZS/5+1PqpLdUdcxmxssWWxM6UMUEs9NQcmYFjCXktTy
9nemZLTBLpVN1yHFu9GnThCa8ZCSiV3pZSlhk1oHVA0aDLR8BvbGDAgqc7pZleletexi77mI0hbq
7mEqEoJOtJ1qtE7SW/r66o9nf1jDRngIO1rlVur8Fd+RaM/qzLVb7X93Qo8n5x9M4RwE8A9GhXLQ
cCvnjn80X+eP5yA1vSlUgtofz5JT5fSKG9F6+bczNCk2XK3qu3yt3D1MU6InFatqPMwnP0iZfUTf
3ZGMtF8NENk+Sxdeg2iEJE4RFjQfS1RNsGaULJmyBNIM8GxQ8ckL9RD/Xe5ZYJmkz88QHRzYkevV
FKR4cqoO2pcdpcB9hqT+VLsOSVx22wcdDa3lIYz27jMxPPvjytwnS8FPBkiU86q0/UvSIeRTPlHc
CBF45nIsuMqf6/XbamT8u1T/3ADK/IrFwx8CgtpE51efoxaqyNkW4hEU8XNzAO/otMmH64M3fZL6
8rIAMChv3RALAkiWa4hYVTPVu6nDspSS2V+pylgkCAxpUkxWCHbwTAfDgEjIDn0alrBKO5QmncRU
MkMCsnkjvX1OFum6XV2nw5ezNY0FfXIctcHvtCQP+IqDHOAip5Xjb7YD8/jXGvT2Bqntj5kYQN1L
BSWOfaVbZVUgVzEO34hD5JpoIAJnFUBPyTrnysgjFKaPyacTxKHRxSPPqWChpQ8i/4mrKB7lYMYQ
ooE7ploWXgD7Ml2I0A3iMHSu24WvPuDwiIrhhQy+2Sqx/GCBSWW/VjQJTTt4uvseIa3PMQe+Jzup
3pVdoPJFMol+YNiHlFEwfthsNK6gh8NtVZYXq75ewWDTMN0DAYVUE8MQyU4Teht/lLxxzYNEVTer
GcTOUFqeHm6LlATBD0DO0m1Zj26fE1Fdk24CwX+2JGM4lpz5DMRbDd2KXZQ8WgHYSU6d0eUBwgIi
Sntv+ORClG5BXhxo/91EJmyzfnDc/SnoHs3oSYq3hRwjZFG6xyHWT8/DM87osVotNXJLk45KN0TI
r8QHAnSgZ5bx8ntPZubkRkSzBwuHbLFNwHmOc8/zldDIXQmqyzV/KqZMt0+1tPWZqJ66LLeqLXMA
27FeLMJmsE5JPauQ3XIGwAVo0/vlasvVfBq/swNrd95LnH8cbi1t+aW/1Dteoaia/ACC04xdDPy5
QIGBrkBO6oR0k0IMh4k88m6Fl6uglWNOIB3c6BmuOGCVWb/r/h6Fk4Ky3tAZRgHdeHGn4aQVyggD
jgu9LY+SP09auKgSkQffdzcmrlKwZhQM+RAEvWj9FYKYwQbeeeyj4ASBaPKMbTwJChciLkit7rNf
y7Z2pSvkuMIi8Lqa+Dn4VZyjBTMpXS20dMl+JOv9I6mFFRZMSQpf4UchfLmqrmdmH+YQC+8+Vp/J
imvRkhWJmG4orYqGvRkUYhiYe4Jvxk+pNAvorf7P6PClYjJbrGOaCTHMaSX4gf15lpd/E/JIn+8u
CuX00QqebHx1pwdb2b1hWLN8j4xR8KF3JjZSP1CNaMad47MDgUBkBIOFiAgi50ulSa7FLj3BeoVj
iukbJ+F3nJAWr3T+MY6a85h6HuZuBeudnLGOxlX21mxSUHR83+SMD7lVLrbGImWZKZv40NnHNXiw
jFakpI1RVBtelDCacOt5G7F90PzZImhuySn7In4QWJLINy8/zUnGQifKFK5v5lb3nNO57hucpgA5
8eQVTxfXx0+uurJMqLVWcxnlnGjAb9mt4z3u6BiVl9xZfXWpDVTdeqXENUbo77MHNx+oE8kDrnTx
fMkN415EmAjWhzUcD9U6yWhkMshrNCepJzbYlZGrIouY7xtxhwL9l5eOZmoFe7bjefnpYyjWvxnd
+4I9jJh0qkg2RomCCnB4BFeokJgJpZ045r6IwOu5RujjdZpX4/38UA3PiQEBa7tecJmXq0rslZaX
izGPUwDhQGWeQr66xC0+kOLI8hqyP3zVHLK5DXoUH0rgMiZ8W4rbSiMuMYk6F2OjzShM7/k+FgDO
Srh8WTvQ7D8nuDty/e7b9t32PNqSmz9f9WYHCIoj5j68wAjSWj8Dya2M6CgNkw2kY1GqPs7bxLnd
GiiJiWVD3NrYjW/GN0w57YD+dNFuXvhO19RiItoGcDB4b8zWTB/w7s/91/9AHwMKV5jPNSl7xTyK
TKJJ2Y3EywdyJC1rrVPO/IqfX2j/MkKRZEWPaNHNIC/tY6Zf00ppILkMn5xKme1Kd7OPNOCGS+r9
wuTY6p2RGgNt1dq9TyMPV2MIoI1APijUIso1FvWgTRIqdKe/07646qxbBilkN6NA4oUqfEwBj9s5
yJQdH9JGYxChdNH4Bcld2TQDLyNRJd5oScNd1nUAWhZDR2wEa5uizb7liVVxHMuDKP4QtkmvSL8E
1/vQ3JqYXB/qZggeKroQp7p6SB+oU5ey6G8U5XhVdTog4Kex8/omhRbr6Op8pCop81wNiP5RmjSY
DhJTs6bJMQHLxpm988CPmsL8PMYic0MHPBA+a86VFGgnsGTAJw0AtS25dZRbaGVQnkG5JTnFt3t1
i1r3f41uNbmrx0F7WPbw24MSass2oD53Czjh5JeRB5h3sIoDtqXI8G1yrDNaE4maqU3NyJDq9I5G
nIDABMmaAY8kMWlKW4YMPkiigD/nwH7LKZcNjuX4dqvCTYt716m+cBxUfNg3P4Mvn6RbaOvYp3Ts
Ikf3hioLXzh6/2+uyiow6RRRJoq4tXQzmBCA/BUIIsmj1mocmlYPBkcOSpFZoQmeAtWSATVjvoOE
E78JcDBtmzndHgE1lRuHDEhjBmn77XF0vJ+CHnKV5rI7eX+WStolL7YkB52NyDFFTQbBQ9o58at5
ZS3cInqldlkqAaPtUbEGHiEy8dmStvIDVHx1CDuseWSksnfvT7Rl9prLWZAJByoozlJ35YDI3f87
ztBuefAOpA9c14CUzHEy1HsQaIHov+s04EscdZEGmJhvSm8xbjMS7WPPioIH9ZzxnOmBODyw9bBI
5zphnZa5sWpjZOxL/dlITfYiU2LTlALt4ti8yEyqOpVgYheXRK1r6ZryvBvystnvn5NMpaG0Wxgf
96gXRCFw4EAU5C+YGtGsKcBfgNtQPCUv5ioq4O4zK/ywO0YldLg5I2jS1MVJcj+3UAiEJ9ge5Joq
Q2MB42KTGOkQF76rHOrda84Mj23pd1V8HFqO/nSyrohtRu79fJFjQcKbi1jygvXW1ndl+xWfRrI4
vHCZTmKISpR7pBtheGK+UzRby8+USzbAZRtE3q7DMbY3l7Giopx5uocM4R5dlDOQp2W/G9wKWdNm
GiXIGJhXO1dCPo7EFUV0uNcBuobOjg3i9uhwjxGXFRZ9Zar6ABFMHysVpWWudyHqGkZAu5S+3evw
dk0a0VBq1lUpj6IPqV8J78TorFjQWVVj0DAHamx9h1v2fB02U/b75IigeQntPFZ7qJw41mqBSnnH
dZJiLLF6+CN2dgGn7/9PhPzQ1sJuxRScERZ7ZAsoOffD0etnQwrVoLVGTpyE7gb9TXD0L8vj3TxK
AQwM/6vWwqF6Z9QKYREYN+ILqPxzCR+LMioYR+x8Wj3JcHCNgc9HNFnUVPcody4uYl4q2hxZLywE
cVImsAi4ufNLc1J0AFaUxpyQJfttl2+fL+F49xIp3ElMyVLl9P5Wh8uLHuiG0YG9IcBu4ZJDhtsw
Oa9i42eo/IDF7EvQwqboKCXSPRwIOg3eRjFH+rGRsC3EQ/oZtA45tyCBiQ2jaXZRgyaUzW7xm+Lp
f3VdwLFH1RaEj2lAbwxM395yu/6AftsY/+huBAY2eSD3UX/+C8RUcrxaxU5HzEwUEwQcB2P97Vd1
hw2+B2YTdJJ68kExQlLxuVak7VkWfJ2gCYAgrVUIt3T90oA5Nhs19PMt+V4dIVa7KnfdbYUpTQqF
wjJ81uW4a2X3L4zFn99rLomzBJlHl/TSlKtP4j4KlFotCbI24VPlZ0Kf1/Qsq1tc6bjB8YqsznJu
x704y2JVQF+VK8Nss3Bkxn0XJsXzf8rEuNnmOEtNhlqzkAIavzsj3n7VMhecHZ6HoLp9909DhN0v
IZPx7pkRy0r/2bRstJbBQiVSvGSgXo0rgD7UpC6aSPQJh+qcghkxNEUpeqCVaE7ZAraru45hmWp3
ZTRugiAUGUQXnn/YGsV5n8RbMR2PWSHlHJEC1LOWOZmo/+DKTYrFWhg10JS/K821aut2OhLcVf54
Sj8mWa05fhjnKkm0d8RsMm3EFDxYtsaLwybIBQUFiwRg0T9simX5R1CYwz6SVAuDYK/eyC8M2+DE
XyTmqyBcsXsO36UPLAnwqDwaUgAIhjn1QXTJZM7CJC4d8elgM6hzPgxC0wN+GpEM24odJJaLCpXz
1onKByVk9TBvgr0rnLqDX/X9H2EVVR/jFc/VohuH0Av7+R4DWaqb9RmCSO0iZIoMRGoJqCsjcqPC
z+5VsarnRPT+Cs4lF9rbmux8TlxUc3ytydo66FerK2zQDS/S4pTXwjTqTVavlNUrMdtvL08aNn4j
HvW7AKJxAVBNXLDLchqhquL07aG2ttlOhauffwrqUNe2brrlvuPp2q8CuGhF9BjPsGgZOKiA1UIc
Ttd9C4DeZdHkq/H+NwmCu/XqQavTOTZbBc/7I4vLN66FVgSCt56JB8QLGTPi/z3hLSXwpY6y2q5u
Q87oqQvZ9VPZMnO7EGOUdALDFIRqJ4hZMoSBAYYeDwn2888FmgUuo2qim3M3PGS3keY1LbEWXfZh
vZ1KxiOhMmZt1ymUaf5vtrj402x4v9lh2Bl+6xnExXNLg9MvrD9lYXgoCKV+oC2WqhCFLUEnu25k
maeZUtzBC14Jl1YTf5eKOkiPsx6Eie1RLxQx1w2ly/18E9jMlGupUrKsLaSGkjexjX9zl9J6sFEQ
BSD2fUrCjzJWaCW2WRl9s75nL/4ZDLPge+zMZwJo+XF4KKJTqnOzt3iSiB0tFGJDHIcXImxDstEw
SGVqhyk6vsYBL3iUxJCD2NapL6tVdssf3A1pkRuTMGIsUtMwp7vsY8Tovc3TKUw50An5ZsYvjU2L
SO3se5BudHY0ar47W4hyHszgE8ZAlaTCJw7KXCRzPk4j+7g/ik1PbO8XfKW/9Mozlkw3gzhGBzgF
sDXFIBzKa0R4ou3EZEHLld8lORAfrQHbB4CiDFg78ekmKlFovVrYwu5HutK//uj28OC5xcS9rMBQ
ZPpj7GoqrclW8xbF1MAV+7iR2m+rBANef2Fnn3I3O3W0R9QE5NmwlqV0B6cku7oH2iLGG+MMlXUF
tp31mrufvhIgu3z+n6Bo+4eqV7XH+QIUomqKW44cb4RakRuae/bzOD4LOBKlksrwTjtCsCxV2Pr4
C5PoplcHePAzOu65WKnNG1bFwqdadtaJayV2e/zDrdh8uVUTFOS8X74jQb+BbrnfFSIs51NikEKr
mVnhricjWtk02a31uVyPBCNn91RISfZELuTyrfNyF03aVCs1P0gl/cXZWh6j2wA5kofIZNDdZ35g
BbPWbPCDTFbkWAX4Mqa9DjsY8kLahMCZ1v60aaDzXJhggy2lERU8N53ihfde/x9JGMET42CIe0gx
W5yNpW4YObfr1b10DUCPfyaNJNKXUOOn5ow/omZ8Ua+/T6xd5d3tqARuGSZEYdtaIfFzKwFjJc5F
gBIWnbTyjF35ZLAVkic/ADwjf0mZ5sNCkqbdxZ/MHHIm2TrQP6t5+DUYJ46GrIE+Oo6Z+UmmkrD3
jO2MZ/JUWdQMmlBFG31u+/fUZ2uLvz4hZIe/6xO6VafoWMNl8LmnJfkF9pAU0AFOhvJC1mPQk6Vw
oZZVJbggnsUPv9uhXWVYlbq0H7pX0FWtthG8Z2TBYEaBj3LA3HDycrCRyZjLEIydS2X7ylqziY9n
ScjVLqHeL00WalDDpztJC2o96DdONAWvwfdINpPXJIFtLBKs35Q/31SvEQVfly1zgPs/76DBPQE8
AV+D60Vtm9HvLP+9j7sz+7RcOYHhknbhxgxWnhrBT1ZjQ2sCKRCT+utlfin36yOTZA17aKnmiFzv
Utucmfw5/x316N+L+EtXB6+QK3zFS4TTXBObjWHptc8fGHkSKFS4MI5icFxz76pGpEmaYJfrFcuf
XRmFUM+qJbCsTNWhZ+pd4X0INTv0CeX4f9aQhG88B5sUTo0lSirel5hGfkdYmyFLZUrI3MKu+eVw
ls4FTqQkos22fpoLrpj8llU22mnqu4NYROBIsyGLCgh+GxvpMQE0FEaSblKt6mrq0RYYNNSVhkld
CrnqYsaY/UpaGBul6kV6L8Z+2vIN04ZW7IrSUJz4awVcw5joyVXcgTL3VpnOfUby7yv7RjAxvEFt
M0iZnHD1XDEa2hwUEMdc35fEdzOTidYtWi9lQa+iG3Fa4BjApmkhLx/f7k4VYWdCh9DBer6NzQKS
OzsiA2h4I7EAACHXLJOoDnUUk6R30Pnr8O1UldvSmzm6VJqeQIXkWfz5ZEm5Uh02VEHrJofPY9aD
e9jRPi/Nyg/UHBcm9asQaLGt7mBDAQPjIq7teftYCZB66TkV6x0Xgz5Rr87zNZ9XWk3J6dQ2EmDP
7v04YFu5jNu48iIO8Kec1Rp1jPTX6bFbkrTMST+4ZwJ+cE8HAHSyvSwhdfCr6AIDX31A1ZhJ8l7+
2TFrnW6jybRGNzNPY5IiGx7/DhGfEH8vsW2ICTCWU+Xep69TVipx31K4J0Vucj/BrdwJQNXfl6h4
bA7PBLrQZO6HRVygIc2YbOa8wr/JwzBke0ei4L/Ij8Kyfw/vf/XWycxigJlfV51gF0dq4/LirGKm
YbQtf1Lm44fpT2TfxCUKdHUz74Y3j1oA3MgD+xwtRX0okFBZFOypYCazp8jWdbBLWosVsBJovb1W
3aoE0xwOuJ/u+ZGlEwk1lValtmfl13ImgIXGVNMwW+DwMhg6iInvgDoTfT3IzaBBY0UQeqCf/U4F
zbfj8q0rZxe/C0sIpQsG9jTOT/lndAtacpKb49P6cJlSXCxFq5KnK8R40V9gkRGCQ1rVBqlEh03n
REBR/3ldSRyHnE1MxS+124Gp96VJJP58VK55xjzNUe9G6ISs5v0/o5IevIWoBihFDLEWuN37t8XS
+bUjlO9EVtGV1EIrrg5ZZ1Rvitiuydfb0wYCIgTnPWdZ9/uyHrL3WfiI5OfJ+wq658POMNdKfrV0
p17Fk7KqteiLUI7klBFdoTMRyOrxRKjPP6NXkodyl01lG3B3JKkZh1QR02U4LNdPq5IjJlM1ys/L
VBJHsz61VUPdFaMNyZRqcWVeugwG7k5P+Zds/xRVzbp7yDT/FurBPJ/et86Gt1jH7VaMacDPuzex
BQQV57Iaw8TMgUOrTggkB/+7lAcilHwCjmLajQr4pH13/lRPp6G+LmD2xIe9FJG6VBq0WXi3qlLc
/Nwe9BXVXO9+4Hgh3Y3eAmsS0XrHPCiHrUV+2OyFxtsLz+WYrAE4OmLjOysjHuWfy8fwMMjkWLIb
1wNPHxjbnYwMN/o2SzrIOhMTXJMqEVlCqNko6PHbVnBH3y+z1F3Fiff9Si34wjf8e4/HJ3tW9Cho
t41SzogIJ8uQkQbM42DpuJZkPu1x73MZnDYKX0PhEwd59GO4CKIDZGdWTF2lfBm3jubSfTli0tyg
bD0OFmReWHOFZvmWQbb71PTZQCGS8MMFZwMEb3bAJzIiMYKtR5Hf1EtZQuXtbpOMDVAN449QnXn5
69KPOShLRGIOyvUlVjQ0MxHynegIUEfsrG7CBlruIe0amt9Pq4W5LamvvShy1S0EqCC7lbV6mxur
4kdxYg5uyf2e/mZ31hcTlWQZDuxrAT1yitmrx+5SQM7sgiqwJSnB7DCulBBNpPPOivhSuxA25DBJ
Ek229WhPYX+UuNQxeAASMxoauwrBUFi5RA26suBbR1+NwbpBk/MiDqltW2QhBd5XvN8DwUL07JpX
Fz9a/JqUdl/xA7/vINV8hsL95Mhv3rRwYHCbBZ3o3Lyb37BANngyXMIjj2ljz0gaD2HDgHIR73z6
pNgE+qsc9XIJwjjFMGIPJI+vkUum0Qrxtx/nTx/yNfeS4zBr4orcQ3vvnCytezi2r5K2GGAMaei2
d4kSytciAg36Lgg81pTzgUb9WwrOoryOLb9KP6djGG90gA3wp9nw6xrfNJ5Q/HiRLIDilLt18x//
MJgpZ/qQxYapvipz6YQjOxEdYr8yc7gOFoRP+c9T5gdyZqMipLlMew4QRstLc71TSHZSUKpOlCL9
/K2zpLDjFlYrGHhasXGBqaQT7hBRbmh2VEByE4YGlu0ApDT/TgrKby62PAkBT8lBmyuKTTJx+aes
6xv9hE95UrBT6dUsQDUC2TTpTnj5XRKfxx/WxfxgVBsB5S7yggmkoFuqbOjJkKzUpc+Q/6QnbAwU
f9MheIn42IOOiFNJ2Qx3PaI4qGyt7vvU8CMwiEVYXFXk3JUqTuldtM7qVjmBnPHcHRP/GlICmUl1
AIq4TkiKjNqYfXbD1KAW7F07f3n6tIQhDMQJbqvueP+2CkH2ukGpURPLJYIltzo9GrejidvGkpYM
LTS6iiItmN8oJncCH7MEKDyvag3qoaxActV8i92tj5r8UoRF7Wr7YKD7Zeko1KgJIra+gG2zb2EV
y1m69pst23H5pDk5R4VcT9NfdP1aHO6R0M/J/0LZwb5ipLLsqqE9R6OfHwY1ftelSiUytlAycplK
JHkNFoE5LHqwCFwpjZZ+g3I22pSTEC0FTIT7h9XO0K7VEyh7JRCQOCthI1qw4w0vs6Mym1j29ck0
a6cuF1H1UJTyS/t9P8r+hqEVDhuEwJ8hEO8QNI8bEYAp1UPmoEMWDx80kIWIv0EyAtG6GC9ahj7k
2za5P6295MCxLxneocXf/MY5WNp6NDAY2bxlkAgcSCy9EK3TK7Qs1lFZ+LuzuwxSMoXnHbdof+sN
siP2E8si4FT1VXlj7I6YBD9TY8m/mIG7AukQOK4OaxRJUMB17j0tBVE368MRj2lFF2813aHJhflI
2AFqaRaTR99KNAQ4gNncU7Qv0WGYXir4DykSxuPQ4DdIf0+VG0//j7oHafJ4zQNQ9XndZdA/9SJV
QywpM5oS49FW95QCsJxVrYYGfW7Xdxi5Kz18JUu2iwlyhs8ljEiF4cNDZvdqQRnXY9AfoEnHurUv
VOdIqSmMmNCzUcdZ0Oda8DMdP9nbOhJZjpqBHM0ay9WI6iUbTDI7J93kCYaQaKkeREIMld/Eoffi
bEE9vpc08NzUc3rNVNcgW6gD3jLJ0hHuv07MzXGGRijyemR6BI6Phjyg3DK1y3Zi9g26hSFrEEH8
iDkYgnoFsp8/9KPsmWPIwg5LdG3C1yfJlx5L1+T84hywjyB9BNdc6JxajWd5FwkBoSqfIzXi7u24
56gln30AWsWeLPb713Hq/ZZXrepVb2mFRWMNYhkbtTqfcfMgOYnEaexsUmHUQX92clQ6bopbZhtj
brwNnPT8KPTo7naqNqa4oYH3MgNf+IPqo30wwUP7CEWx9NLBdcLmw+0GGvYeuZ9YiSMdu71Seegq
o4HF/xCc8GY/y2GEO0gY57Tk2O8nXRzLJhbHw3UGLu3q7vWp+gJu7DV+nQyRT+qqeKs5fToAdJAy
NF9UnJxJXvK4Qbl0aJ+hThLSvy1sn9Ie7Yd4w7vMt2WsJqZrUQKy5+gcJjJ4iRdcKXJtXE7fI0zN
hQE5lagmJr/JjTFoM9SpNKuEg1RQKiNCe8Pmrws/fqTqMIIcxW9GkOYMeZdoTPCT8j/Hr28I5zS+
cruFksxwvOh1U3Sc4AO/fwsoMed5IkKdHAZtwggfjMDDUoAMeakRSQXaNYDJfJoEQ00L7L/lXzeL
E4/7weGW6XFvDX4x2EAgbD8kWekKC8uBN2RCvtU5eUObL+flDTlp68RZDcsdJAHbEKmEdmdwnYbJ
qeJKEiUk9hKk1txWWy8tVhKKZ2t4WAuV12WqtVAdVDTVu1/1yL9J4ktcQC7ZZY2c5mdoadX9Xo0q
z8cNjCzq2mvN9q75ADnB75NpOsE6nelwB21SCSt3wgSaPmcam9kMCBIs4yzPFSEr+FbrEa4N2A4y
9JbV+E2Y+J5EGphIr3E/oy3rJQ75V3I0s12UgbFRLQHTW9rZNZW6nDn80KYox/0SFsnSQ0x6v6V1
KDYrXsxtVQzPiHyTxkqPEQOh3qEcuUlpYR3K/4ucSH0R3nzLroe/OnEBMX7Pmg/kg63Ib0sR+jLs
L5E5TYNSBxHjoRinKYWzhJHQhZ0FJ/+HWD+Jpti7fCUA1+C9Aq7lKySS4MIUtuB9nvpFXkjdND+h
iLaM00MHzG6/lqb/n5e4qZig1H0garQ3lVKmnTFYx3AkgtRtyxzV0iiGO2VmAhqeG3XaoyMvvREY
fwJnG8ZdxQgcdtSBcN2WXO+zUobDkAMgDALojCUtPVnv9e6zpTJPZW+RIuPd5+Bpf/4P/RJsdV/Z
uT2ssRco8TwKq2H6DBD5dzBPNd47Uru7gDAmCVxV4ZM32iQNd/pzR11chwfoK/HXcGigtMGmNsps
83ULnm7Xm8mSJbhCMChThr3+w5xbINrTINYpTffOQ/77sCzuYtw9TKThvckqf/cAKT7GJpXYU/Zo
zXilxecpVYOCN+fF24rexlkom/aeMsnQ4C/aLBRqts7bKocaJNQoJEQpdzBKRlekbh13xgG/4m5I
PAQbvfHMO+0IIBgAvrlzrxzzWWSG02Asb6zgmZzogJOVo2D4/DnTT03rF4qL0uVQD8Mmm+jOo9i+
tbk7QWyMwgz4jyd/IpbZYP3eiM1o9Vz26I2Z4ZaR2e61oFwrFe7lWECFHDQ3fBE0WFwtAXjhI8uQ
gtCyRSRHzDJJ4X6Ndy1JiNzP0v45d2uzg9Tm/4crtdTa5mAU8C5SHrzYU30jG4v7iz7DUuj9cwXJ
7aYacgEeFJq39XwAJrZfWFsbAvJFlI4IRCtIXXMFT00aFpZ3uZAA75rzYwt+a4W8lj1iVRURvIOL
XQrKOCl5tBwzQqg5Vc3NoidqUbkInBgGDYjY7H+iqn8Wo2/rflwLGqe1ki7Wfq91Qg7u3N9xy22E
OInkU7oYBB++/H1kt6zSZjwLKcztZKs3U7dCfHlMLoykbBzf/3DNO9lHH5Vg3VxDtHdpx/8XZ46t
ufevq5jMm1s3HiyOwlOsDZ7DuDP9+N6NjCy9iBFFpqvHlIgwYswvnYZXjLQ+TrLdp5zxz9nY4ym3
oAypeIC8j6Mp4Lw1hGEDaKUR4B680votGSkhwN2UUo56rd+HtKXMZJDQImedhAu0J3eElyWDawpt
NYNnMKZhbEgPe4xI1mU7zYD/5ctEniYZsqbay2Xi7QTTHuvpam4OYKeWdSsVYNBWConFl5AI3odf
uDqawHPYF+px7S7j4SUi23y23HXnGyuXS6sguvgATDLBr2FOusQn+B8RzPQoqIRDdP5+J5OJGRuo
Q2FlOAXE1l2JAYdgECB+EjaDvks3IOF7wVnh7lSlNkeOGSomjqclLPCtFofTh3jSgfLODF00/Sw9
F9zQiN5uV4gns8WyOXa/e3hQkpy9Xi4fEI62cUH9GEa62j7GBLP4m6Hf9KDMqAsKQ6v2K9V1Rxcr
YQFCbSZX2aD4vhYWMRNHTE4kJ0KbSMVizqSp7u7ZHERDeGJTZtjsJS6N+G0V6i9vJXhHdkPDCkWR
/U0PGvXbFAA8HOEN4RfOqoWJFtLitVKhV8RzbVzrpRJTUi/R6YfsgQIBr+LUTX/qXAHmshJQawdM
07XuwgEhUhx/kyV95ozzTc0oAOCIpUsrl/dloT2WXsg+P/cZHlo3XrwMT7peQO3FqJJCbVO57eIR
elbPp6zvhayG1bJsc9oWNRGLrcNlbsvAiUkVaMbcAXpxIwV+ZeaqTvv0q4DOixZdMh17ZpzMGzdw
GVcjctdTBIkZZhOCsUNLSyD35fLBDEGZOfYpSmsLkBAjb2aYKrKrbsTxPa34ZMP9Wuou+jvLgqJJ
XQqOSUkxWfTiolUlsyXKdRfEx9xkuwLeeG8ZEsKr9DlL5G52TRl1eaCHTObDh5GeVcxttNN20Q4q
N3wVr9F9dBsnDmH+ureItI/bSF8C8vTiUETTn/ViFrDIDKo5uxMphAvNJoV5a5PDrThISrQCUJN5
XJFFtVXXXEIo1gK38szgRO/RuNeEVN2KSVih/0rFOQR9eJ6LKeLRvtj6ry9XURXJ3uDhUL632G/z
7oGBhv+ueDq2cI+ISYf/nhvzF8+ob1rYW44YQpK6yNbU28U5mlcPf2oUfwKyYWDszaIHzrwOcQvB
77czKpJkCS5vVKW9+u7EriO9ElQG1vf3os5kVh7NOpLpz8c02GBLWo/AoHgV+7HOtnYsHdmlTsvU
k9h66hTkx998ZY8zL1C0dq10ZBC7O8lSP5YzFSuiwCrdD8Cw2lQaHoEFozgN3FHmpl5R6zH6wFXg
1jKDibWzMB6In/cGRcBaDwyr49GrnSAckCZwv8aEeWhubKpUSbhRZQwLfNVQp0379n+T6Jhs8WLz
TzweI+IaBJmmXW8g/kvsdiiWXdNg4OfYGXvipDOFTBir7SazNHQD7K+VNHxPo+QYxVNw4h4qipJX
G1tB+rUwW//vpV839iIp5holODKvMJWHqMMjgEoaOAiAzQAFr21IPQNJmBJc0F6W3I39xKREWm9L
Yxb3smyztmUPnku2PmFQ4UIhp/8LocUbDbpvr9RLwSt/1CbsYdfCrKsOPgJbUiAxAohDIAY7wVTq
9NiUkn8lQn+87W5VdHPBg0pcOW25I6D9/WAM1L0LO7v/c/t3L/xC4LvKbFWXvQDcgPISBnh9k0Mi
E4a9FMrLlFNv9byccGiECRSIP8XOh1GKrisojUehTViWV5sAsV89oWIO4yEzVr6hcoKJizMHndUm
M7FumYErOJ4fwKXLiW5NZbDUI+HA1/bsjVJIU5xBToJR1FPHqJByKTFrCJ2u1aqJcjVw/jUoLLDF
Qz0U7kWyyR96+Q0fJW3vq/+K5Qbg6O2tC0WuxJmb9uj5uhM9miT4aXnP7kUg0haYhnpV2sO00qGR
wJiq0Y1+/74ksI3xIsaZ6j2wnXNYSRE1T2p+9D6pSgN7hIQm8oZkNX5gb7PhSSuq9+HSbIy/Xgv9
vorsNNQWPALB6zOthtBERc9iAFRx66gt5zIFePy/ruyViIMIXCf2cly14O4pA2bfPLRPB44CP60f
jmzarkkKhSEdTMn+cZX7FGWWCk/IY0547KIOsPafSyLz8naxLDJWvukfSzwTLy51socAQ69tcojK
GCgO2hoRDl74coPGk6FR2ykT8fKs9wXG2n+t43TJL4jV278Zy9Esep3HgVCBNqHsYhtxoEjzmA5+
hR2lcITlSe7F9D2kDCKOoY7F8ShPo6vB7fh3uEsrZVeHlXgQYI2A0WDg520gFRiy8mlGV0cGSGOi
5OQPGx21hs75SWbK+29j0NvXSNv/E5u5QawrOLWkZ7tkWKattrKPZGwjZdnS8pgq3HmsL9LzfZs0
sHnDy27W5Ur1UOrTZapGhyorHVCxN43L3t8FYNEycHi9NDGesdProXRvjNNfKonOTKzDn+YRGliQ
kfskiymLbbth3Zg5hk6AsZaYMWjfH+oAQsMM6r3awz4UpeEUXwSX4Y4kBs+WhJPkvpSAYQjWNIAG
k236y1PY1455EA3NXLj02oPy5jksOF8X72GobMWOFwCtHhsUUZ+cTHVmX8q/o3N7axnvDNT13AhW
iZPm59JrSeSPBicsnBy0EZwLuHfukBx841WzUqQm7/4fHhEmY+UUUT2MFOT3dqFIzbOm8gx4Muu+
x0DCq9NknYM56xQt2S1e9PMaaJ/zDQiLrhz96UdavkYVE1qpcJXUBocWFhQGKdc+1CS80tnMsJZM
g+w8D9OjJIVIQfRn7fUqNjLyLd4HvO0TrrojDE7UTWn/5Uk4nqypulrxMZeWj+O0EdQB6VC1uKZU
DwXEdzu6BWI8tO/RxNazGnZy5LWGW8ps3WzSvBJLtBoYwGwwUUDcPhfAGv9I8IoB5F7EOZNsQ2w2
ggJb4RNKcSbqugjJnSEQeZ9hDsf3rMaHEvF5d6XTwA+wJtJccj0L9FmdtydYacVW1hTibz/LpbcT
RahQC2JakwULHsk4epe0LjBzGkcX9200oqa3ojHZUP1uvN24UuRdjY0AtKdKqGm9H4xQLsuahMvL
rE9gh55l4iCTALtfI5Q3YPGqFRpbs9t4hueImjrWmzGcnVW4ehtpnFP6KfxCgniyl6gZlNpijlXR
/ZSjf0xcdRZExCxyHGaz1/J0e/fC5zKguwyrA4KlsHwrxqSUYvRcfmKtVruYcdTqfA28JExdodrj
QFPY1T+ho2nnPtLlf1H237IUCO1SM7wqhnIWZMVJz1nxkyxV9O3+BP+G/oZDf/FtFixloBVnQiMR
kVYAsKWlrnct0S7kMRJvxnJ8M32GydM35e1m08L/iy6RhHl0OlAPTT1NoS7u5M9meRl57h8JcL+t
oUjib74ATHbEbNPbhP9pe+rseKgLCz801OvvBqz7tjemyXFm+IHNxS9x6r1V27/hsjgZnZb3m7ND
EjriJrH6PrS35CUYz3YiBGY89ZYumwD+1A+lYSjRFe5JQ7dcqsKg+0UGb7h8QRm7VcrvMkZPBB/G
j1b/YvuCYsEVkfL/DWX3iwKunFikqmsrKG3dGd92IOd4GnsLfaZ3Z1ztQzxRKuTpMbAm0jEqbGOk
/+68qJ7JNY8XKTGYqoiTqXag0oLBPmqLVNEyN9ujh295kFfQlTAdOTZgQ9q9/0jtH1aJguaWf8bb
F7ShLjGQnz9rVCs9JF8OUORbWeFPTV3gNhhBT8bdZCNFW0gML+HkWhmErxOKSqRh2JHSPojZJ6v4
xDG/1wsDXL3jc7kju6tmWrZR398U/1YnHxdMeeCAk7OBeCuevuThRHMEu7NR+F01aU889GSNw6lo
/TSy05y7JzS7rvU1IkSPkGF240Pn2EsNhKkMsGKwhtYVEoqTZL8V4IinUKzGtldnD4kYNfOtUx51
DtlwDxLuuUG6+Uuae0/mbG86lfxIBmZCcj6xzk0dUn6FYiSzvDxXr5e4MJojgzpFfBkEw3f3TItK
/WtGqDR0tuI8Ko5xt/W4l9jTJ3vKkypNFMZuuAKKyogJst+xpUFE0nGe6KckyCg1+uvIciACeQkY
a8kP5TOzgcvBgA16k8iR/DGSH2NkZCP1Q5A3pkyUftLnUmAqTibwcdnGnvRmo/mKVs+LGmaenpcZ
KQu+oB1X1wPZbuEWAKX6SrAx95r7aTg8MRoCXwtKapj2NFyg9RbAEoDq7bNbPrHV8mM9pv0M1vEa
tyS7d0YiCxAQjgV7FhPvaFvlFtC92tTqmGnJHXh8z9tg5AGHS9nxR7t7nyjuU12zybolqAVE9kmt
zAhOinw+bayiNAEz1jiUBtVgEa8em24AQXAiuPHCsO5mwyvKigGddTApErNEGPNSHAaVKus1Wrfy
jKrvfPNnldgaQU1tQtnTdjExV9c7xaPP9VjOn96nOv5aESY9RPvaRv5/8A4drCFPjRw1XZ6tAwwY
t5rE8okE/zZVyHH4/tKtCf8n7YDSjtCXu0QVO94CqBb8HGl6JWzFAGW1qXdLJb4NfoYfB/FMkSXu
k5WVv0g3F1SIwf9Y8WecYLL4CnnA0qQoQTdbePONX7L/G4SY+iPC5nWyjc8ni/fEXuCxpp+9m601
3+rC99Gcln8uY6dgAG3TsHRvWd8qH2QhSuVjOs5ar8dcs8RQZYaH9rO4meV1lo5hVEAIOjQkdnXO
1akhHVuAvDd1PnMPWT9U5yNfMOV6a3VIx0Qv+Di3TnSXRbt2DSRz2PzD5B1yBlYh1spbSlpQ3rEk
oZ+MwUggqnmy/s5qdMTfju6Z35Zf+9JT6zTn9jgSgWA3ktP6URv+w24rs32k6oAvCfjli8sIRHRr
XtnqlDgYK4uCH3vK61Xx+n2S4uiskKgBFsmbE6HygPLRTTl7pWQkqnu/Cqfit3RMCQXys0biq2qO
pn2DE6LIHmLeOj2QSnXLRfhHnLtqbDmwC4f7FgJ2mM6Wva3/D/+Vtq3UG1lzNYaQ2Bd3Q0nnJxXb
f76Nw07bMKt9+i44yzS25sGS9dfQbSzRYejoNSyUHUBNwJbYOWqcXv8bPJYecFCWpJnFI8HoG3h/
vvbYdwxEZsZzkdzzGxKwo8Tt4UJW97vnphbT2WMv0phklF0BQ/0PhvULYlj6W3RonHytqR24ze2o
OHw0XcA4Y2/rbKtYp/W/ONg9KjsU9aX0eKK1eNMfkws2lPn+mpaf4IJNpneDHGQkjRgVQ28WL446
EaO6ENR/U7zvuPYbJjUojZIHRZzNZL8E/Juop8mA4b/zjCNFDhIvoWSoot+QaJZXfs4Oh5i1nmeH
jrC3zdPkz7ku74s5CLzcxPYmiPjY0ZUtqmTyrtujJsiZ2fZU2ucWrHViEfoHQdiLsD+8/AFi0xZe
5YcbTx2lkjlIbwqD/7fWOmU1nHOrW8QhfLD/KPR0+8rR29VZB/TrooYSUltWdTfXNonzx4fuUaVv
rQ1aGsFXFScWiF/DUCO+uCrBwz/efD8e5X7lcGhmpM4373UKlv40uDWqLQN9K2+PHALXyC8LK80l
o8XrlgP2cLGx3ocMpa44hBo6HoE7cyP+g88qgvGc35bFYae7psKtX3+wB2Jr2+MXKkgQEJaRv2sh
a8iziKBCS1yBLKggyCu/ItTHk5vQZ/sUwfMPa/MYip2ei8RPR/qPRv5UGpp4ehjlisHpkqGpEvIX
WUV9ywdkMT5nB2P989IOg93DPeqtKfWxX0rRDaAoAhqI/KP9WVs7/Piffd1dfuN2ZS4vv+VTS8Gg
suTf0fDO2+xbI0f+BofrrqtkbdQuz20olvBKSuNJlGknv5qdZeaBOQCsbF4Pim343YNnpDutaVjl
HqfSol4jCaPQvoNCJw2OrJWGPTsrhMR0frFGzwR+v7/55KxWpFURUty18Dkiv7V4XafKpzGXCmZb
tkzREBojXkRupqeea+HfGyh+fd4f8QyUwtvFewkr3wcdFvjZCJj3xGgdbpk/Ztl/rila0Vs+Vn5x
n9Ohi/daKVtQ8uLp5X/1EeHcADOy0MrENKXArstAOxn5wbq+KoNLWZLwMrnT9Z8422dVJEF3O/wO
wUXzGVAULdTYaREFZNuhikqzS3H75HD4LXMFBxmZfEHkbfd4/vpeb+vGi5wmB1hOMLZsvhDIDvT4
jIC9zeoN0UnT7ACryjE5Tbv1/1trXxdWtMikVSDRHMladpBB1IFdhWMWqPd0k+cHEZuAYKtVY4KX
5BADmP5Kcn02XUTVJK/tJwXnmZtfwamlVmc4Q+DxdXzWNgSXI1Uq3eFgtFKTojlK57sxFv980m5d
zAlZloHNudxwUo2U9UjqQZNNRHJcbfm8pA5JqpAepxjMo9qD4IQiHEfvHPtNLdFIdGb0jT95AWIH
2jpyfqHc9uKGulssn+Mw3fGCBQ3Px4T2mGVXMtB64fdkbHWX4YjEK/jhp86ForPzrKjyFQt0KSig
SBrKTx4GFsM4jASCKzg5QVZUQL+2UpWJG1ifuR3DaqEISjUZMGKGBY10gaIy5XNfw07Nc1v95OM1
ry/zdNCcH02dSuNKqRkniVAHpI9OCX/nfhcVKZ8CaSC3mTXC13nodF/QU2jPeZEsC7jroJcnYH3C
tDcmBuqHc2DsJDkrvdEDa4uPGHaJ8yxAIycMf1WG0GZyt12GQ8q6fR1BXf6SmfadUmsLgsCNx/vl
Da8d13N26jbXny6vOBB2hmi2utMBa92ZNpZbVAcHuV7KufqqVwloDX9v54OsS8ZvPYptW0J+jfsG
MQUARsKWJiqOc7miLPbX2AHVJ17GtF4WYIMRnjlkd1uuRsI91OLVpBeqgOb9fsTArqVRIv/7Tu42
TGRpjwQnABj8dWnwl0wVsqmNuOnX3H3o9gQJWQZmf6p9qvfxaytx1ppo8mGUMviXAMewP2SnzZg9
4D//vg6mNJWTv4WMVTaGXC1NWlsLdr1DzSipJtzAc02CrAnm/LoJg4dUCiTD02nhnNgkLy5FBytB
hsOaLE29j5ONFyQED2vpGNYfFqHqAwN8TLDkcrqColmO79U6acmTa+oQJjaBBK6LNYUekTwSnMky
guIRW9hdlnZdkghQib20+QYfzhJztqO6f1DtXd4Tlkn0WiwQnyfS5caXFFvnx0SHksHnsTpA0lp/
VrVno0F0t490sv1xaeLykulJf0EdxnkV/pRG1beKIlKwTYnNizwEqANvmbV6WeejMfseWB4ALV7W
ASKe5ijRvQx/pMwoSiyHyFE+a0q+0s2cncA4RUWDZmP8T6OG3DR+fYpUJTfeYNeeho2MkKpPBZcz
gq0nZV2DfqAgvL0/fZjz91UYxlcZ8H7flk25FfBNZMizDuIvjKbH1t3CK8NO9RUVb9cSWYiPfqqf
cqTwyWhriFMf1T1pqPNhRc9hTGvf03r3HjnYYvLfb1Pnstn3aMDDDF8/ywSs8HxjHGTuJWvYD3DX
KXB6QdgSikqQ1l1UQbZEph48TvHwyCFHw3cOY6/aPZwSnoRKlrvS2RoXu93OP4x/Pn+qJBgsSwSm
9gcwsS9zbA5w0cXhqeBi/sWPQHerJcjm+lj3UzhHraCPsxkdowtBIAHNv58W4S3OXGyns86mzEo7
X1nszr1stxd14bstc5vJh9dxsQuMhgZXgpET5DeRGx8TIDttc+39Jf8QT/U6ynrQcV/tim798FRP
EnhKFU7xVPD2744EftB8PvZVohjMaRiFxoNzv5UOGomFhOiIpOlo4J9c4UmQl2NFDj81DnLK5vDz
6QmfiCdwFLXYP0xWk5TKxcMEDclpFQVVSTqYb/t/TTTgx22ATP10nk6HFTY5G0nlvIgzTToeXeOH
T7gKTdUEDE4XfsvLlIK/U8mGmva6F+MDywWwAhVx9KsNzliIMmk8SBBw+KgKKf4tCVE6p4uMK6jv
HYo5OxQ4FDeFbn42Uo0l9W9W1KeGEpBo0xynu0rkXYK3DO5u/INU0q4BUrZPnLN375c3EUE2iC82
eJYLgsI85Ri/la2XZaJGCM8bcGC+XLakAd9niCv/dLuNErNWL7zEEE/LPrUCrPWQbNvZ14Lac4Xq
70w+WyFXRRDhFzTCBLKtwjgGY1FUrNDk5IBBXGfbJ+mLrj7T6G3+R2QKGLwCvJZRuMJAI/iScQCL
QZnen3qzjMvJZ/uHVB9KsaclsBdShHdXzeF+vZuV08dELH5wopKDLJnImUFKh6fv0Ja1BTvWYvZ3
6Lp7vj5obhoSPvGmgF+e9GnlMRJBgt1d4rRDrM/mK2NPkyLTEiRHEF9+wrlEuwhU/mh1BJt6tIhy
VizsrycliyB83UQUv3EkwBvBQOXC0ZHf7+0qbVYGBE1nCHuBbu7BIDJBRLhfBVn2qC+LWhoWtpXo
fJWl1KSjXTG+14U3UcVy5pyzy0cf3uvYBU/5vhdgAOX/XmnNI0hJ+9jqgWcFFzfOxKLRLVR6E45M
fS8qbOBXWkk2iYa0GDWjjEQpOuphaF1SprPq+uAfQq3DeKP1imGJS5gUSCHMCpxmsvPNiXksAxGy
s3XYb6OzoLFFX2as/zbaYgqX2SCEx/9Kdup6m3S34kHBpEibs+i5N0OsA4al8aMJoerz1496a04U
zQRBQi2LHRZTmIQ9Oc8Y1Ghzuwx5a+rOEzOcUirLSkMhc6BIfgP3l7AlWAJG8dKk9eBpOlVuKz6d
4G8IRp+fUt0H4vOK/54MBpDwNpw0gW/op9DKvuGn7Sx1iwVk7ZK2WapAEpaL4IDw7AnVZss+ZLNB
TklCi6itVvxKuUTHoBq03horVTIBGN8QwVe4mYIfXbqdak60nPH3wbF1V3XIIigGZE2zDs5N6ryb
wd9Jhcf9IbF6SzgyHyixUjNJt/Rk4jxXBCjwXZbrzjQKQgsLMl34GR7FY4V7jBVUxXvZ0NuSsaOQ
JKYmCu720MLAy223D0rXuitKBTYMxtcl1yf1NuDh/DOEhN/Ms2UZ8a1u9jY5ukYail4/Y2y8Kadw
Ugk7TZLPDWLVwYQaPguiOdnAKaf1fFZ6ggV+1vuYRs4h9bM8uTXjXFCiS55bQqIzlZxKZIMAh7gx
zMUOLrh4YcM7hODI2JTHWYV8D2SttghDSlRFCiKSdTXXoEii3voBCcCGPSd/EPKz0mprrddPiFUU
kRAu0ltQ5qAz1rtdUQum5MDK2qCSx3M3CQkrm35wdpOsgUcJG5aIGBpvlqaUlAC06XPfRnbAGR12
AqkKsyMOQTEWzJeGsuT3ieIqfmkkuOi5eFxX8h5XbPQgZ9QUm3YfRTPI/Ea3WyiKwU/tHnke5QmH
G7gCGKYrYDSoEYxNqa1IOCD1WyKOIf45/jVkQwRKXTad+JYpSOTuCL7FPlRffAd7y24DkSqIt3bC
U7bVe1YSDq8MmoWwEjKz6DUO5zOE7X0wniYN0a5QvdqYuXtlQKSZwh1W/6LY+/Gec00foVDP2VvN
EPVrg5lQjCkegOWBGZr46xl9hI/3J25n9vlQSRPcpzUuhuqrMWtEPsBs2z8U8N1ljkZaOfytnjvC
pl2bYt4PBj4q2lIsddDt8+P+9T1IydDi2kKbnDZLdfpa1eiWWNILrjcqi9hPPAhRILaIKHhCBc5e
wTvBMXTiO9cWUSAFHMK3uqGwLaGWkx4LfmREU6Cq/+fnJkmCVzpC1LcdE57kVdFfWc41Rpa8iY0h
EkVzZHqA+BpdwtZ+zXW2tmk9CdidbDojqVjgwjEnh7ci41ePdO0ifOHPHPfVBcdCDj0XjOAJ+0EG
8Y8sAj9JWMjEbaHghzytXfDlQPN9kYJRtCU1H7+/Wv3iU1+/ovMSow2eGLbwAPlJ/Awq5WlppMZO
DZIjXp/bFLl/r/17zt3nFLtj794A6hyjHSWtnM3KH8GyNIcSrHDKODTsl6qNxjFJ25LjAKSyHh4O
ox+0hR/ogBCt/hAlCJhfgVjvmF+JcN3cSntq6keAUeUIRrE6LtJQhXZyUxBPdWCasl0zTvf6/vt8
WmHWWoZaw9Mn3atz3yUPPcrlJKhEiHxNuX1oyot8zlyQp0ofPyqGYe1RloWAOSK2ZY+tZEV1lF5E
j/XlcSAdc7DGHFG3uB1vnI1VU81JrdhqhlVJwVkcqivjG8s1927Csav+secS+nRY3XBHII+Yuue0
zu5tQTTq9+riaR9wmBCXD6K+G2wfm8s5YFeLK9yxEbTKYZ762yFBLDJtBs0bzCAA6TxVWd87QhGB
/leA+Y9z5zA+UKZOUspwOuOqik7+BEe2UjpgAqjDY6qa623a4bD6OZY0C1hsqyT0ywKPn+XObHUp
awou6mtXGxZxDO4ztgxZN+wQL0x5nWbXwSLqQC8Do/vEtqcC1Phfv0pjDZ5Tqcs32jBZ5RKKFCkN
p8P0K71Z5VM33fZc7Sz0zY+HYTUOLnjoyHrSEtJpUKfk5E8eOF+Hy3PZB23cMou7Q+m3xgt72XUP
cnFjWUCsyCDcbzLNQ4QRFWZzjdUz9vtIeNAi2VnIHA9lcY5oBVXgvVAMC3rZFljLWH5t3+NnsgFZ
MW55/iLjtq7IHAwVdPCPrjGDKrFVjSjzeRQfF+bxHpJUsZBeah08Unx3TSEIb1HxoqG7L83G/E62
Ft2L6fwnND0kN+MFMQa5WjLzY8rWzyb+9a1eaU/sxsKx2woAVdvIT9oWXu4vLMYrqRHSPf+a+2iV
kWqfonhVUBv9kCJj/92InEtnLnMT4OPRrVb60sEsXUmtU9NYoWBwmLvaHnPfN9jf5vOG3PQcPfGe
fG53MRdD5Y9aoCP7+3SS1L55vh6Z4jHpcb5h6v4Vl4JDryDjEKyoiQUi7qX1skz7gEANGWZNF/rZ
zlz94VvBk4g3k2jW587ukmbbHqU3wa/qYeE+nttXptSFEVajYO3mkCRF6kGs40mGHIrTTF8AJ/ZM
aEw/OBJFxRHFhaC9EHaJzE47kysUIawG2z4PME+X/07lE6hVzvdwQ/R4CgAX1ULx1CVaxJXRLeEm
AEOX4ZGZyRBmt0TSea93eC7walzn79P5VCHqm4Keh7F6azmyHw4MvPLu9bWli5IuF3VOKylvX/uB
jEZSBw1ZJ9ym9QaVN2J3PTzhMGRzLLdDSbZASk4DSjwOm0oV1FCd3WusgJh87w8faROq5kfzfBzd
1KyN0IBoRskgPgDbNA7UUryMshf4+CUpTyqu10k1Nrwv4aaqBcAFK85vo6INYOrKlK5JUO9sxo3w
m5QAuR+GeXBgyF+Imwqv8ljV7agrD31zGHbpjkS4DLZwLeyrEpotyFeUjLYtXXLiRpxFj3c3Wh9b
ZbUkd4H1kGKjyDZxr/PfabzykRLA0bYnij7dw6ktrMh9QLtUo4OkdLwuPFtqFBPylI1UHoeN7krx
jQq+hHqEg2gGK5VrFeLi6Qql4wQXqEx+FKZvbqOYF/deGD/TEV6Vjrawt/IrktzRQn+PvL3gP/sR
vQCNnxRB1P04eaBZRLyBZlUFtVhQuI3+i1b6RP6WAymTnbRfCk32XHPMZSylLrdEmWAhxQrLTuuM
+ldxsdWh5fa8veZ0+BGauwIPFm6jX94LPDamsnZkX4bBbw8RVkacmoDVTfH+CUMNMeMtMNusNPuz
DMVJQM9/hJYIdWpcb9fLTOteCO7OFRuFcenRqriEJYmMe8oBykeRqk4888Ac9q1rz0lWL6ScWm2h
+8hCwQya2cqToKEasM2Qef5tssU43yZIY3MGh3xsxOXthM8IqejWBQTaYdvytkgjBFJGneTam28t
eqwj0xi6uAAH8zjRhV/EypB/2wU0/ApmZyJ450ur14fA8VcuA7nC2eRgH2jXUL6wSb/hKhI5wYZC
TlWAU0DNh+ZYMn/Xw0LcZ0cbBwUTki8DO7SgxQPBkmZRuJOggfnq0O8JSIXPkKzH8iQO2Ty+3qRA
Z6pIZSw7n85YylygD86sPUVkZkg681SLph/rJARQbqd+mIsIQn/mWoMYd5pLqXJpoHH9w5zG+l+8
aJpsniM4oEemXiPDYCFWWxmmVcDy4J86uJBB7DCQPai9HPfJ6qHjw+W4T2f7aO5StS/7PaQHKZRT
+txPyLt+yJI5brvO0Xhi/eTblu0/FnIwP8BpccX3SKCCxISQNAPxslG1lUZOR4VidCuK6J/S5cz4
ZYjcN0kFTS+NlKkoYqIlMA+Lam9eXq1y4RHC1zopuOLuAccmdD9rqZCO2SHbSNcxFTPViwBdsPYT
LcimYQn0DCe1gLStgZrFyEoceemRoQi0VKU93G9ODmP7bsAyZeVZQ+3956NYrEVqVkBBmW9EWkFS
wpv8GgaJ3Pp9+7vGnl3YXIf1+hZEM/qxbD3e0UfcdpBC5sMcauTt33P4Hv6UvQSpMJTqrO/f+op5
9uwEiVbj2YLFcELDZZa+XJHnO4OW8iMFWprsorrIzlCPqW4L8HpCOSJAjenkr5vO8yjhtyHG0QLA
yHb8yyrqe681/XTUTQV7eKRABeVh4ev/zylREIrUkTlWgVAhYb+qg3ZsIxq2WPUmrldg3jcp6X2x
54PdT5z7P0yeMOpSBJHbccZml+ZAFutgKPzDClS1MzxLderVbmAnfLIpRc+KNSAQcdGZXxtr4E99
nPHa5fLKz49JGgov8CBScLLlSToL1syRAyb2tj2DtvFAQQWsfrzqpQoUBvlYUrbbHY4gIhMLq0+2
Duotv6e3xGTb05zYnVeSneAKPNfLv+6FRgXFno1fri7s6tgZ5bxMK8HIn1KJtJG9pxL0DrauVc+d
4WzvEq6qhM6nzP6OFGe4SZRxokx5eaSw0ZBjVLnP7Xq+qjp5XRVefP3vsPf//dX4b8diJJJsg6hl
CxOwk9d8yTbGhgKAhOMuWINhuGT71yGOnik+BjXZp7+lkYd1lp1Bg8H5vPdIJoDsUtTsaKjRZoED
NdRlScT9zKAXlnrhA1GFL72lcAyg3yXuuhNneVgDRef7U7M673ZgO2llgiDH/T18OlpyYYF/J336
2jEZwS86OPtEXaBZz0ZxPKWiBVMG/d2LwBQYDyve4BCmhQbuscsAdPEv8pUUTpkPFai96bnRF9H2
O65pLq01ZPhYnwR17w/NwjnygC5LY8xADta4tSSq0T+4sykZV2jXsmBTnEL4vVcNuDafMzzFcgKK
H5bJ/eoXhdK3zbMr5lOZEEhie9nj1R52LRhh7bHi09mwvJeJJWnA9fkoxkComfCEIiGl1hcul6/o
MlL6wl3mqK1nn/19lcGDKqGphnqZQ3llHoOEZ0RhG0P76QNgXGN8VyKMtArLsEwgxyhKO74NYeii
MJfTgW0ym2QiUTwfGqk6hGJByAtjMdBpKKoqLBnCQrVFRiFDcJev7cILknJuMWff4NSE/KcUYgqi
QbMWx0EjUVvXtyByGXcME/CYBXsyuugPAK3EPThsjvw82aMSFzrY0r1hWZc/BFbZ2WF+n+7NhM4y
5/lSkr8Xtgvpab8bPCX4R+jF7KB+J1soR0KNaUzdIM21khY/681gceu6+N8Xmp6fIKTFyqlNyAp1
GWHEIhwIDCG7lX3ev0lUTwGmglq9f96+oOp5U6sPBTpJkX1sROsyDoIWrxNMTpZaHxKuNvenEr/+
YeLWdKQ7L2aQkNg/2L3JW0SqpkMlGrVTDDuIFvxfkblcO9izCOxkmja16TrW/7P9Gwj9N5dhfc4a
xJn6Fvv8zkZAReCcl1DSzotMeEZeg4eS2SJSQe0e1iEJQy/C4q4EyQaPV+fERnG/s5HT69bE/CV4
GyxuLqTdL1YQnUqDEyTwlNKntHzQRxYt9Uo09lke8s5zsjdiIajxAAkK4ZJDqzFIqrp1EYU/8F2C
Dzh5MuO615gge54koFNQrKUO64S0ouXlzSsSILO+RPM6o/3pwJZqH1cJKxpwR4eHcCSNEoFXHcEB
aWQX03hLBN5bq12cap9IdpsOtFMap/ovhqDeiSb1U3qg1rnF2JLtR2WI7h0cy+PLkNil+2tyJpfy
qQ+A6Vuj4nxJcLLmgD24Kedc6Lugdobid3woFm2jQPPd8LBjYod7lVkPWfWSqBpQA0ANY7PY223k
93/zUXCqrTUuDLiif1jkVdqNZq4ETVGKvd+Yz8JzVn3gzAwQQCEaxIap7nXAVm77FuvyEi7XtbJd
rKJCp7YaWG5A/W+1Ym7SbLmJA5+M0SwD7/HkWjDFH21dt78EHcjEYK2owYpzCvKONWDp25SGwsmx
89DTrcbypdm+R59tQ2+Xgcu6MDgbLw6URTAgwXy5nPLEkJnEToNQ4VieLskeDHUHRoWsGzuUi7Yw
MvQ4jo/wxJrdkjAr+fNf/rO8DhEdWg9FCcp+oNt0DZkiFhThfh+dWymrwK25cWEATp7m75m2Vft4
lPsvyYODb/8EncbP5uq//21HRmiX8rEP9BXD2ZaCVzlLridybfnJf//WUDlSv9PSp/m9GzwCTTLB
e3puxBHaLBElHTX5YwTFB5XgORYia8rH0s62azs8BTjkBUBAJ2WMGQpgIrwZEnScdcLjSH+LTZit
elez1vH46DQoLb1FIFAT4y+pUXd1x9SAY7bDfZcmYGjy3l1YsMiPJzsBXpExxtoSOPRUVUQEv/4G
Gtz9AYur/GE14Rmw2hwO9ufFIvGZpY6TNOlW1hL1lTYVLslPf+2b0YNlLUOTz0pDwabTG1nfozl6
jhPYd/lhlQ3N7jd5u463MguZbg+pHC9IvSsCKxTmsC9OYtu4oKd1GEJ5E11YuLY44TJ0zS9iEy5k
Uxt5R8BhsNtaccwpw17sRw0bEAb5BvWFzugKuCxmrkmMgjMCSUmhBKPOZV7U+r+8Z+CPbxShtjTp
oOjcNQeQLbqH7vzUjfqEFVO4TngdE9uCiS1NJ9Ne6XOiMtPH/W13fTqFgSFJec/Haw9cEd1rlcfH
rwaPdoU2dcvvDGriFj33NdKKkMpoVyCFyFY7U79DF+Nh8aAaXIBCXPFJfPZoibx8I+L04wx6os+t
5DGhTXLOUTGcrpS5TgIJcrS9E3cfbSnUi2Mi1IAyxt6nnwoWRfrZ2FmWVy0KJF3sWaEZXskr5hto
ukjBmO+PKI3n6saycnNg1lrxCDurc/H+tVYiQxVw7tLMkSFHfxAt6Y+IPKyA0ofAWsdBPfsOQefo
bA1V15X0z1MlKhGO02PeAehzzxppwwKsEjYaYlo4z+afw19gQLirnRxi9b4YckA8b07a6Ua0kBl5
Bc1tnA9/6DLLXYCvxd7+pp6f11c2wTqGJNTcqeYUnwlRGH5IC8Tsslyimlalx2lBM8W1q/DLvfHf
qTq6CD+3N0bEpLwXv4fCJJdrmWZ+Wx7CzrSB9PvH+40Hky4R2cr2lbO1ygSdSOtaEnyB/TfBD6QS
b6aXF1Zyps9Foa4iWXCjvMvmbK8WFw8z4BmefDO7Xot1dd5KaErho1LZ3tR4qOcfFmtZqQ7KhIgJ
BC2cDBeiSEw9/LdeiFMZruoc3izD1lWFYqzgRB4wcob11MwC1ap3f1D48uHhK7+c+wonTjpftVan
mynFQvTe8m74d2QNcQ9NmpQXBBYOlZlygPsjsptSGD7kDHy9OYbjnlWqAqtZBTGKajHTvj4NDgEs
n6Ua5xqE3/V2rSHbAV8TyWc9vuok1pdJIafURBnJzPu9DIgMcvlhyuFYtoCN3mAOOhJwjTa77/lL
zwzyeHE7TDoQjYyBziyMe+DtuivyxdjFSa+lyVFt0MaoCxrvrNLdYUeMVe4ydxDa4QG3W3mxGFwc
v7ZMTJ27C9r5igzeHkUW6W1NRgElk9hTWntZpBlju4V3JloYCe7pPA+og3Obl7F/lN9asBcdk9yz
wAUMQSjxvmdgYdUoH4xEPi2Y8Bh/Oj0oiD5HrwNMyDo9Xzg7qLxu5kUqa1X96fDII3xMJLuRuY3o
Nyh5LUEVQwuHmjNYOJUUN+4Iw/rF/wt2v2G6ZmZDLPHJpmLX0z39thSDu8Q01n38U6JDKIRXLtNd
Fc0IhU3I0xTIPJs1ooBeUU/UYrDVpNK5kgQK+/oPf+C6QCI7+DqnAU5inllqPLzByW8oTznYktc4
fOoggD1QbYjU4vA0Hsp2Ers918wlXh6XvaTcbAccu/x+/1YA9Fxxl7owRB3je3YYBTuFXVnWwPef
5P9mrtGGKIK634QoOKHFWvlJv24mW3bn899nPInW17q2/6VDykwS4r7hDefb+3qdFWFjqvFQegcH
kS9wVatKl9xs9agaQIVuW0pbgbHt7VF7EpiV5N6KW6UFHKbsdlSqtTScMq5ExwwDw+QE1bf6NPTD
4DwfFw0+q239IiYrzD6Ot5GsCLoiJfHRB2MTk80rdi3seDgP2Rt7uWxi6hWK6qDG3bAbw1SRero5
Z71WyIGNUiPttTG/29OP1SVx6wsCTki9QbuekPgaaNTxlJKC1SS6Kq1LabHbAj2f6BsInHLdyDRx
o1IUyp8ZW2EyQTs8xUXe3/Tg2uK6j3UVES4yf3g7/zx1ExoN+9gU23g1nIyvcTQYvrPXC+QZ/AVE
zXNNnsrXGkOq42KK1fwKozq+jvlcIAhpeHMq0sNzcgd8LwXAy+hXt31+RCu2Oz6sEgPXq1K1EF4C
4oAiP43EgXmpEn7l0++rOSRvqcoqRIYKFtxqDe16iopz3mH0q3NN5QiQKzWf/X2aL+zWiF9LfTUy
JdS+6jHhBgOOG9k1fjX402TZki1wY4vDW1smwUH4MgmvqsUPDLUTnYnzBZnrsOl8kSJq2wcxBnF4
rUThRLyd1BPkIaju9xLSgjciKxN9UVzOp/2Ue7ESWCq25E4YIog9GRbteVp2SXossWjSn3JjsOe8
tnof7Yx6ZckmMZ9raMHxki4L/2dPPxeEzMRxjUwWgzf83AYwQIp95tNZ+tqCR0Nc57uOhTZkCKQo
RVGxad+0Ki5Rqxmqgv2ucCnJCWx+4ueOZ48pCPSkTxVZAukWbd0LlGmsXk8JJ8lnP/SoIueWJL0z
5X0x+rz5YDtaVCZPwKlOs8vKQf0fg9ZqEUMGcNElDOnu+8CPJqgnn0N142QJb2wCsn0Pj3SXcFRZ
Q3bHUMt83Ebfpmx12WzcV3xsBEcZWNiA9Lrwuv7FGKoq8Pk5SPdq8wMgydHA9QlCJVBK/XPeVlmr
w1zRkUTCx/1WeQL8y6zm4H1ADnTylUHKJGgHAlZZ9Pr0qe8ce9JFiG0z9KxOGT074HZo46ofNHzy
HTViKzb0Qa5vHWZdOaXSP+ZKwc+1rJjCBybRDJc3A4iXmgxkBHk0uDHIivI3Akbt5iK5mhQpI3/L
gQz4xA2+vhU69v7A1L3yjeQk7mIyQA7upfdeyubnDjXuHIvxskqeSlWwo7662nq5GZO7Sj2dCZs0
J3jiH2XH0A5etURZwRjfcopBOEpSw/4bNZkCnSZ0yLHQFEY38D1NPoZBDrKwQEg4i23a35aEKMD8
0i4FjsOIU/6UsFqmr4Gyp12A4xwXR9HXYzwjLfSbuWMdEJq5xdGLxjT4bDfEZf6h54qgmiDLcks5
Dz3FWuWZXlF5suNpyzgaX6OrQ6a1XuC1whSwGrZe+LM9e/eShsFwyfbGw+Jx49jckmd7/1fSMXR3
11ccTI3OsRTkmf9cJoTcuJqA4cCueK9KMenjq9cfFs1CJHMaLvZv22CQGdcqZSyt+svq6XiMF5k7
TbPhSSilUQx2NhWWz95plDVt05/pgmLymhZnOMYIWDhgV+uoXH5k/ERGJsPQV3c1JYzz8nhlyF/Z
+IelRYflBSgKd041lYPWt67SnGNuEybFfKw+fTvwAg9FOq+dvF+Pi0q5CCyTbgVuQ2VnjdX/Va7r
1h7RrrABxx71JfLr9Ak/GXJQIhqZ4tlLFM+9OlGwCA0pIxLwGV1+nVo0GGw5EtRzYUI/Q+MpU8ja
8sC3pGZesk8Nczvd6XRcNZXnRC9zrcOnEYj4Ho46ZzZs8uR/TUvTxugNDV4RRlpELK/S0IKcf0aA
68syz3TgYpNp/heV+b4hExzbkRWkbarupiBDfaFKTsMj28IaWF1emOYDoieewJVgVqpBkv6/X9Lh
DkSGid6pMZCzI/yvs1AQcn3nDYo0A3RsneAzdnPtFzfs5aV0ongMgRl1hgGyM+hWa7X2o6XneU7V
ZdmS49t/EbDWxLldEfDFDE+Nugc8OtcKoPFMPQ86ZteDc7HhwPc4uiy696RIjPaAgK76E2YSYnQk
tW6FtYEvZeo1M3d8ZqJQucks5JMIapUM/mYRVrs/soqpMVCIUu/bv0OU15lZjU+7Q/uuqh5jJhgU
qwg2klEH1NcQ1MAI3QOJwWhUu+LIn63/YWwB68mqVymdBBvF4xaGZ2SX1xAF29iQL0uBdr2rNAIl
87W4nBCY4TQw2SGr28O8Un0/gqZm5P5sMolFF89dhkDOb5zH2NnvtGqwFmSpxjasPTQjjwvkZe97
sxSH2ldWdKGsdKl9reZOKU8gRcB64fK3OR36V0hSJpEMOIWAFFSfXRAeCZxyS3AbqnFkceyrsDgz
eTu0ece6TAT8WI37ul/ou1enoK0NRkyxHMln4gbu5DKpjsKiSE/4fpE1CJQX4x+Gew8UFS2duDf+
Qjj6rIFbgOA9snzmXflu6dlq/r1ZXDXlTo2c9lfxq6d3A4u6bLJ0FbiyJiBVWLeRXVjOFo4IrsDY
2JroAhUlCBBd+YqsDniUAdhfxrkMUyM6g0iU8ncC4zVR5OMIeSWG/9EadKCInKwZamAjSLSipdzm
2qNSnKWNebXyHdqoS9HYsuiBAAX8/d2pfgvGizMJL7p23ve1x/uBHRMz1k+eh2bvuczFbicG1tq0
ZlA6qjIblUwrKWsV3gGFUAxvVlzoAiPTRqa21UpbzHklAxHodrjbU9Q1dGUhCCGVIXZXObf2BZjf
YE7iPeD0q9aMItxBE5IkC58zHiWCq8wfIHy3akZ16KDaHnXYfzrJz43JowPD5DEQZTTNTu9+KNOX
fZ+8CHl4WZzWq8SedVUBHOFQ2tp+b8v/J16ophONuG7tlEAVSfJ6Ci/bi+ZvXzznToDKr3D+aXR3
m383CEIC66zzkf5toEMjXERabA+QGw97easRQ8ZfUfsJRMGoQr3jcUbaps3lgBnPiBs8QQ9lm10V
/U9x7YQLS2OlNBSxbiqELGClniyuF7dzJJEJaOqpSd5vTcNKrWpcObG2JkGsW5wut78sH/4lvVZ2
19JGhBmdKHdtcT20XG1dkdFkZ5NtUXjuLWX8BfDYwoNPec8NExxb8lcwHtFw0nu3rw/Sxa5Goend
uO5N9I/kS7bm48GsJl/22t72G3lgL8MbupPFcwRqm7I5sl7XrcgSazssAHUiu7cWNVkG+NXv4Fhk
z6isF9zLoGdnV9MtmtKJcd0bh8LFTO78caYoxe50r1PG4NuDng9LpF3n8zmU/zShBOmgo+f6ERlD
GEssXefTpxEGnzvKRQPQx7C2IfhvTjKaaJEjUZ636yE3ckd4XQXNioT84e8pF+xN81i5/eT6v0zA
xSLFUWoaKo8WUgA/o9+AkYy7aJHrqDBtosMxIVJ2vfSLCoBtPLvTxQ/8brOJVh70SkjriNj5/j2c
00QixLd89u5lAJqXoEwNc5FH9pi/JfOYShniAV+Kk5uSqF5Gr7Aqkj0Pebfy3SBpY/vc8F16l5pH
OlUEu8QLHnyBPB/i9u5qhCeb7C1OdDT5soDiYIZhXjanb11YN4F7LcQNPIQpjFfKZ7p0hms1Ft3K
1l3LGEv4ADY+ABLYGKiYgzg1P71c5EZLMOMe57xjfNmjYliQvN1O1xx7KkR5WmY0gvgQZZO2beAD
SEKm6gBiWhrFkHkbnNX8hsOfmOyXPar2Ye4zOiTzgRayzQhU+vn63D7Las7RJ8fFHXE69OKBDkuP
SYnxX6we67Dyb8O5mQDByWk+q59jukllPyWONWjMeikPIPgj/25dkqN9eCDq0iiWXNp0fipFKgdC
RkJLgiKHaDhXXZf0CUdwGECgnBo4w+ccBO4FtH5h5DABK81Rhkt+/u9tnfVa41Oy5e6nkp0Tuol4
3nJLMTc1wxJgneUOqSlYsWiR8BHR7fKigd6Q17cloeYK+9+jvnC05Lnu9RDFA1gixBLsFOSGiGf3
oaiOjrfHzhvTTOg9W7evtegOaMaPniRxAAKQH5AVJp9ehALn/5eWLMtEEG1pXdRvb1jyOI95JRbO
X5NXR5RyP7Xkk3w6bywfDBGd3cIAc1R6BQqE0RE2sQdTva+gKASxo1h4bSzFCckEDlvv43qGGkzS
OuRkfnO+2ylItvHtQdcP45AEgGYSco/ABU8dF0/G1HvARJ00vP6Mw8SDs0GtIDjlbv2W+9++PCY+
FslQaDcAZJ/9mnHlW3uh21BT+UaKu+a3w/EFz6PGrP1Xtjrs+lvbfu2B5Z8CG5phxipioxfjD4WJ
yWzAPmVhxeXh2T5+w3VJ4G50GdA5R0rsaX3Z3dzrHvB5YcW9dIQuM3wlXlIB+4Hbref+1tGP0FpK
v7loRTINIjHl0H7TJ2cF/4JbIJcwUXJTAzO/6pCh9utbWKU9AHNUC92b2yfTqvhIccrWRbJVsSHk
7TvlPp3yr0rqbbB5HMCMvOjEZHMzmBMcJjpKvFuCVGmSXyIXfVf29DZJV1iSRyHuSC1pyqXqSlgr
e3xvD/O+WvELydGuOkrdm4lSO0PTzLi+gXWt63S8VdgOmCIEt1vKhgbotpTpSoMdgGCVqpPvTxnz
iMYcyl38EY/DNPaJzZ5oMmcmut+XwuyMmvnmcr0Oi3UsN8qZ+/vDtvo1R8wmUzi5sFI2yeIsP6m9
bu+QzToI94o0PC4Yk6fPGr9I9nuFlbzcX8ut58zWlX5Hxhe0vl/wF2X4ytwpiHBlhCQGERVPl02U
zk0bb5cx4dN2oU7zAgz6PAqOy6cg6BWKqSNLuLxbRpGMDKrAiyTOaedG7lSYip2wjb2tvvZNDQos
dIB3tcDOBu8G5imthOJDsNukQ9MFGhBgSKqfx+BzLkfidHTqs1qG+f23zfm5e4+s5GO5oVcGqX9/
eCc1QX+tznDAaabNGnyhIMYdZH1wA4ogh+rWSXmzEPrJ1WD1YGWiubaRjvYDKgYOA2TKN/GqYvU0
IdkDmSrYtVM89VgvkQsZj9iq0cjl2McUhwBRMfJ/n8D/aKed/JJakDS60BVxbXxcA2znGvUnN2b5
CcQagIc7AR7wKbmp11F9VazpceQRe3RPdezqpiP7m8IA8hWW3l8zActRM+UiYZXjcchfeHU+434K
B/YIQtRcVd6yZhZOh4PcJxzVJjXNbhfYqLefYxjxdSMpnV+PQa0yVUeX7lpOv1tS0Zze3rbd8eWJ
78w4ph2lFQZ+StcMz3I0lckGjAvQwkTi0py03PB/dsOuqcKI35teU/ve6WQmfG6Z8Rp+fzMz8RVF
X15O/qelpVFQuerT6GBWgSEGw7yQZUZnkBaKTW0g1Q46wmM5GxQaCAi2wxEb4RHmY92SJS0undtL
OL7ObNyWIBelGG3MZZzgJOdFVATQZ3xVTMWROrYaCxHgtWJQ18ll8yp4zUpGpl16pi1s0+5PRFuS
N6NUemQfB9KBf8gHxXzcEqvjo/QwwQDGuatZeidiZXNyQ85xs29vZ4F0XbFPxuBnQAHV8OSpYMxU
jTW8JcXRLUTHsl9yO5CdTxugPL+B3WMPyQwAxi9X7TfIhQiV2W04bDBwdnvERFg8zipMQzvbSKEw
YyKfF0kmwIFjDX9KwHtGqlqJ2GQZdnGpuVNWZU5juifAetGyMudzb3T0Y9PjBsr1NScCW3BnzB6t
5XwvzDG7ogJF/D6hdKWBXm8ZHB53n8FXhZ9M+sESZsZ1BM41U92N0oT+gKW/htV6Wxfgf7KUsspX
4y1gvHlcWsvFpdwIc7QlL87bkQ9MLwbXvydjQwbjRyLCQURkS6kLQr7XfD21c9lJW2Psyz+uo3sh
1y7opzjU2vQAYpgshR5MEkeakXhwkwnREB14VeYRbMd/tDO+IHfZByk62lhalzxLO47VatsDyMlQ
VpMVH4kKtPVDTJ0dqRU10/jF5vZ8JDgepK+jtGBBfJbsh/SiazagoJ120IXkC9cUF39e1QO+s53b
Ewz0Uaxy5GKeB45yuKHoEMzVBHLY+Ra4QLpeH65st74CWqvgTECAByGgWXlM9xRC0Z9oYwyx2U3g
m44KeYSEpLDOxQPvc9yzlpCVB8q4zLLPmBW5z4DJvhTVNRIPxfvlbUMpio7Aa7Ff0HFdn8ktV6Pb
LIKjcCKbQZfLFVtTZvWBWqwZZ2tG8+qKFVWQQFq318UvD9YzwUG6FCDxkrPUpy1J8wrhl8q9bJ8u
vwXmMpNCNxnPa4nnY6Gvm8aUG2JPcn+yQp7usSKMnAaUl0t2aRTna1wjjr4738DwGYKr2GWtOMgJ
PAtth7PMJOXdg5szX21jHwNw+OzIp2iVa7cgEDjYSDJ2hFst8J0WFTXZfn9iK+ahjbY/ArI9WCsq
MFApOqS5gCo5mwi6moh/oN+t4nfY0wu/ElkZkmHWgrZdIuRII1RpzZSyh/G8oSrDxhcYn0pCn2bG
VfFW6FC+05ZrGox9GzgXObwJGBnnTX+b/l5JplztCdDUwRNk9IRak3J0FJIl7nvjculYVbi496AN
nC7qW1lqQMY/jp8ZLgzsnKQKBja3mJtm/PyDqGEMUTp/ngFgIPvY2FS8pHtwvsJb55wCVpwLEQIG
9BLvZ8Mk38h7YDfdXdh9K08O2BXJ6PtP7BRYu95HNJzNR1UEel4gTY/eqc+hAs7h5UYR8qcDpI3Z
kQ1gM+CrZsM//TaKSej+Nl+hnccfYMIGx8mRTWNGfokzuib6vouANK2aRVUkwg4z58fLu+r6sLTL
cNvOsqWS0YIDhjvHQeUx1PP/5jKVNnayqUPnPvJx2EuI/933QohFf1S4RSraHK/mtNHhis5RqBAQ
zKpHITrxoSvp0HAl/imp69dT1DphBmca7R/J0Z7EAoEAPSQrzbr/Dk8S5KD+vBdyVqyQRixUPc+Y
dKKdA4Lb1/2BYJE4OTXJrP0207P9XTlLTM8rUd72QZ5lfT/VusOHX6rNjNeZ3m3bt/h34xLQGGXX
qcbetkpvtFPwYPTzM7PKtLKfRI4lktAWVzCkPIQTQKM3q3qaJM2KP+wIa65UuJiDELFt6iNt38gK
ER76XceItClcEYfZ7+thTku5XKiviLbY4KAhIBkf5+JvKVh0r4KfdBl8KJzyf74rQ4vqmIjagU3i
akM0jDeGyxbXEK7MVPcslJbjzzuaun/2ZzzE93HXv5xOyNbI5dqXkGFd0RkAYCLBR5euuzK/VDiD
8hepk0NAapNhsvIT2zscQHAf8PkqHoa/mp6eIj/KsSHFF5jzzkpH1yXuf6AROZTWtfrWx2qZdWbq
fOewN13WmrY11mJzQhcqwarycLUCcJUuif21A7nxpxnVJMgfnhoGl9PW9Lj+TeyOxA7sKpvOt523
zc5HSzjcOzQmMbQlrM7l8PS5tptuM+2BP6So/s1H2IdpvmA/32XqZiBuRIBN2uAICXXMyioGSk1R
vb4QnjQPdqx51lkUzqjSUQeDTD4QzrAqBvQ+RS6SZITZ/HhU6wVL6E0xP98n9gevCdlhAdG++IYw
FaR+X0dXhYtB1t59JP8NoSCCjjIArLx3cHPJG9ZD6sSHEiJ1UBp8hgb+KAxALubQ9HO/th3+6il0
nCizC9DszK++Le3NmedF3tSX1j06psWZe4RGNviSjrX+GXWINWjax8a8WRsksj8qwy1IF5GQzkRO
kjYrEopjaQfSa9CYn2IjkrbIcSmWJuN07yjbKGdz7KB0oAxNw+MrpAVWWMZIHqyNPi5hpxflETG7
tiOWhgD3i3vX7XADdxX2N2kGi8cCYofBoWdT6kWr+HZC8Mxiow5RxacUze7ImOmnq8AJwJftZHO7
40Non/tmfbwUhBpa/L2woh0fj0XFD586leSHLgJn4tTme8CKCXX4Bg9A4Q2kRPX4GwZoZ4dD3DdS
JM8j4tvXdZAjMvOOyFhVSvXXDL8p3z9bN76eWsZbSAR5STlO7Mjga0bY4iB05D9h0XV7wAyfPpEj
nmWbJogFYByRxCkqjGJjb3p7LT8HGGlKeLwk6gDDdTXmY4NBKLx3III7nTwM9CEOp4FmHO1WTqxO
FcwPNa9DukwMabgS67h9tFzYZ9WzDRQwf8rCbSXcsy3B+rnyl+X7BzyoKWGrNbRCdCzadNR7q9qI
ctZNGeJEyT8ztUyedVNT+R88jE7BOTI3+MtqfBb2FriOvr7+dOjUl2tSAsv6n/jwUy3sYQptIyWA
VUCMzgxYowCOLb2ZiiM8nk82ZM69hBJ8S2a78OUQx3E7fxt+4MaHeKH6WR1m8i680DiBI4CLN3wa
wgmBKCtFe4oMtQgzWyeq7ACnOcIcFcJvYDyAue+JjMR5faPRc2AVtzOT+5hmGux/wwgW7tAAaLh8
vXVO3duciGQxXi7w7uzM/mQGXe0eGJ2SBn5hSUFLIzSsWR2ThHDFvvKH4WKGJK7FWIeApufBKZ5Z
E3nIJ91xH3dA1YA/kiFM1KsCqms9H72ueobPD4urrOd9bN+FkoAJar5DPypMbURDUH59/syVlBg3
dyu0/upw1b9M8jWdrRSMLHUxjBXufN+eRGuzOKyml8+MJwOXArir/BFqOrKwDdem3asjcbUMfvKm
PX48roafrPsyIAhceyetedUAPl6iwLFwWpdOGyL1/Yzf8n2lwZnWqJWHnJEfTEDjrWZmFtDrbmk/
sBnuISfs2G5J6BnKmXki73mynMV2rp00MvXJDZ/MMe3omFP4LkchH0YVQ4glqc+HzxsG+fM7ez0Q
NY/3wfkh1aNKINaCgmcFZMiS1aZi1NuiAzPr1wgezU7OWqVqQzYOGm9XJmeWwsc4tS6gDGpnws8D
KddgeQK1066oqKIXAIXPfh7p72OX4PZM3YbkWwtHjcwtFYjlBXsAhve15vJM1aItYJDQLrlMGCYf
cn93Q6QR9Nee+o5CB/Qiq/N8Y7Y7kDg6DUtE6FBZ+L5n9XvfI+/2s7nvXhBYFI1HcC7U7jWbcoY9
i0g4a2N4xhs9pD71rmRjIUg8k0fehvtg0ifvxURxJEIw9FMWtrYQ3dPpo7LaETQgIEbg1C1Fy6UF
viKG2lbQVntOWOyPrconm5AI89UWCImNL25qqwyKH6GSXU4Bri2EsOU6lboJZo7POKaHjNlVU1JU
9MAnOJGObofZw5dpfZ/1GAP9lnyHPunTo0FVCkY6iHIsZs9oGyXiXsaRl8r54Vz9ZSZ7NYl2dU9M
q4J6eZWGYPPGGnh/arOuXm0oBfGowKnpLKN7RMI7Y8f9lGqF+cOshHOlEHHt7qHsVqjTdyMfdMX7
tgCTT3oJqggx1QJlMo52CqTZ3U3HxT8Yo9swTEUYsGAjV5TdYVnqDC+G26276c1ZJw44Xj4PCyvC
Xdzexe98o/ThhETGFp8vUZn6etA/f4stfeQdB66HqTVw8Hdny6P5fykoglIVpBMFt9fnzUQ087tO
2IERBgArwcWOOgfhBcPi8EQOlEdqq7Y0m3NJdUEhHHAU/RYSg9fuWhVUCf9JHS06w3uBIcR7eIZD
topzj9UIhSWeznf3LYpgDPgY0nrW1+zQi7axVv2wdDvUtGmtoaGsul/pAj3z2gPGNfE9N2Lb4gTp
jltV2EudIlyvxL75pHpg3Zg4Rs/BnmzQVKr0ahg4iona/qB2+Ut9pZeizbjKwnotMAuqhUFAi8Su
mnfD2AvpC7fkjvhXMaOFT0AKiheGUI9ZqOIlh7BCtLIqtG8soKmZCoqjH+1a83O7cH4l5Z+v/nFw
yA0P/yCgwDH/Shw+vKK2SAJ/Wi4IOgZ+eI5rOL85txBtZTxazCh/rGhoM3QD8XCf4g/WdM18dyG1
3tIV7S9lnr395TL7wXhF0kLoKn+W9Z/NbFLa45xWdSkhzeIN1KaaoE5bOJpqYMpjIRoMtKpjeOtR
BHSh+GVYQ8AGZ813RPdqg9hilkMU0Zq+4lx6U9CVxX5Yi3EZTVXMiGS2vENfVvV3VmW+/bqqvqyx
Bn+UC0GAcPcYKRzGtO+w1imZg8N4efMmQqEJnUN0psiRMPNfQXJBSMX08iuACaCcmVt5c9CPEhqa
Jdt9xC2iHXhqfXEk3s73j0/mT2Trw7IX6xH1K3SntWARyZKjM7hc84syvN2spLpg9UvmGlQax2bq
ottsO4kOBGaK3D0mgDCWacMK8/2Pr7ORz7bLxochCog1iz+A+TnXZIlEDkQ8BBh5CEai9JEMhxXe
P92IuLGD4eMSPCFKG44pxmYyME8GAqmjnJjVP2rvBAcHj3XInFVcohtBHFO/oiahfKixZNVl6e+Q
39u/xjm036i/ICVq6ac74DEdXMiXoP2fQ0mstR0aTFocJgLyRVpzlFnBBvv6porzZdbD8++x6Trb
gDo/+tqBdvfwBD9yOh5JHom4DLdQsvfUJD1ppGEFs3sLD9LnmDVinqmLc7gfMxhFahflU5zkDE4j
RthzFB0MHYb56/bfxppTHXPidBYRcDkJbdrS9WTEhWfZe2fm/tXwCBEe1yaTErAbC8SlJH7NRomG
ruEtuCHGB5/AvmUPhAsnB95OpByrwvgNEvNn0Jg9FmxOojr9BO8h/eJH3JGa+ryM518C2poyimzc
IrHPcVbXYttIrXf697NB16c5ZE9eW7LXipkRQ6PDwXqZd3+0YxA0FhZO7lOqGQ9Pdm4+kcrWTtJN
pKVmmou5v55Bw4VDA0rXvSL/yUuDCe/B3ts7ozppApOET9XWSvqCEjP3LnrW8Bo7/L2aVmlf2jRC
lBAYsx/oLHWJ4bV6KmYO48gLFw3/wxkcZtt3jNl0DvtsSfSjAomBfbva3WKnBWI/Y1Evb2mH/Kx+
U4vRAWOVwI2HItfsbDjp0Qgyw59gW+ELxAhRQF+hJsQHi0pwls+05+ux1NzOW10ZNDyh96G0XxJk
l0drpLK1/YGbZCyfM2R7WwYP28pExp4OkkbLp2T+LWhxGpEc07pN0AKP9clxAR2oyxzizX9CTZxu
/Zcq7Qi5HvimNPp4kxR9Fsi4ElkYVOWVHr/Kd9RXoel4PgdelB6EjKOGKS+JTG4xNT7EApriw8+c
81XrR/23hWlhIDG80qcC3MmFqcJK1B4wN+SZpI08vaDU5jS9jRZpqfU0QLSgPILxkGJ7cxQ8/ZpW
yf7onDp45ZQ1gOHcBxUibNgdpJ++Q6NacrfQEuRBYwradqKiWzsYVWjW3a+89tcXvZ8ZdseE6N2j
fui6sNGMNaeeXys4ZD9Ma6oRjVfNWbNGuFMIMxZaL1DC1XrT7CBAj873KY6eT2mD3O3Zf1bc3ypL
gCFhAS9bVGRAgD4rxz2omCF0lPue38ZzVk0Q5z+0vxSZ+cxhU2Tq5ZzQ8pmNJ6ks64NLQwItEj9d
nG8Qx/TtBr0TYmbaBR4yQ9aoFBZ01vsebIKi13MV45xw0nwbDdVeC1erALVHARE0IlC/KxpSTD5X
6AXq6CMV96Fpp1eU1L31GqAbFjnCKyg3TPXOql1NfK2xtGOKG6rFntiQo1k1tUS4ZnKW21dCLkoK
wrqVHWnsqh2rSBkP6m26ITEw6u/wVDTGZrCGq31KzDnfN8eI8aOU7I1wmRDxpA3luuE3EAUwzZzJ
22C1VNa91+tnspPV1JNFtbJn3a+irbqEy6rXw386OEZkAJBLRpXBC0gniIWWBwM5otAOHkH/m7p7
oHPAB+yl5qEK/pH/gS/Iy0Ehc5zR8nBb9gsFKwRuw89YtxV/MuJ6ITZYUiakWXCaj67TCqsmEBX2
Yp6WnGZhrZadNwdZBgWOz1WB1gubcaN85fwLaLbTThDEw0cJtFVdkxVnoiFPlnPKXsQJjwzbHshA
eBzufGOREuW3nZwqginnMaM416MEAYxXzN0AfFurVFZ04M/YGsHIQdgrHfw2x+BEfP7aHRczBbtS
bEYZlx7WLFZvmQKA2lab7aWSIKwVR8hbZ99AWCEe5ZhwHUI+pfHThUz/cnJVZIHPrs7Lxv/wg8ST
aT2Q4fdZJ4yjyLi0StwGzEnXBU1JNsSCZvkJt0dQsBo91+jJdTfa0nGE43yhEDBIsSG6rA0TIR4n
zXJPe0nsLeZ6eLiCpOQ4Fw67XcN4D7G/HcoFBZEOaD2GVjsoXtSNWNRO8EGMfgmlmkB0vn3Sl6u+
VBSfwGIB3VusYJYsajHF4s8TrDu1iMoSdleXGwPzv3o7t26wucdweShkO8j4K7SQku38nOzyTGyV
tjztvDKQUTK2mA7W7CknKDMp/Ju1aQUIR/wOsoNMN33fmmCP4Ed4c5erA7srViLiARrDGnYqKC4p
WcIc4LZM2i1hZ6WkR5pNG2Mjn2a8q436C5Ff5Xm+K71RCCZ75X+23DNT/uHbv8ihHD3/kF74hinK
j0WHESiwHOIuCCyhCG7y2IjRaVi1WPT/W3HTv6pq1hpdlRBL88CQmxnGPELjWByf9plBEU00JbKn
a0lmVEOtuWuiAmu5l4YKGuiEKDOb9+bSyHXpiBOV75+8iTmwCkGUMpqLOOU2kR7h36BqNr4ytIS0
FPpw19DWLisfECqlNhSyDMYJqHvP+FFL2/or4fcnZft0HJIOkCUGhrt0oXjSxhaUSBkQhfRPvOTY
K4dgjai0wYbnN/IL+vnBJdt3KQYNJi2g4mwSGX2S1cDE3XHg5LKLISKq/5DhSsCn8YpyzJVmqjyy
VKP0VBfX0+/8nzdLpS/niLeXizdguCCZz1Mt1XBq4XhYswJcrbni4tnhTwMQ54b7Ha83RVkQdwnj
iT8Lk1GmrA6/raOjHNxohT38Q5hGoEDeRv9NKWbPlvX4TF7+2i5jn92KaAlQ6ovMvUUiz5/gVNz9
A3GKVLYBn6jXfG2+Vfr5b/DrxnK6eU+QJxesS74TI+Hty40SF6SBNqrRCWfO6x8v1q+8rSo12bmE
T6cSUPiDIhmrFReewBzhCG1YnzHdZooITK/IW/RpvAn50fO+wJUuN49x4PBX4XxDIE6vM1RcN3Ht
R1gDrrh3yjvzApK1kuhf3DSSea2Cfkq94454E6IupaRQqST/56DZwRQxbGcbo90XQ/ve4RbXUTi7
c/FfGMZO3cgtgo387p3DvmiEmkpg+dRRJMQ9kBRo9XevOxAsvf2ivI4qshUQcAWKPgLy2fEaOKxh
ZiRNebpoeazCFMxWQ12DgojRqIMvwFOh1D6y+Il8PG3U9cmVM1vUTLhjftHXMm+OY55sZA1Ft0pm
w7esngVOrZ3RL5g1yJ8DGQ/mAnELzSQv8aUnswwYVu4la6W5sqHEDJmnvUBWfJeF/vP3xfkJur/6
TFO6goH9GCgxaNSZxkdDKfMEPa0iUm8uzohmS6JvUtCXsGFzQuiv3JBLMuoyd6mLV9wU6SIpeBMN
v/zg9ZW6CfmsuX8bkybwlERJfE5folmfSH8Zb3j1Oj7gvrGx+8gSo4BERr0nOwrOzDJI7wxs6YtL
w4DJLyfaIVCtmhFQ/Pyvp99WHK7xFT3op5EoiRM3JFjOL5kRZHsKFYuAIgycM9Gjg5RQ9hwR0/yD
+dvZkbiNY2UETnjsT0JtsKRWcrD6V9LCVLkB7QQ4o5cFHc5BKLezqCH5ih2BG+D+dmUQVszDCLZ+
NDDNPSl8IwV6sjhl/q203oGbVl/2Ghyfxg7/PrrMMAFUAzPKruhwcz+4710qxJ+qaNlNJMp34i/U
/5u6xZ/UPaKUX61GWeF2XVB7ndPf8l769moEP6SVHRwq1k7X2w1VxIQ7LBSqvWVS+XnCLwW64SIZ
gidwAxXVyUSDJDQSQMljM52/IQTKPgfbbfWHYGpbq4LITYruGiK5ih3iFJ4C8m521431YVPgXrRz
BPWBYz3uzIy7FT93RB1jFxe4Eh6YXEYOn6WGDgm+xvGqdwRgw20wV9mNcWrmYLNoBu8p1a1XWGfv
byHpMyx5MxJoUX4MKo6GVSmQYrJOW0JMFExQK8CStf2Fmk/MXeFl+nkYN22uc/lfFlpSLqmoT+SK
fFx7l7JEmj9pBX7ZAoMV4eX4CBC4NL1mGc6el84G5BJOy9mX9743ptJ90CYw7d8x1kUam9vjlqEn
9MZWGvvbZxKYUnpF50ixQlZqRSGARNFJIHU/lo3bj9dCmH1nqVoTUj+NU/IVLJn7CW74xIgCLS3y
VuEmX3lYt51LkEyshaE8u3QNO4pU+LnNB3xvJ3ufOQmTq38JGElmoDVTYi/Onwz5w/9YiCLi+DD/
VC8IGU+cK8G5kYk/01BJJh9twvmZzzO+Fy2v86baflgKWqsn0HY7hqvUlddq5TO2SC7rXvHR0c8i
e35anP0hbTLXaEBXqXuGT2acsCfzJ5RSBGEyxKVp71UdARF6OhYmZXp4/vUA5zXjpy001uImJ+SO
reSSAJjOc9V2qJ+Cf2u/b6zF8FgIDepyUcn5WnejSoeU9ZEcPBCDmWYgaKITWeiXpsntmi+/WO0G
kupxB07kBJcUHW2ICuaENO60DCK9ywguqeqJTUqc7zBZ+BtpneQSpCzrzGLwdlo9puU2fUxEZ+at
dV2YlOHFjF4ht1ArcRkyh0UA19VEym9pnYYUdg34Q6qlCj4KKIUiJIteS7P/HPyueMDhUO4GC5IS
0fgMPBkPPXJlnnSJ1LPCtoLUSrELma+2mncZKcXwub8bOkrN3H/XCfOV4rYuOh/ApaZZ9B/XcWTm
NjOk6wqkT5h4c15+MvDqpDPDl9hxPfFXRSTq+IqdgXi6y1i/1q6gTPqYI1eE5VW3wS453kTUarrk
28UltFjZZ4babSuCEBT/qIppV01vtKDq3rqZGpXNOFeDaCKR3+ksRC/JZbqkPqH2sObHl6iecFM9
JqySzzDVwA87oQlNMXjKaLWS5W37N2IcR9QIC5pqFWv68laer6RXoFRqEnDIoTF5L8BN/pwWszZ3
DhJf7THcDyKE4MOV8xaaOAiT1S6r3ia/R7qep7xdBsgk6UYL9inEWX7N5oYn+ND1NQig+xUkwoTC
AWxRJJi7X+mExdCZ71TiY9IYgbnecLR+W561HErBznpJwRTn4MhepLRlyqvhXdGumPk4AEhrAgDJ
rsES1ZJivkjAKS3Qr7a0oUNZtTRmc+/az+UkV3BcFkuDJbnYGb6AELfot4HFDChavoCNsj74AqAP
XnjidWDRoJdPSRFpchBnK+x+Z2AB4rN9lsdmWVF2bkDcCvvp1sbZFkTKkorIbbzGf05AVRwylpZF
iOK93RW4974PAfzfhXAtjLB2x2Brl6MCAOIp5d0UzFMP4eLEIWhjEdlBOP03cXZEzZLENDcMMZG7
TbmceKnOmtBn9PEpuMQVhMMHT1ixCBnmoTDoXlJ0KHv+Dascaux8MOMrS2LOwaKVDu7dXMQK9YWr
/5YCfTsQxhfUQeYsMHPznnMcbAXLWnNPcJotGBciHx2Ni5/vPorNqgaVJDL3U1tVwL7HY6NxTrUy
hYxz04x91ZFY4O+uMDzqfaBDm8JOYVI/N5zf4EGBITxIMJmWh/s1iiU/htgmDU30xVY6GjaImu0r
bArJUMBIesovXPwU0LX/694P87wxm+hv7OiBkX3cQiNbdgUB0UMrVBu/5CJgiZPWlm4jUqaMZQsF
opVaXinfbDQOtgs4no9uMnVHG8x07EKzEj/0ZEe1yJNjo9/G57dTpKANaMqkmgjUy/hOk4Kkz377
vUC+CmqiT25gW5TsmnLOKhznG2UBKAfdzqJDA+Vjyor64fzipDszmXIJ3ZG6M7FZvplWe9aiDfUy
ttunUJ8mhI37DUx4UAtKaVZhNTVECdvyHmjHGEadBcoy+R+3W0lY6TTnZu7mP0JWszvysJkGTK8c
ZNs8sT5w9LIInFJPtTDOCmFUNcgZ1zh9SrIPFYfRWDyKu54JEBFgsRoOuFgyngZnI2TLohpsMhSJ
tOQ4P4eHLm74DtVE2YoNCZH/y3uIhSSa2bwZblaO93tlqTykm8wB95ZPhbjb6rTekSA47wAVBTTQ
DNlzazt95R6s1vs8sUnSHFnxxVEU0+kNbR6jSoN1yCHPfNxUjUgzvHLspAJDzk1Z+vqqOe21e1nr
+NXvOWojOiRu+6ljlWlDtsahx+x2BiMAfeE9PrUpVo9n69BWhTzQDguf2Yq9gTB9eAujf00cfVIZ
F45A2uGEs8HJg3DBnJb/Hmj3WmRnUTu5rjX8qMYpUCbrOOhPSYqQYCPmSgI91s96s322N5mWWN7L
Wk34FMIFZJJC98YvttaPgE1fJfOx8SsulXamt2ksnxgrm0S5+WL8Ama/n5j84X7tTlTHA0T+ugJ7
AlUjJ3srvwsNuqDAqqlNCKyLRaITcGMQRJfLc31D1O6E9TTB0DTDAWO0jzcjdcJSXnGK3joPTmI4
3OeOYTvTs6CH9GYGgfWfUYPQY2BmxvrFJ0DvmNXH6fk6eljpQ7+yt4FUv1L5/Y3WmJHpymm09/69
lcjlN1YrAG0C6ef87iWkhcTCkwqXwk4fNYKJLMa1OkvaIg5DycuoYVgPxzzMJHqVKqR/9WFQxcDB
IXYcWTjq/ghg6wecoN6NKVfv0aqQXEJB8JQ601OC5nxYxlY7IFT51kp7itIfal/I1xoVFr8vE/if
v+WYLQM+iPL560pvuyrhEeoPMhINermzHFP69lhbT1Xvi3zqSt9USng60L9D3hupa4f5W6UE9DTa
5+PhsdvBFVyY6hkHcoDZCwS15Lg/wG0uM2TuqLXLfIRBMKSRsGbKGmicC3ynhhK92zf9ZEqS70pM
RAFAvHkxT6aJGGwbu6mvVDaxhX3A4oD2O6t8jVqttpIcoSFX3gXyzMGCKwt/vXrwoOJpSrd2BVCs
j41XZxj9B3O8lYTGcbUjazHQoycxtqslsVWLJ0InwkBmIxHPVWrv7Xu07actNU5rISi8pxHzdOqs
eVSMzyalnT7kYnr9UrgDTKC32wqgvWgfTNpoq2Ty9tGnvb+MWcl3RiKj2LG0OXx6YG/yX7DbYiYE
lfQVO/pcExBnVhuhu33wUKLpJ2WXIORq5nencI/DY0LNiSuUSjGU+/ogVHCecqPp+KzJwLIsh6/I
agTzPzSmBkrFF1HV0E7OrlL0otPpNlcgWYcyIFFQ2yppD+nwNe4dh0nqudKf6z/dvZRJLCyIfzFW
iA1K/SY+IDgo/RnXpyTpSgPk+P587jJI7Y5Ynrz4oiU/NKuaElvTTSmFzRFKwt4CbNiQSPTOqLiy
PhxdJM0tIaHwA7gjuF1dhZeKW7zfwuazDmffOay2lGt5BLnQUKOqx517+H09mKD/Sxx5FPpOqigR
Lx7t2Bv6JBeRwH3kgXsyYShj4xoeGHD0LZ7G84MZOx14SQ56GFBl61FE84vWnm539ehU49EAk4XY
vQiOT3FRiKOR9/O+ztyRbGal0S0IOsABT9kpoRnWJHSZ01Pl+mYH2jXbZD4Myf9S0jL9MLFUEQqm
CWQbzp54nigc1lJRckhjLdOVl61FxIJ0YhU8TR6ykcyoJYqTytJIv8c61+bTVZe+Q3J2aHNwpcto
3ApxRpFFuyxAwi3ilpG7n3rxojBgzqC487VkmjVQxbctI0H9sS1FuR9+i0NlbzxAwujjKTjEQeee
pO07qGYTgeKuuEnxmmhMd/v6tAe8Mdb54T4u53UCBNwwwXwxsfV5hc9GCYEuRuhGYNRQ9HkwxDSl
Tu9582miRj8wWwl4TjqkcL4fscV35wFB2na9TJW7kLAykZydRHFXMsGnBP3Z55rlQaJDhkHRZzQb
CELO/NGhWk1S9ZAgJqLKCLIqliVmJ0NHnUJAK8wtr0+buBIAg4Vk+M84H/lw4sQAF/Ql29rWpeXa
5bhlvVHv2sq6OhXB3e4B2sHTPP8UvSPxqrT0rQSysZZGVKjjrCWU0EmJRPg52w1o4NMiz8jUVL4b
UT0gQumr5Iy6/ItP3ic/naVQghYzGAqfF5AS6SxLmHQmblJcaYmcQ5s7jCwrUlhwdKvgZIPej+71
2jaDoBz5DhofD0wqnw84OeeYVuhEfiyAJbVOV3BsnhEdnkCQ3VygUnXfGjjiKq30te67sO9AFFZc
TgOiD1u8SGxWLE37WnVpNWfB0bZ6rKckE2kHNHfY0nUIWDM3UigxmzfhAve18ZuaWhEwbSL8M5yN
Czu3wSW0Swp1JATB96Q+ATXJKSq1vG6/E+a0xJukfNJuuXJSRFsq1fbAH8lPR0EkzdyH2+r7LSVv
Z7SrhE0JbTGPNzCO8TXzGdAFKRsueqtrxmKMyd8klBzbduVlTMiejsiZGE6J2Iqj//c43lP3KDyS
aAHvSRw74lS00Qw1fnFeWgz4EFtleGjyunlpRHR0Y461cxQHn+m8Ef57CLryadDDi4n7DAlUDZBN
s+wnnHo1xC2bK+IDnD65xm44vRhi6BCCTTH2mRdW4U4X/+pcbJRglcF+EjzpXCXdZWZrAyjDKhQR
1NIfktruBzSBXYZxiIedrBjk+ZllPHC4cJIPVo034GWjVMepeoojaqNMUyr5HtibkW678FLxn+oj
xT40fLmw2SK0yMWGfWSmdSmve4kymcbindqMp2A1ijAnIvoqUZBg3rlwCUoZVsreAkeO+XO4X0PW
VxNGe2kyW3lrfNOo4QvnMWCMHM24x3CXGL6NOQWmwne+SyJpTjrpxwzpcxXUvN52s00V+4KphSoU
g5eUgQcmY6ZYG9kMPhQN5qjJDyRQvU0/B5rZJT6Ng/mr9l9ht6cxuofFB6EBR9hhQA9+GSWeDbrc
rADYCGxKqomn7tjh0KDpQvjuMgXCGgwBLXrEF7tEP21CPoYnBRc6tvFSnAWF9mJOtYCJrRV+9MvC
FXPN6XFzbfwiBGDS8MmILJTQu8d9KzGQYU+ogCjOlRqBScHmVgw04w3dCBWwlNMJeA4WdEyeURnS
jxSpEQUCPCSi6hTtWmtq7V13ECplPJrXI3OezT7SRLl0BK25WFfYj/5nd5fIuofsQAuXuKwKDMBz
DCuZxLAHkl7VN57SluSR1emVZkvIdMWCj0cdUx7aP8pGoHZbMsN3QDlgT9YNSu1AyObaH/to6Ljw
SXLvFP6fzEO6HSS0SfzhXo5hHq2f4VFPsi15JzzlHMYbbj0VFhsxVgD85phaRFD8lOY7EXKi+VB3
v+jyipKc5VI2mYi3bs0eufbTf5fG0xZU7cHcz0uK9yNX5hr5Xoee7eo0RJW45RDgFzWjrU/Bu1oy
CztyCMcYsr0pH2nUZbegCZrLfG1A1AF2VEpwjQAeM5AA+6YyIt6soky3T9n+eOe1OyQwWGR0rm6+
yOfMo6sPyCW0OogGHTzGHIpXUR+zVwDGhqvYKQSG2U9EDSAOhRDHoshGRxD1wlW/gOtnR3Jhw2RL
+WZOxtOzd5ePTDy1piYuGwTTa+HI5loax8835y78A/frhmZUtEBxF2VWIT/IciMJzs9NH6az/kSQ
hZ/hPLkxOUfOMmuaqvN2l3DFWr2hWFUvMCcHkf3o6l4TRSVlG4t5szUMb0sKLkU46XL0v7I3qEXM
Xq3LK1X3EOxYzOYSNTFpyINDXm2PBnU2QA+iQxH3fkKqlbtVHFJuG0yF0OlvD/iwP37G0VYAdQwH
kELoJ4uekZD8tdj7RLL8JMbRd+M01lTscmOeYZmgyvmyi5wLEI4NHNU/2des7Z2j2f2KtpQR/YX5
kWfcHewc0LtRL9jzL8mG+SY7KT2dzmZeM+qCbMdXPFV7iBQbqE+RwvFQsaRseIT92A6/6MCIUO3T
OkZ3jLO0pSW7kcG5sD0Fhpj9E/7pu7jtAYAsAi6IWfAex6F7JVblDD0wKF575q2EtNxh4wg2KHgN
2kOehNvaTZ71tsuGSuwkBOxku6fkIlDXphblHhsptbtCrNhdFt+3hruACHucnpwYPlnwsUdK64i5
soguDjuMf4mbf4voW2S7Kj5+3rZi6dPLWIzCHMAJMed0kDmJtR7u+lWX9JsWJ5LqPJeKrsxYKgf+
qf1oOKwcvUmYalu8RpMn7AmIxz7fNn8OrvOHwOyvW1V3E/9tL/a0cS9l7064xANBrLtiUXterXjB
i5xc31Ey7ioeRccIjVfA/nLaNdD699xGTamr1TA1s6ogySn5BEfHgfgDz2/KP9eIIVerP7m/vSTU
7sZNtJntdMdYDw5URrL48yQEX56mqurcTrgCge0IoAHY0htrs3jeyZgICA99tiU++yQKyaSXumJ2
jh8zp1xqQjArWCCp0KW92S678R6YS1Qw4u6MDUcDJYyBOdiyG1I1el9nUMA+uE5rPm3tR8HHSEx0
WIDR/1qSJR2ZBETYp6hPsvA6kznaH9954tqhyje2QDVqBLQd5aC0Bd/WNeKb7eJDrrUPMhed0+cl
DAhDSaSbn0KSnj5HhiS8zh9lWnunrI8eSkRmOI7WVkWIEq8WmZh2zVh/PTRLnoa3zGlsLCjSDwbx
VhpMdT4NGO9qlpk4W0haLiSnzEZXIokXAwkzJlgFZO18hpt7l/pz2X4KHPjqS+Iv4ptI6llEUVUd
jioVdK4eqU8mnrRnudA31q3ePU3E7JsQBHMhMRiMLGXRYQ+d8J6K+KjPOXheNUSdEcGTjGu4OnIY
/EHZRimT8fIDfHWGaqZFYC2WSswljAlO9Q2mwVlT6wuTyIf2tOeGRiz8AD+x6Ax9njOpOoFQgxT2
nh+bYM9aLXnLjXXB2l6PwFn8xpKFR/UOnYMU51WNFR+0rtZtKlNzwuzZiXEDzB493cEldT38f3i4
nN/N1PhMJCVjbICOQCpWhB6dvF4fmEgtAy50tlZcmC91K/fnlwXatJDs7DaZDJrhZYv4pzn8+Jaf
s8sc9A/JwTS6agpG88vtCGIQLjaLDh1qwCqGhyRG1iSGgt8ptrzH9Hl0HdT3oLrCfOjmNKthSIyA
xUbJxmZxySS+eeYr70zBG0sJWMZyDmDC19bQW3jdMBHenhxjbHzCFZ/caC4xFBVw7QDT+gCG5g/B
uTXHRtNz7crFKIOIPHWUetwxSKMtcK0TMSlabd6GTd513b/Fjm1G3QUpr+Hq08moi64F6cL6lWQi
jL7gfkagpkwNROUIIVisq1b8fQ8N5aGvsELn27KPfxkFW/TvHJWtHr+C//lZ34kPX5ZhGIjndNzc
iAAbq4CtflpU4zUOivXNXnL1+uLwvj+j/ka70v08az2H+0HWFAFxFW9m8bpB66s1L9UO4cfawJpv
z9FsPd5ELJSHPjGi1jrP3NAvVm5S170aXjIWKmqT3uWUTSQXxMUNR7faM3SGkFu7gRB5su/TweRQ
ROVeVt9YdMVZ/N4/NFlEiA/Pw2c0MXnIjHiN8Eg7IaRLNXCpmxMyRuF71nfWlI0ZpMyVGNGvGon9
Ul+SsLVw8oTpSyrI90AQLQ6iMLVa1+Y2v3v1Vsq7mGnD6m8FSlNiSv5pjCo/1aiJeUxikkS8MQ+8
3bKEq2H4w9qFR0lrpFu9ctna+q6+RIYtSd8MhgYSy8+F6YG6BYhNVilkXIZf6prm0KFL4e/bEpbP
Vf47m+y5sNK0QwYGV3+YkY7O5HWKhQ4V/uUcXtrHW/Ia0cnRZ7vZ3ShJLXaBR1ylcLlBBdcndy3q
3F3c7UvGP1rWGcPLgAsTWdM5l+ls90J0XgcMuiSDbyMr8usQKxmR1iFox5qnzQJJ8KvtLbUjbNBI
jvEF1OJm6ZGkWq235GJN/Lr71dr1NFxU2Iw4liPy37ZLf6K2lsMIq1RmkHFZkTos5FbYRrLsHxu7
OeH3LiRnplq1LJ5HNXHs3KuLmt9FQw/SXGiShiHCwU66u6a+DiAcOWTXd0Rk/GhtQxf/AmVuPEgW
vfioIKIx/Tl8P2z+wl9StBEitQUJ3D96A7NuNRhIonAPtEYmA34xDNL0nK+Nl+fP8L8KRdMngL9g
NzPO4OVQB1KFYZxl6dmbsFk6q2RlWvqFqX6nHXSjzY2x6VVKYdjyuFvBgOGcjTjf65KGxyfqTtmI
x48sF6ARPxaq9/SCDQ24qjf7npDJxj97UuWi9PWaXUWf9G04GTFVjHkye1VTiMQzNHjI5secGJw+
jVYLvFYtrpd6Rv1jB6jpFU5L8LwF09prUyl2z/Igbv7t6fUYDi8vhD5ac8MLy5CEghmgA2WDaTlO
o6UDIPjh7JalyKAq8dof9n9cPh8Qo9yjmbnU2EoSSDBSVSqYfTx7R7ZyrJTlNRYf8YT7x0MeiquK
uyhfXrzKd5HjdTEiSNWkJkvtY9nLi5Q8z8JveJYCRz6bqaTHKMFhMweW1gBroPJ83sTbWGcwtrxq
Fo+1CoJQWbTiS/HDIRpCwRffe7JZLLl3NJMMSKHblvlQH4TqWjrJ5PqAPLCG7fMAQEfu2Ybn3lfo
Gx64w7L9pjwxMF+o4+yQRPXYJgr1QdfqfT0anIF3PB3vzxD5qwvDa3ROcXZ5luH3neqj9JDACezp
n9OZtLhhlIyjTqvWrFbHFzON4Ln6pR3xMR0jGINbIz2fnVyQYvpiQVX3VfuawKHUsF2FOyogcwpl
Hvkzr5/XimARJv7ZHuQr5WLuUnidfmq9od183YwJ0Q9Xz5jUv3X/Hxt9xQeG889/TLWV1aZVjNOs
q50FtbQ64tinnY0UGCkFYJoZpxIfN3yplKzT0MEk5JiKRThGrjH8OhaMXqTMy09MxpHAdGyheRH6
bHwyYsIibK/ro1Nf4OG6kC3LkQPOSPn/KVy5+yDeXYtop9OUyIUY8H8AZJYuTjIODtKtDGDYibJQ
JT9416cBE/D6MbYxb8u6l+XjdB5sg6lgsTZE7j5zV8fwD5+DK7Or6vyb9T8J2eyHXIRq4tMwkhkj
wuGJvIhbHgpatbEKrKy5cRCouTyCC6N4c6k/TvxZ6ask2ItlEhJ3GvKPRIl+eQd0UPVvIKAO9/T4
YVhRrZGsROpETJMY/dxgQzY0UR00SUJBSHWhjeg7+4PFV6CW9EEJWHynNz5h/i6BTBIRYUn1b1St
6pHJnz0vX1HJqf3l+BSlOz445Eyq9/+G8RRA9MjpTCkn2jadQp1QKsoxN6v6TG0i5Z1dch8doXea
cMa7nP8/mjHvu5/lnGKRQtF+nRdF94hE7MJUxFldsl6/ZIDneoDLPTZf4bLfhXb7rKPGji9SNmqx
UxaKbkBm17usgbT99qr/9WwVhAUhrr6d5DXsNmUmQExbkM5DcaLifoJcPXQRSssIGEuMkE7KXCTK
omv+spJ0mKjNggsJskmrCGwCuFe4qRl6o/5JCC0tEIMRtaHe7qNC5+s3hZjuY9odnKEXA8YDNk2A
5cip1kxP0tLnqqRJhwLaH5fodRaytrl/1JIyhEv8eiZPHmdYyaiLAid3Eqgtn9aBFJV6rDXP7ugt
/g5R8OGQB9FnhMKEWPSc54PNr5DEy0KPdKnjXeYq2JGqi14qafhkxPEgMBrWzGwJoLTVhSMaYk53
PVmj5MBU/OFWDlEh+Y8TbgGEyYnFg0agO9YYaqWtOD8vbZatJ8pAssTsxOUa96oJ7938JWlW6ZjZ
Xv973gdUk5RRbARuYngHRmydjnF7mxVVMsKGfKEChkS8F3SpUumfPToGMOQh73nAad8kmEG4nPVd
a3apesSAlPpyEGcf5MW6AzdJZyKrx4VAf4xuTrtZ2szEFTPqF9ajGKBw4hMN1t6wd4sPEQ4BgdCD
sfD2iHlEWpz3knalD3ES/3ygHN+NYp1H9ItCGR0QaMzFPGFUfsak2vLwy8tNKZr7MHqenOJAZjOF
LOIOi5E4gr8BnSmqgUtgBlgGC8y/0QBQ/sb8To4Ki4qKFiXZ1hThhNZnD3bsNQiPB5yOmqikVkHc
DzhMwkOl4ESEMWaleQQrFZGm0cEdrJPvZ3zLv/IK2Mgu6Ojsf1jWPnNGxp4xidtx9uy6GIHtLuyp
YyJtXTfeK8tXbOCVOlSDE3+n7YcDRnAyhMopPjn7hmNlUZ8lPhVIujV/YssG/H/Ci50UBFvu+BdV
upWGScleMF1rZaMziQk2l24ZmaH3h+vwAX9PrifwuIKWObjJWG2f+m5h9d7vrhw3rotUZ5OBBKvC
Z46zouRxsApYaEsn+ktM8vf/BvzfKRtW+nI7dYfn9BRe6pCg4ywZ9JEFkhTlpTPZ9AfWuTNklYeZ
ATXWNPbUf/cKXEyRm8vpJL15G88ZUxLoMIB9WFNnswV4MrhK95LSfBImTxov2i9yIVdhhyD6XKrr
bnqNCqT/jc+hBFWcb3jQC4ce73PahOW+Z5EyTGcGn/7sdagpD8rE590nKqmOvF6A9E4u1Hp3x5N2
MDhGUUVLXQPa6km6P9h7zDQldqz7hr5HtM6wXhsxno2bp9ZvrwhlpGfPh3kfJVIkhNA541gusGKw
yW6GIvvcOM0zR/SiZIwADUOL23DU51cm1VkPMbuFoc/pFQFleiFBUmktr1WjcgvVZQUQd4XQOuve
/oblyHP1UmlxUW0/MZWS8GHlsZ+EpcnnTms+colPjejxqlu5daW/zE5ZYJwX3U3CniPSFjCHryRc
Gz2fwPkqDSy0hE+YDOJJdK80AiywGgggvG91CgjLwGVlPzp8VsNccsUjnr85Os3jUdmaQc1TmHMi
xVPk5JnRhDV/LJLOrT8TcdTx+UHMUu5/TZVzBQ59ammk5OtobhkPRa7SmV2LhTYGb/gJNW+28Sly
koaCheryDZLoOSZ50GLp+tl9K0MVcjhsdFoFB2GAFi7FeCw6uN+lugS991QlyVmRVNaF/ksmnT5g
aDHpXD9j7vSWTFPRM8nby8qHXHEErgJlh8hCYkx8H1+oaYAVRNFnCY2NiWvO+5kkZVASF2UOErm2
91dIkx8A9vIr2n9VXjpBY6vceYERbp37oD9tINU9j7Vz0NDBCkwtPoYNfrByNr8QqhmWYJYa6FSn
8qycgIxRlXQq72VicujXzpM9aWQOdMgR0CS07IIq/nvpRWYdSjlZKptpSNdbSDhmXoLXJ6Y2xqWI
UZj4sm39HqwHM4b698TiyIhgrvhSyhWOopbgB5goBuGAeEervxfN5Rj5yczH0nlWh2MSCGdvw05c
fEna2s5Q1voLHNyg8k2J4ZTnp9neTce1+A2AF+059p3LnGXjuEm/ct92B+xEQpQNFD5kIJmQXM12
jVeDlgv4gB0BJYnagQfpCTOrW9rCURXH5PmwlCRrbEOskFUOijeFbsmaf/g7i7GethM92BbyngJS
ga/uzNIwFhZJm3EftYKld9lln+ydkjmG05BmZC03QfbB92nuUUGJq/0lZWIsx+ZH2Hvf4vixQZNd
CqU/D9aOBX4V8qx/p5wWzh+qZ1P9ptlQHR1qgqjtTVN3AgyqzmRW7ve67SZ31QvVEMhqutkrDguA
N0Ij9hmxJqo3cKkAwPyeZvDRxBw4GqS0SJMbgi3oA1LMIeTREYG3ZnOrZT15REhTaiQLrtqcNdU2
MeEstJ0v9Y/yhaTkSnfAA8ru0WnsYHzNzO2HLXnNSHvPrIRAoYvgg3a9WL43GUC+md70Mfiz5VIf
teqtZRQIsRBFIOlLgE/PzccuOcz1A45P7qaMD7SZtOivVQ8KoXOs8g3fgIyKtgmh6/GpMEa/EQ2h
Ybk8UXSrlaJHS53NlyEbYxyGvjxdnjGcKt7Vb4YukDjiuRaPQ/Lka/uSUgwwfRq/gyVMCI6MLcjx
CTc9LshM50QJdRldm2IxikrXzIqoRZXPg77qQtFEEOlmWYJplMR15LaFcCfcbT4V1Ur2Tju6J5aR
h+pXPLXiI4uQRtQ8cibOtorm9y463Muz3iKLR8VoFgEcOm4S2Ca5XxsalLflY5pj5Gvcfq02jr3n
fDbIfiJryGcVOG5ZlLcw4ivvH3CdKM+KJImws9YGnsBG1f7rQJ3NBeW0QPKDLdog7+K/BF+zSfCC
Mh/f6ZUu1DErDf/RRip37au7mdlkHf579bIUEx6zfgJFjTwkJrUxR70eKf9P8Pl1N38ZV9opCHm2
6gqNPZ9nCfQJlAe1n0PeHRSZUhWwWfIB74uNxqNiOf7dKEOIir4ArMSUGXYM8wtgl+dBBJGH8j4K
408r+niEqmUpXruv/4GgS6wTzAe6NGxRiRQu80MZ3E8pkOrl97EGPYAowr/H25iPtJe0gbVCYQan
aBG1pB96TTsJw4kL+vB0nkXXshM4L5v++Y60B6v116dw27EqurMofNzGV+anY9UDXskCdyLBPqB+
4f6nmDTmFdJho07RAl6Ax91ouTT58WqlYeKbHaNkXVNKKo46hRukVfFuY7dR5ZAHQ41NQy5uFaUp
QEVsCCYXVWJHkp9PUYJCOmCrYQXz220iziMQlmC6dZN7BhEHLvofnVLhjnX3uNOelLii7Vg93Z7Q
qFQRq/Oj0IEEWhkEersbKTK7Z3N8QsaApzZHXwD+5CI2fNmqYDUUgQ4mmp+rfothnQWm+5K8AIwk
fBP48UGMld+I8zHxcwEqdoE8D6MbR/vK5U3Rnx+f7zLHmw4SpkfTS8SYnxMPCIkKWo2wNGOxPAKr
+DD4G+riCMPUunslr15X/8rN5u6bkRipcOqEKj9I5mf00vRiVtSUFw7rI7sPzvu3kuYbMagjnfuO
OF/F1pvWg206pCHE0figsZ938jan87Hz6GsFLB5Ql2wHnp2OhMaEgkuWE4Zl+F3Eil0dblWWvqib
/1L2Ocr2rFG6J/Xse7OHsJ0305mejEyBjqiqPhPorEuiG6Ojy7tpFBeECWXMUEdkI6TqyLBj3K3O
BpMJwTepeBX94RNZMAvqRCrzqGZwJqaOIF0TYZvK2CdokLf8wg+08AVWLDhVytqn/QLbPsASwaJe
vVAs20DKk4FsiXkj0F5fpDW3GiII09jQa4C/JbDiYkEBkYD5tLmUOG+nhxOyx3VNAY91SeK2okQP
2woKMtPXRK6Aub1SK0hcZm2HwidSTYL8N5uRIU6M7TwgVB6tCiG1tACAmNEeACMdkX9sv7hahDCg
GSR2gJ4l/hGVzauCLE56dIpd1WjmbEV2e7kddK+89jAQSgwQNJLapu27LxpdfMcjG+8r7pALBFXV
tq6kaMonDna+1uliVVSZk8qPmTwsG6nqr621xdgdGOWtyUs55xUpMPgZWh4yNGKRSS/NsFPjGDHq
l5lXvJcgYJW43KxgNmMLy1oUGeoqffZFiltBvXQlZ9Zi1Uoy9W2pOXYWgPU4O4V1QYfcMOTgmP4X
IzOcrRZdlW39RrhltGut8ZUjqgmabWBD8GKyWE9Y/f3BHFtXzgzarFdyVF4C6M8xGgNoDnqr/TrE
7VUzDlHNTjmiGsN7NT3uwpquaDXb8NBPZ59og0JPaX1nZkjxj7isguL6rnhBqsG6SSZW9pOSjnSy
3fswvoh5ofZLRIkrnUEQAvYVRs85+0+4Pz0v82Eqh+xtrENST1Ov+QJ48mdjgB9kgnTVgbVlsKgD
vnejR2aoLPHPmAm7wNx94oWhBJcYQ60Cw2o03I8JrWh/we+aWE9+vGwte/lP4IxIjspWXJRwOLxr
XNHvyfP7ew7IwDIW5q5KGJrh85jiIPzFXZziTCZLwb1+nTn8UaIu5PY7bUc7Kd49MDvsE/HwXAnk
wYHJweZqUn+YkhovbhzhlWgROpp4eQpZbRwywVhCc22Bn6LvG0ZxltPoN+KTTpHdv47OSWeORsv6
TVAkTHnFjPBmPMBoXbOZzlAvJhTxRmLuuu3j7VoJQcKELWBgb6rKBSVz2c39je0OjpKUNj6Xqc5M
ChpvfNaVvNQQr1SFotOZJyivU89ikiAaD+uH7LASfGWr3pSJa64NvncJMLtkU6kIWi7AV4dmluIY
Jy19rbkeQaAWJbHFDupp4FI1WR6gvbbD3dHf8V8aC/zO3ugpZcG5JDBSjdpDgzn0JiworK5iPW2g
w5cN19reahFfIe4KzB+LaHHA4WG13Q1rLo8LJ2KUbB3SSKH+VkKo3TpgQ6VNk++9Y7gFIqLmXB2h
b4RLVdX5lYLXClkd3rApsF6qrTSNiY4oT681w4poo+dJb8TdrjagOsOk92BC7Bv8lfarxn5RjImK
beBHXwMHytGGRdPZurZnfZstVMFcIgwXnMkWY0OQUOIsQv+dPIkaWssoKv5SeXOSscEMD3wJIe5/
ucczJVg6RC8aOBgqUPlaRnSj+m3nNBmLTygcnwBXAjQWjkq+t+FgrjgN3B+yZHibLQqxFuFAf6/n
F8WvjkSyiDXKBLCky6ZetCODlliiQgT1L8EzxAz1rxzdGL//MRdJz+KZjd90yQs7QdMeesB20TLr
Ubl+Hmv448JjuASyGiFWMv3lgf2+O0nUUnMxnxsD8tM5XNz2kld1HKhHZf8JeA7iaNnXEN3PAqHM
iL5AlgyWkKtoxBcut/nykjX7iac/kXpHjeYkLiV5yYbwSu9ISI6gCO+zXHZROya8ltdZa9GF15c1
C4GnNA4TFx1ouMcGA5DsSBOk3hinBV/DeXMp8vDB4cPVVQzcIF3XEeBl0gvCbg+29cWn+F59NEoH
y3phaqVE97x7sUxUT9424afe/yCliDGC0BdNagiwKeUUBkfsWaodtCxQg3SC4FXMyjwlGKlb2GOk
Tvs/jU+y2uJbhHdatErPadg5aj6trxz5ewfxLLTGqRycJ1Pd9XwMAySFzB4UUwDxYgJ9Tfko3gOl
W2iJz2JgJDt+QAmhMaf/zSW9ryA2H6aiHxhxTbzy4thRhknTNQAfWmk4f8F2TRaZqwn8ijD8VK55
nV+MScnw6v6v7u68mXcTmnAGAjDwdc00Hhk8xxc8+LSPKk5ChtGmiJLhFvtYMAxExtHWvBpyow7Z
N1Rhf0rZ6zUjjdFcwf+K88cCoYeFXMpnoYTiWCsSitbfxkaIuYvs8rN6QL8MhC3FKjOo39Le7LXz
ePzcoUnhh8qyBe4+1G5TYx1keSJrY7SUYiZ97obI5RrVGZJYP0SIa4gYZZX7smy20Vny2eFo3SN2
3Rzz9V2UhIOFDmPN1EjrtXbTtw1e+zZ2WHybiQ1CiaEQRMR3TSo2DH8rXylQR239YztvIBT2QS1i
aXuCv6Z9PgHR0OEErL5bZXRc7+jdZy9byi2HQ4v/9jLXyVcFt8EbZoHVmJbmNtj8W7btj8fcl6kn
hgUr4W3ppQbMI1Ig8w+DE9J+cjm8of4O9aZ6F9aRMka2h9GIoOGmjCFZH3WeAtOuzUCcSwm4SV1w
8F6DAawwMLEj5NBZCzrQ8TnFmRPLHTTZMSm1A1JV2/tYNEPXw4QG7nK2MJcbR1wmIx7cz1YlXq15
gURigiRuJYpQ1YQfTC+4/GmYNzL+rolfV/sFEs8risr/J+OQ97oGpvdkk21UI9dVgLWsFjSxZ3nh
z2Wz40xFm+n4EzHYY9oF5q2ePZrYVb5Scjy8dF1746CDYDrpgjYaeurkM1Rq45dGM97hMz5oII5O
kAr5GdQSf7BET/XEOHCZJzWKDkqA879KqJEXgcxQI9RBEJJJ49tot4rPM7+uGuv8tt03KA5LTxku
fso4KErXRrwEDu9zIosQJ9FEOTvsDZlEAn9AFRGPHC0om0Bg40FxpeaLccVKYmKE88uex8XW8UYh
VhuptdoEQjku8O3jSKUisOnQSrWjlbBhMRq1nXyiS/vjhPgm2g4lIpYNDM7TDJpTD5XS4DRj+P44
RbZ3zWr9golRzUovE8IHkd2XV1NrVWVOpUcNWCtaU5avWUGthBT5DbwUwMDenI4LFt6Je72xdvFg
FnDM/KLTaxUqQSaVPdH+/ji0HRkgrMIIvwR9zALEWgUihx9UMYvJJ1wdoGb5kwIjqU/2KYF8cCUk
Omr4EZaWVcv1c9uTtv6kq7eZo6tgkP8m1e8vn+4KQPSfryZzvVdYyijFk7dfTYmwKSd4k06MlFgk
31ojZ8ly37/PRgEiRU+4+8BEJsxRoGBsTf76ZdkilAJPeo867WkY9aFLNGV8pI0lyskbBULRJKAx
mBD5MW0lSI6UBl7M6S/t50aY0beqHmLAXRFxE5j2d/vCuz49iLmqjWS/xmAoWGA++PHZ00S2Of/z
+H4FuDj+sKjxeeK1b7uce6TIXdP06nkqsiruG/sW6EN526QJ21ii2zNmudyukgE0TEPDnPjmowwR
DBI98fUrMQgFOXHysa0ZeNw/MIf7tUQOXJv7fMl1uxiT2jDBP/RgDVcENnQMMRS+MYMizCRLhizf
5Vyp0259zlJ1sfK/r932gsBgWvr0x7mq0UVmbrAZ4Dz7NYN0kmmoRAv0OA5m8+5NrM2pE6oLkCEX
mRsEF3J37ofG58EvsgKrD9PYb9pIwZmV2j8nf09rqto/gazwAT3kgxqw8q850AXLhWp+H97iRXHU
uJhuL0fnunmIYDUFsqXuNxF+ZP45yd4mKH+sqYDbvna6o5z8WIkPgG5rVLaTQZeQd14J8N5sCwmq
YJN63yqIwk8xdEtH1vFLkuZUv3eg4O/bWE7RYbMLtDGZxZEy/ISy4JvfBrETd9KS9hqPhAAOSQMX
yTxJYZUxqnS4HiJbKcxoZSXmqLDxiAxAw/tP9ETDm9xkHsmLIN3YcuNA7InUS8C36HLsNV7Lixxz
Ehnjr/m///g8V8Rny1zdF5ywiuyzYd5PqzOwyCBTMbc2AQVUsmdY+12m7k6hMTRSBdxZc2mrXd8z
38DONrhE4QhVKoUQ3DNQUmvEScBT9TuwnFNCc75nRG1clQ+9W4h6afrefcHQuU67zXodTdSowSts
vb3FdsnZ2MQ4HlXZn+2Innzabiidtzhlbk9oJ07CBgZ5yPPZyYBMsHFTFQXf/c9uKQtfYyT/6mgG
Kpk5U4wu4FGoX/h4wOBhwkoQ0Ap1DRPxkXj9hDnikuuH4GVbCFr/S52w4oc9IVSnDkMiUD2Gs00W
P+pNDDmkg5shmvo3F2thZliAvpNNbJ0TyIdV6sw5voT2PsA+KcfHoLD5rYRF0fnab3yN3CTThMkc
mPP9TyIrBoZN1I1IdYQpq3hUHi+lsIYQQxeCKbPN2r/8sQt/3hC73zffeHbz9naQVw9IYO4JRvvu
4Rqf4SfdIS+9N1TbCfbnlQb2MnqRX0Dq3JHCsO0TRUTCegBdwHnAnADO9TdaqODboK2ePbYvNV1A
SoK27v1zDJKUbVHjddRHRXF97xcXIkmb3QYW0N9KZ2qW9BNBr5bGEFvqWwp6dCENf6Xzlejs96Sh
+BXXp2ode4LzmayB9+vSItWv4o7uNut2ptuNW5bq4JRB+DeKArmKJF6Rar+AxL/XCv76iPs182+t
oXsU2ZLpYkN9hNJQ18TJWxmCA3079+eFf/9oWnZQB6Eu3ID5XmpWhJBPoKFyDx+qdAqgbKqiqiWS
21GMn6kb2RodiFKI7y1Maivc++LsE4oRkFdG3odsJQMbDAgatBgmbUs74UJS7q9NYzp2utBPFyuI
XZhscLC+1XLnxE6q7hBe7sEF81VL8sQJ8ATjtvpVfopnUqHHJhTXP1BvkoBLzCIq1a0IiQ1JGnH9
qLPS8Dr53r3w0e4YLYQ29T/5+5nbu9ybeIalt+XAH4lT3tgfA75rm5SMu0drVDX2fEeCBlLenxBs
JWP2fDvB8l+2T9TjA15qXydMllV6uHJBMoKFCsbWQURWt8em8Uyl9mIVj38zNBuGazsrfCvDaQx3
+68e2OsR5WfCRA6aSp9BbNiU+d0G7/YRI/+0EXenl4P3FRWubVZTjUmDsGstPXp7sLApOKJB8IZE
ZGQhBm6IXlzcYYelh11iDNasynvD2NoOSkbIjpFC/0N/baHwbIfNUWsEe1rDcvs2OCMthAK0DN9o
e7ic6yp5B/o0qy11G0lD5w4708HXaF4/lQhJ5C0+gisvZzrYhIDYIsu5j4Vb4VpwkvPheoqed2eu
3D4L3IE8bJK/NK5TDlrpwcwLo/DXVHTAdUjJIOtlaQrd8N3cKoJxqs4f6enb6MconUcQ+rWyu+Dc
6rdtu66ZSH9UCRlRijxsyuIJM8OBW2fijOngPOq9FBv7uHwGez20O4A8uO7XgLcVZ8j5OuTM1o6X
4TwFZ94Ls+aap4VQNsclc/fpn0RxGoGhAvc46NvA1Pjlw+SacJYKAt6ZPayZ+o3oQmRwt99XfscE
mAz47dUdk2B+dl/4b9/bikXy7Tq10ZyUdTqrOB4l9fmfHZaCeWqBZkWxR68JsuC3nMceeyAT06Bz
+r+87AJZ4S4VaSNQZ4w5SmjVrEYnynjXxprjnM7yAPZoLg7/3gq8oqGBPxCwRKAgbRK0kDjhxMe5
PYNE+vZrgtbuwoh1A7i063jn4U1JKBlSjNNSPgqLBtS81dlvM3gJACEaLp/eZqJoqYqoGa6CyCFU
A7xVVzEz6uvUwCPnbh9XvkJcvIn3BmoGMFCKrBfMNdHFogrCm5DLNddHKSst62nCVmggc8LN+fj2
P0QtVh3E63PMbFmCkixnT5Kl/4iLGeLBdFWPgypwfg2iE0cGohQwQHMskhNcCa3H3VAZwtbtB2+E
/S3RZ/0mg8xhJdYADPXw5RAtZri2wVU/biE2VnI+VXWuDymcptmsn8uWCOn80NArZ18It8+ZIXJz
4PrZcPyyfGO7C6d2KT4Gek6LfIaGk/1EV4bHY2WGWKIUlpIOMpahRMFseu8DSajiGa6PmEytDWsw
Zi5mMH+45/mgCHXdkeJIWrbNpYxAVzMIp7HfJjaOFRfDK+OUZliIc6zgJRpbGcXorgSEJpdt2+qo
pFvuyQkm+7a92pSHr49uFq7Ke5jlkZJJGzUIw/wAwrCa9rpJQ0ML1R9hd8VPwA87I4rnwX/InkiX
EDUsFhKGbJ2E0pN8JHo4Z1IstXoT4PMcOF21NfzfD7eK/rvJm2KbZv8tVirf3J0Us0VX2/i3HmEm
5LJFsYfEbpj9pOWAL6He6GeDwSZiLV3KxfvtB8+9z2++ezJnD0SR0tDuKOT9NNXhvS4nQ2BrACVJ
1HRhby1uvzIB/19JSCDs2KvlAIioo/MKp+ZHrZ4u1nNS+eBw7oWacKhfNcHvmoDgd93l6gtcngMR
TYZkQS7/CFNbTmO1kdjzc3Njd3NTbwlgyKldVXSkTqaPBs/QVKdrB5MDTByxG+/h1OzEppM6vb85
zkMXq8wLHvTowKoLayzew1SuK/vaZnaSAXfMMqU3zZjQ6p1uFTdvMvoLCAJx7xaLQGCHkYPk45oV
maUHMHbeZPCDw3/UBiC/QRPEXFb3LRDFM9OtZBVSsRgqitHIhqXusRCIuT9yclIvt3a7dzCoN5R8
+CL4x1auSVNMoTDFCMqrwQJRj2LA4w+6Pty5SG+6Cp5Olq3K45AJTfTz2ngJfryJpt5IYkoP46OY
3/8cFFzU5AjYdtyKhMBcDzkZpomVz11SjlLGiwAc4SRTJkEVyXmOhju65HZJuw7iH8k2yzEvdxKS
L0UYGF81E9D5bbd831CT+YWgPVHdUKEi4OAyq30qEzwEyHX34T9oBZMVOr9YjjdR/qsvb0cMGy3e
eyNAmnRuBwk68stBBr6/5NXauuX5VLgTtWzrVmQpNLDE3JoTX1pDCwS2Kyo0P4/eh5N7aaJyCFjw
jwFjsnEW0BjFM++xt4zM7C0IWisfkuhlQuN6g0aWYERDY7oT6ndLhsx6yHsNB8rPwgSXFqxdKJG8
hMgJDLuvtVbirVfd/6W+tgCz16qo//CffelAAwlZnq9xijpYxvuAQv/K9UGwV7XmOyHXZdjCXsXj
OP4+NjRFUdE6oZ2xanS0VgciQs4Wi/sKtQ79MgOvt9h5zVaDuUparNriZvOesD+0JDYhLXDFq8HX
PK/mxtx+SkfxMekVCLgfW+a31UGdP6LTVVGbhpnsV02mAGyJdb7/cWZgAveE3FJb64ISWCqWZtIv
FZJQwnkOwy/14UQ8KA3Ao3WbEDsexKQkGCerRQaVsUSicTz7adZgI3Q55gM/dkTe5DErr+L9H5eM
c3OZvYt2Fal/4NZn9bF4QYwCw0+LSPJricUfzImvIYh2WiggYClatzAPJoQGV074rvvzfWtmI5Xn
NRDIm7AuFxbYtTER22TqLQ917N2u2Oi19qroHUYJWu6BCNZNZ9pxyJ37Srsm9//wK6RrIw8RpNGy
HwQQhe19nnn8TAglrxQztC03lZompGltByY6acpxi4ygmmUjQj2+g+pYD7+pqcI8/8BbghwnbGt0
MpqFULii6z1iD/EwYL8KAwl250nEWjASplyRiz9trB5QeidtgdmOaOlRV4TBjogfHzjd0z9Wd5L6
iAvowtwlrqmhTLSdKt8JXxRY4bPOgTmESkBJT0zfHqTyQm1mYYuA9ucbbBV7+vwEwSXYHgVFZtUc
m3X2gNl8bmDrGRkbsD3x1IHQdveZmMJqZ/p3bfIzV9uZkru8hanvfvAYfEogV4+W46HtIv6EZjRV
YGJJI4SkLwEO8uvujHUW4lizS5Gcys0Rp7CgH/9woIvvamfJcs/cI3DCkPiBvSWV4kGb4IwJjwbk
Rzd5WjR4NspZjQITetaqEqvJy99KZUX6i9nPlKgdUu5uApx6c4dAfUyRFoSlDqlfv2Yyp/VbB9kx
KmFretTWjcPNQoVfapqrALkEZifkQGc5FQpT7l5eMfXW1YetT5j1glgbK2Sh/4mOx9gGaofAbqOB
ncGr3YS/TL9ysJnda7Aqr9vWQqmwgpPNZjWzaA2yycaCzzrZm57MWG8k19Z1uE3OcH6RGjDXB3BS
ZfeWUdF3K+TiTs/WIwtcBMYfiysNQLL4cUPfXhN/0tFFN8FUnVriytbuEBOl/gtTltVI/dOrDim6
qbtN6nNp6OLiwQC4Za8i+wi2Izs3WBs5IyWGX9cqeshFIoFOq7goDZPHBNuHKFhrJ4Wpr00j7N5E
jZamY2F3QgrpkCH57z+m9QlvMn1kBkqoTkb3XkIBHcc6SKJtu07OC+p1QST67sa+/2BiJIoA5VcV
vI/AidQLDgy9UcwVRbczRO2qsWfU9VjMCyGEbg7hMOWMai1IjAfhUeMJ8DQ9yU4wHwmIO1sFgMu+
YCS3nV88y9HrkJLUCnsevTqSv7aVUXa6Seq4HHr9f1zCuoo3ud/l7S+wlcm4zp0YrhoOpgL7+Os5
pYn0hLSRq+OwVEpa+HpmqqFIPVjR8ZeJGVw0ap68mN4tBMzSaOD+CqEIIl6TvB8xFLPFmzGC5xn0
86GsoNMnAYvqzZ9+375zBDwpfph6AoAooJ+X11QySNfvU+2zEQP1M4uQKo73crhi3HPB7noPrtIG
7q+AkygG3KsHaP0W+O3+QAe1707Jp5wO1JrKiGcsGhbjoCK6lAtyhEWLNXkNFitjYKiHFy1d5COA
PuNOfB0lFIj+M37jAvOCF+83ioMhgNIwPbgXb8ndkTmFb1AE8ifmSi4+zKiyOsXck+hbWvp9jaXH
9JLHLkW614+2rQ4kq5Ekb5/yt0A9XKpYEwjDrfjSqMkgaRBFJEBwmWOtpat65aS8ooxMWUJGFZWS
nSywuvvcfzJvRMbvLupZXDs37y25TUgoxrSMa4IcAVe9OO1B8souNiqCDTlRxZXBAQ/CrznrZcil
hQqW+nDN4GAfdWBZnHa7oF12wQhV3Po14CpsjOLC8Qb3++nqs4Q50mfWpP1P7+Kju7OW9EYHSBhV
cbdAHJTV3aI04WYE92usLW3NlbjHf91rqdqF1l4dwSisKlkWBQHR7hBXb3RPmtprC7d4uH0R3Lc9
R8OhhSss2tiMm8Eu1JGzuvOxNFy2pAZNGUz7dKHyGnYMYYXqRr5qOBM9TK6XnCpjtY0zoAWrj9ze
/ONYfWPnx82Y5eH+4X17pKmD4r33DzqTA4AXyHhxc1aMKXVPqrNhKZ72b0l8rB/QM+TVA5txr8mP
N1PWbdvqBJamUCQCAlwlFgu49PS7YLMKy0qsF8cg6iiOOH+1LL1RwQ1L+RFFUC380L96OvCY8nXv
swbYxnU1yzfuwPCN8n0aMRiJOXiV35ehB5Jj3GKw74acvCc2PHisrt7PyKKJuowuEvDwaAL1F1JE
3wukr0RXRG+y2J8eVzVxe7MJB1ZqveY0r8QnSiPVngxbF9zFOoBIsTZz2mvpKWuylXnNz+srqRrm
QgIEoi05w9ht+fLsVl0afwcyb98ZxlUKdEvxI3AGtS0Qk7lZ2AUhksdi52AJyKiKLcXIiSpEweSU
CeMTy8oXFYVK5fSC4shiaxiLzj852uo9kInqjGG2V6tV/0LT6JnapdqfzSlzWeQX6hSVe3rllFU9
o8C/eU98VYCtVuRCLKd0cSp0WTDRUzdjLnzhObkUGblTw3llGynlS4pkuXiaBef2sTVABbb2iWQJ
g7lNuopqA9TAbp924aPrVkOgf4dHldZy2XMr5RHHjI1Sm++sshCDDxSGKllbYq3APi7OBjyp3JyZ
sH3LqSIxHX6pv1aEO1nY2xz2ZuvHm+JagfjYwJznk6zbZyEeLS9cpDf1kfjFDStkDDsgBXz3+4Dk
FNIZVIwbtHJD5i8ZDMMvfJ39ubWTEe9gYAHzvSDc6Gh1LTLy1DMZq9Iltqvrhqct5qtowQxoA6CA
CLwoHaKc8+BsXH6UlK8nCoNq+jGtK6xA5SiM2C9beyi5DxTPI6g1xtLaCNrqnJZihZ2ms0QVPRZy
rzxlRGFqC8hlzUw3F9Lkz2H4q0kQ8RiHapzgkZKwr69yW1IrR3mCe5Vriqx3Drn2EjkxiCau0M0B
gIs3trFIeQYimP0U3FhhIHU2L1Qe9EoTWLK5BWujIH+BEl0O0Cr5SHvGj2/gRhcQFPR1G7EDsc8E
/5tlijqHYDcj4TmN83JkShXHqD/JU0wQm20f8Iqx68/RpjKLkNFhtgG0nTx8Hl35fG4y79KR4LdP
Sm5vZvYSDdl4S50YgkVI59YgqcmRNcd4JfiIBSbqI0FUok7ZxqYpKgTQTQjXBEI7zCyslz2FDn9U
kNJQJJ5AAvna3Gv5ury9Hpz0j/aYN4vr48alX1DC/2FXDQElKtbelqumRUPWA0Qo1jwyqKdMefUs
UU4phxDzjaiKGdnw2Gtz0lptFJYwL6QCj0z+jAHDZYUpI/+3YrECOCFWU3+X/EDsI+JUkfPtpYW+
Otr9yRvcaYRH7ex+CGiHvglp+mUGRYlgZfmnOJvnUi2YthsaOgJFUvZbf7asyimEYAFXW89PTnOW
FN0GhePVqDWrAYuuIUsdEDxi6qg/s931CaAiudgu0T/oAK2j5dx29YNYduu8k/1FHIGwZb4qYxkC
BJFEQvK6D9B7L7AZJeKnqpgP87NuLjQOJjFeatFJJl+H3khswfbAzAuIP2PEaoEdkJbsq9KOOvDQ
N49M9RuWu9ozXqFt3ZC0YTlSMqz+Z/zG2vs7KMVCxIeHlqVyv1aQgNJK8GKzxJUz+Isk0YANuXFe
ikWZ6z2oxgyh+VXEeAT2GPlXPW5kROSZFqQn06xCnu06YRRbrSh9PC3RaYmYHl9rg7SWBcnwC1pR
VrARPHvPxscXJBPOS7EsuWLpJI/l7tJVSOEGVXhPzUw5Mmj01dYaWWYuFhafLWddCqxgYHDiRe1b
DcXy7FgTZhg7n3VeUvmHRCaMqkjXZsD3u9CKpRPl+SzDnWSlBUWLx1DFl8Xsv660hjYfUU67JU8/
j8wKhwSByeKUzMNRBGOz6DL3A2LwyRaR4SBLU69xJA65IBR83xRHTiapMoTomPPtOHLpSOZ+PL/+
3bYB3TAClhDRuTpOCPfQ4q5CZ5lkeRodoGNK0V1m7XEodEqhTqdOiTKb0NFDzjAxxrFXHHXvJBrm
hDA8MD8/wK5vV9gL2riOQ+wBsO4SB6Luzt43/nKHRs1l1pOWVHWPX7ZqyiJRkj2gORl48N7eWwi4
0kWK+9tKK7HevWYp0szCPba9+d/CV/YE54er16ERMp64FRYNLdJSxXJs0VIP4RrxTEMjzQ4XZWba
HZh4vR2/jINymtgqVqrozgiuzy8QiR66EGZElAwBr9+hYGmgHzn0RM2iynHcQvvP5r0lJ8G7YhqZ
MRGpTdtKFV9WIB8qUs2QuyXx/J1tCIOZ4mphefIjG6lqYLQMA/mvo/dnxgPPU2Id1Gd7ipZGzwIe
FmxBWryqKZqU3uT3+sHo61mOFuy8MPO8R9K2wcu3+lou2CxUefdatLF6sDxViJBcMq4mi+JCp+r3
K6U6OhkDSIYvOiNNMB474CoGBuuJwI+f1Zvrp3P7Onl27RbqPlm4pDf9l5jE/G0hrP3BWJcLpkaT
wagCHy+tV698Q+L6lNWbTjaCtpV/XxGaQfuhYYPcsPf/cQHKq+dPYZbe3p9e9wM8fW57LWuFadP9
WWxaPh7gnRcu/GHT4GEarBjxtc2O1SXoWqCUtrhsx5IHalCUQrtKfTvSkI7iMujSlczCoV8dF5ar
C+ErAyotFclc6AUcDGhagpS+IZ5BrI+ChJu2dTL+dmiMzRAEBy9+IH3b1OVPfRh4nrQpKftPdWDE
PVp6QGwL8m+LmkqJ4kGR7g6J3S1+SZCcx9+GKAnkoogeN9Q3R4YKKF5wQfjAxXl7dtq0VUCD185W
sqriBSTfTObnZvPMlRRx8jgLlh/8spw7HrFzdHX/h7lrZvzhG7O8HTVCbHSK7DhoyFBcXDrjek79
8HHVVORGl4xKnN+qnOrNN6PtopfWjEOojgNUUWLJN1Jmg/o3R41HGX35GXXSJmzcKSGpHe9El45z
RRQU6oorkZcBO37WftR9gMpuANmLecD92NnQV5z5+W7wUjpvYG6D3cpVbH/oPeg1/swFjtbdNmK2
Srt48OU89IDwZnPtx7Rwwl9w6MVWkd1CNq3ER8N2Cqj0Oe9XH7pmYlZsaXevBUwU9a/mPF2RB7d8
kVfqJsOHhG9crCl8QluagI7/elTKMsm51xTAuGFNrD5vxZIjIPzOvaxZuQT4kby6umiHkPtjoIww
pdVHN8KtC3mADpND5tr1cFeLgSmcm/m4YJf14eJ8+b3P/bNJixMwe9S+0aHqm3djhXGFGX+nBE4d
IH6ETQgo7xmeL9ulZjzNk8cx/h1V0ELTVhjg5Jo51aDFrUh1EiXzDzVV31U8BtS+UN0qO18N0Y23
F7F1AhplUw/YuhS21yrpiD5COKE5zIeJKfcNmKQxp+YL4PBPzZpdBDB6V7zMF/NDu9qTAW6G8dgj
uycLyEYxtWUtENFtqi+HhTENffa+Gmug7WBmV8H0D3DZ4i+VhN2YGHrrL0Sf4BfWvw1cuIUt4F58
uPXnIzSMEDden3ZQOH5jXLDh80+iBlNf/6VEfdtqdh0h5PHSnGja9jpeDm1cl8KiwQM5+/wbWNE0
8f0HrjTEdt+/y/NLo/Yyc8qbB0QACtpVh7e9qOZht5nS3ikjpiFD7rMImjSuAYoAR9gz1kHMHPfd
XuzNACHZYkMZZ+k5FILXN2HYmKpcODzM5BP72ChZmAHoYoItRdY9u5NK6GJQyJyHp5EvosZiTHIq
mM6iJmF4yZTItJCayY+f/uKzewEkwUSXY2No5MrQUfSmxE6FuZVG/mNLaBko80Xv2Ab3g9AKvBeN
FcdUoCTgMblCuVjB42or/Biaqw9PsGjlAbr8sZ5kxDzxQnda0QsaCBoanJNhUCU4G2sJ9gzKPmYZ
jjdacX2LFRrqO9UbT5JZwWq0AuVwpP05UpPeuSu5nH22LqlGKOsppKUE85jdrqqryiReOFBKmFvB
1OfSMSY4/YSa9iQBqf19ZJrKOoWXhfCCUOA6xSfkSWKY4P5/yK/vtRbPbp5j56aH3uCi4hc74G3g
+HB7Mj08fCOs7d0Ebl5+jb1SF0wf9LLG9nQ7V6pLeTIQ5kQOBaq2oG8OaEa1aKknTjvd3ZZQh0mm
hS3Trxz3nLynEXSKjq7Ny82Mq1jsbEQbjeTQlECVhd40v978a8/gQpQT6pJQez8PhzQ2Gsf28/Dr
H46QkJgpYAxgt21iFVKPwqyafw1K+pAOWcvuft6EtrIb5tJjykNQhxMBMBbiY8q/07vxkJ9h+tCs
Q+o2sE06HdEpc3psuf3TjbWvWLeM+uK8bQYSMvch8/Zlr+Bua/OPNxT4nSTa+CIJNTtD7gix9Mng
2GH4l8MLXQqzS51prL0fCRuPhzKNS9s/lBQcP+wqDHVS6FfSH0aVfwMfNzGN7HEeOTPAfjoWEXfB
UbsH/1XRThH5aCulsxQrWOkyySMZulf6wG0M7bkx2IYpiJYpe35YK2ea3FfrIngJqPjWmafgaXDb
cMV82ASycyYvbzUgGIypMsAmNFJ9NK3hHMGJveI6yowRiSPS/6FTKSqiOpIqU0Oj9p07KVcpCw8i
6FCmSQbCQshmwJ/xA4U8uq5S9JUSvHSAJSS7WaGEscaISri483x9mbzF3QqBu1+Y21xIqEJyXHGT
iQDZEJdviUY2GNwvxLUXiPIbEFeLPSj6XxvD695kaZvAZcF1jqZuRomCpjkhORr7/8ODgyDFJiCZ
kQy9ivK8omXb7rCvkJLUGX9/SLn959hYccCUlzdnC92sYgWMO58nLvJY+9zsY+K9GpeBqw0X53NO
/rcbt/dFqzTQ1G9Me9G0tZ+RtiROYAmDmxv/6ru4djgrZrHRv9nJhV3VvSf7WvM8y2M0bFF9Ysio
Hycii/ixxZHcyYMF/bESOtA3UJyxvk4U/kOlbfZTFpZ48y64QOOijdMWxDmLkQBeGTLVw7mrdNXu
bkIoYRB4azCyoSUr+qPcLWMe+giGkfLnLIDh+HTW7HEUTl46HPrK4zU8mS034Ul7GBhmjUZ8aTQ0
UQZi6eJ+hQHZZNmzSYQ3dWF1BjRaElSJ/dZ1bN04gGaB9ZJkdOpTbl1oQNL/jOFA32Rt++wp3mGX
FV+XGugCPuTVkENSIV6rFy5ivosgN70F92XanqS6WYswW9yyaR0BmxjC1sjlbrD6+nb+bfqs/va8
ROCZBKZYu5PdiL3XqPUETNwZV3+3dTmIT8lBFRwJhDtCyKG9O1SVBxeM/WZ9eQ+XOUsMxFK5w/HA
FxyOXqcDU9PUCemV9SxiYvuKwTg6QKLL5py5uTEkTa+PWFEA5Qn8McTq//7MJkWJdTO0JGTBFuMH
KwIkj6lrj81GGBN2x0vBKdwjl9iKof290NNtpQpLWcescCwuFP5gwlmI88hQ+nZ3NfJ9gXL4jdNB
Qi6ttqIhaj+jp+mNubZeDIalAL+fbSwm+lJA3ymDTfl8cTsf2jqquK8serXLsj5aX2XKPj6GcKDe
+MUnk7OF2Y0AjPkqpJhJ+7XXOPMRzTJiEybidxr+U3fhraGnQF9O8l2Cw3nVK1X8RKab02Ed4Cy8
9zWxhu+nskrytdvaGYSuM1lBs+OTwqGQy/UoNjNe0JIgfWpm0EgaY5ltX8hLj9kA3lumk5Wmb2ft
GljmKKdjU+8E0XKX1lnf+KRoFYoUTMNw6nBpbb14qt1U+POjA8B7pvAUFV4FQgC99UL8bWWqPEhw
9kum8GON4dqXfWDuN+TOSxvA4DLrUl+p8vkZVXiLoYpkU1nM+VQ9TIn6x1OSM0ZkYYOo1XyBz6E8
gnYtqtJdOC9JjXKcVLd9yqiaGRGg7OC6WO2tqEfgb7Pd5qp9bomQ5SavUEVLJ7TweUFWRbUnozse
slK6CwZZVfRtsGud1h+B7en530071UEL9JmjzS0312L+yQFsWEbTA9F9Zx6MwYnm2GcFmBYNazKr
KvTCf4NRLjEpEU4Ro+m+F6gyHY+2Lc2Qda8s+EMvhzyaJjc+M75S+ugT8bPXL8IsxbYBBw==

`protect end_protected

