------------------------------------------------------------------------
----
---- This file has been generated the 2020/07/30 - 18:15:51.
---- This file can be used with xilinx tools.
---- This file is intended to target xilinx FPGAs.
---- DRM HDK VERSION 4.2.1.0.
---- DRM VERSION 4.2.1.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinx_2016_05", key_method="rsa"
`protect key_block
WMOpg4SrMMlHqGXN8IHlKTDWrq7RoKeOP4HRFubh8x+LzOqJL1UTvmU5NhZnJcAF2az45D8roVvN
uuRBPVB3/eG1kLJ0Yqw1oiPsd/QIgQ84W6NO/Cd3/PJKQ5/KSZ7uKJTS5u/EpjRjS8al2CCA5s24
aXWz94RTqzGYXmXvTmXggN63K5DiYeWXqOfZE+a8kZB+EWxt0im3Qb4YQIDu6kojz3KrxnibwGgb
I7eTaToqGb9V+DWDBBuUYLbvArPOAJ4+ezYtdblyU0VreEw9TMMxn3dTXElrPq6O5LCHolTUD4B0
/nFh6pWpBKI4a6jFmi5mBhr6bq4kS1lrh9kHEg==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
Ts8P3uIXAZCOBJ7oWxAxaTxXmWb2AOTxQDjPOMl/huR597SGiOi3HpVUTCSbChwydezPSN148Z/t
D3DemuyoM5SYU7jQWvE2GzDWa96/pUxC86/6y0NIIh940/uMs9aQeTs7HZ0Rfu8te8Jp6qs1sIUT
+b1OCyWIb3wDibKM/mntM6mqTEnDktvwAGUH37DaD0t6Tkv4AE2h29mbUiSMELvNcQGcVEtt2/IK
rHy0x55y9cOqcPO+R3dC0zUVaP1rVqrEPhuPO2HpQMOlZQv7xHLZwzHCi9xbGudC0F44MeXtU3rl
w6OW2vznq+5YhXj/DODC7y5J0IUd7zbd8Evo0Q==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2019_02", key_method="rsa"
`protect key_block
UKGjLME8onWmp/H6BPIGq2Wh3CN9PL2FsJtkOT4MVEywgKykJWrd529BpgNWW9dt6/WqXmrN0Q6P
o579KxG/yFRZd2KnerJOkpZa6nY7i+yDt5RvyAU/z0a/LYJsVWOG7CMgUPz30kXWEZ8L1JtvJWVK
QnMk70gWnUge2WZKMpNTP15oUK/yp0ZJirpQi0FJ4ylfJ6+RUo4L7vty2V0tIIdLmcco82HZTWMY
r4hYmS6FBf2D68HXY+s3QC1Qrh2uVikdRNZu7X1Fx29v6H34sLkpclNU2hhPAEIJMY0gC2CRj8DD
5iB7Qa8ob41BjGFV14JOY7vkE1ywLMmI0MQ06g==

`protect encoding=(enctype="base64", line_length=76, bytes=851872)
`protect data_method="aes128-cbc"
`protect data_block
BjbhbinR6Iqx7guPrU2pg0vq/GBXRe8BxFb3mO0Vdwb0K6DiW1ftIYwn2C9dX/HFD4kroPGb6d1w
367qPcMjB9ZmxMeHoNJFOaQr8G5w4jifganm7Km7jD3cFdvSRtAp/IyHnGusUbPVnCL02WjyEFol
PfPfuZVENyDDXBgAasekwsnEbHThbALnpr0PggCg7V6spKXDqEkLmUA925RO37diVUgAK1HrEjUd
RnwkgWT5+O50vk/8mAdIYdJj6dWZi7++iKk1w1gvMRibb6Eg5LJ9+hU2//yaX4V+qdtJG2bzk4z7
GoofXyAlADvedclcxSNZNdqVHiNMr2sToZ/fiYa6dSXhfZ/Dj8ApsWSN/xAzCs14tIz7LvEMnCEU
rn9ROJUDUf1A2Ae/worTrNGu+sHit+5+m6EjPlMjf3ZjTjI0/4ThGZsCOQg2qcDA1Ewad80ZuUVd
ACiY71DN9JQiP9BPDq2ibfXePvxDtWS5VpzT7S/avGYRtudxtCZgaBH/k7H7058o3Tlj/UyyzLDv
tdIf0hVvCpFtzqFwoM9ReKlsJOLYzX8eL43BP/CLTXoo8rmBOD3WdXLeE3V8VNF90aAeu+4jnhey
SZpsQV6CfPHxIpLKQEK8WO5rI1xKbJ6rGE9XJXCnxcuy2gxwm+AJj1bx0XgcqLJ3FjxjkmAGT9Af
BSofYZvqaktKqLByr7MKFOzD8oMkyvIwTIkg4xMTpwi8xJnXvkNLySDs1WKKRvfs0Cgpt5UYTqu/
SuI6za3WD9l81DyqcbSbny/obNM5orm09aI7PN433tMaAZBmrxDifMnCmrViIGbr7xFTiXX0nJ1q
3EC5BnvhRmSz5l88YPJgSTlDvDxHeM7vHmURrMp5OXKMW8yjdPixPn2ldd/juCU6ODGgy1iQLUBt
ri5uArPKbSxxynRqfQ2ziVd/MkoXlVe63RdCm6LjbWHJENCB/g0z3X5Xpc6VFAwb9dDchlA77011
Bs8MlqVda1Kw62qdtSVyClRAEF9ghi2kKVDV+0BpKWzPrxpwz4ZxLWrhy4F8omN99m3TjG87uCqI
xZskY4OZy5zhZRgLB2L0BKg+q/a9KP2HQd+SFCyStbWxZAdFxB7ttN0gSuFV/esOB/k70AcR+cE9
zCZfv2mI8++vPfSkuTXlAyaYXvPIWsuW8OSKA4fVwG96O1fapUkICyVe/PUN86Sy3+uUyvdjvadh
OPuqncvSNBZspCOX4z5ig7OsD+MP20ZBX/z89Anr+Ne5c6a77h+fFym+nRcJXyWlRGX0o6/bfUau
u99E2J2osvOMIeYKc7J7Ci2QrTOVtXU3lzGibXV8DE+gHkx8QoV4kFzDbbj3LzlQfz8sMNjb/C5x
oIPBWb9ug0X5ZWF+1hEnZk8SOLh8h9/uQgdI9rXOwx8bIU60QuvrhliSLaQwAyYtMXpFh5jjN7/2
PnwQESN/tFBHJNTd1WWWX6If695ucUxrb6cpF3LG/EigTIePFHKGp54tuzD49vMW2KKAtRQyTQ1S
PYsQWamEhGI4xPcbIKe/CElBfe74lJFo1zHleihV7DsmVbQiu3JkUCsEnN53pGnPWVVQc8YMwfZC
99xHg2SDzqfMFXTyj1x8x12mk8+07g/HUV1CxMeh++0tHOHfPVnSPH7aHqva0s4E1FpRR6yyUkXo
5bwDIVPEIkJp67+QLy7IsjF9yQGUDyrBa+jWb6ilG7fFFxspOxbh85oqHpeIKovIzjPWPKjlYY+6
Iacun0Jg6efCj+MY6EK1UXumiNHzMtkDWSIvPlyz0pifwyOJ70O35W6bQCCEE3oL5R1y4aV1gGtZ
q2PBILkjSpU8+ILIHtl79yb2uD3D+N0932zPA7ntZPD/QZEHg0VeedUvw1BqD7VfL0uXdAaxk6Dz
FdKNsF5AoR/mccMRGjDvmdFnyDGxZsl55Vjl9COiQtu6gMb7BkybZSwy5cvqVLJUHDODPPSBDMPR
/oWyrdNSIX//R+JPSvAez2lf9rLStOHENXmen3dh0tETUA2rs92MrX0Nomi5dY2ds1e4scsbmmxy
MZ3Zdr8RsSj6Sjv0nMOxVcUzDPGRBfgRmiEFaNQEJO8Ljso8Kbq5QwAAQs0gt2NDbCFTUcXIcvYa
Sa2vinW8+BCaKhBc//PzWLnnBdGXY7rhSqVau3T3LazDeg+7Jkn4Kh5DpCfz8MSyW06huOffcBnU
BKaqGwXMq39kFiwHvoKiH9Hackx9Mj8aUks/Lf5b6QvYWEJBqVc9mJ21X2OVnZP27D4PmU9orYzs
XzI76Ij7R1OHpHpv+gOEY8nhejgi0V5MYk3Q4/rRLIWc9Hjo/+Mxqu4Ws0127TltlWSRW8oMtEFw
2kbEGHxHZJgoqJlYGf2kPaSgEJUp75sl8TeO4TrBzZ3+FctSGG4pqOxUYi9P/nN/DNZVBC7LenkR
xLB0fF7bPpk1XFoHMl66eU5OEp2VEkj7BA+fOEd9oXqD2rCNFESLEx+xnv+MXt4J2t08LIKwMN96
IEseQbPZKsQNuls6Z4tBny8qeIpphWazkOd2nbvvntyerzihgmWupp3i3IDhKjkP2ERd2VW69D9b
QjnPnMSD9HZC4NBvik8x5bPu0xM+IlOokwsRk7umS4sp6DY+iIx/xRO9CnuhFXRdMqkuKm/RClWX
X5zXKMt3mABM4GyYuzA/oesEUkV6IyYCpRWn39vt/XSoqaP4L0pgg0rp0vbWTwbdid3Pc8YseGWx
uKPVAyGTi+vYOpRh48cJokijbBtiRxHdulYwUsLEMJUNbWofAuxbj6M1Jz7vZ/iS+sUX2rexnGPK
7PbZuCq2GT9EgrHaicjMXIFWMj6Sjb2mQuvs3m0LBS7LkrxxTcELIjkhyNcX/U5xwEYQdZNwQnZa
67ySVLMGUCm840S2EJIwxRxuaKOFHjdHREPSy31+wQ6uxKHmfAZp7lWbfP4V9KQCgAreeRhvdvq0
cVZa066iSQzjNlW5UT8rJKpZXuXcWqxmMfG0hmZD7FnT/XAAC7KUd1GerzGyftSvr/GxorbFksHw
xQ6xVdxqFmu7uh3ZPl0bTSpMAKhTtLhfMu3SXLY+kT46mPThpE+iBheyrQK3TgJsMtrNUKkhk7gT
hYAWdf3g6Vr5KWLP9tDMINpRPA7aC/qLGOHG6g+658hHM/BbYFVDP28wJPmoGdiHLjDCfM+9hKuy
rWg1YheAy/uM9l3sYxNuhDJIFCKgmSc5z9plbENqHP3qxXRU5i/n4rigQam5soX7RWByMkAQxWBG
A1FQ71larLYgR07hOdh22EeceV+28RCBA06BZCPGrRF/jRH7wKtEHLnppsuMvAa305Bgqhm0SFVP
nEwJGbkYwwN1NgLCB3tT94nkmuCmfpccPzCHSbpAKDUcDNBm0VjOay/mnk0WqXTZYRNtjqu5Me8o
L33aElQ84O8CgMZ+p6T6T/Ovt+u+eFWUmQehGlEWtlbfV/1pcZG+GXkAISYecjxetCNem/stqQn3
EwhP4MXH99SDcwbkbjV63d2OR0TcxqcVeftLptZ4hJRsvIMv8S6t1aIUyoE9OOTTiuE4xQUpK6Y+
wYuQ0iJGflFsTIdrbYl5jzq6VdOxE2Dx56fWgz+cLxhqNmWYDkwNZQx5g+RgRIvU7AkVprDAcKLf
E41v9Fq3UJXzrmYLebp6GKnPhFWKShFLJ12M/uUuJApi0bcnEBveVZdN8rv113GNibKHtzOAjCUR
6SFnideR4xIe8APiFCXw07ciy1MKPMqPaHWDavYk3h1P0xtzkMBWvWcTvKP4XAY9rXUlSZ9u843U
MnbSBprYN+1Aq3uwwfFTiJVAlkExH8KS3NEMlsWcknm2/csklPsYZAuQixTuhvYKRIoP35wYidkA
L0f+t11HAT0v+wL/L9lz/n7SRKoDfDmtTVmunoKVdPrcOnvJNSqdnobsXh31k3HDO29wmliQ9xDW
eeGwaM0fdg0jGnB8fs5lJHyS5/wNpDUMPH5q7YyIuERDrmJWN6lzvMSkgVvR1LUQ4w+16P0BXWUF
LIIEXNcb1bIWfFYB6s/IwRlvx86C3HJ+fOdnp6qsqe1dmqJikCjYzKiYMAfwnNiuMAN/LlLIfHDI
Nee7bY+jgkJmxWV5LxNWpYNuzR38nIpj/10+2uRCQMdBB+71JJ/zVIVm2HZJDC2HJNBilA+/Tq8L
puDo78/FR1cDpDJWChsEdHXInp2gJNHTV2EMFAOJvMwsbjg+LGrq0wylwEitZ3jhYf3ZJvlk2p2w
10TaPNuYK/Qq3fhb4GXhXy0s+pz+zhwes7ihGkVWesZW90wrq6AsXEK9fmtXyml9hctnGkTOp144
D+o2qDDTC/KVHbFyt7er4GhBgOW3IQP89D92J3GeZkR1okTjBHGnnLHREvjrRjK6Pj7XPltUnwdt
3bRnhntxfbCRIjTw8ChqHHDN1Y03riokWtuO89XYQQoIhM92GWxPCuwwloEzYPqiS8rmNkFbCWCs
fN+j6CV+8wzBAMoWdEUTmOuwAOoBzkVsTn0QmidK/7rCCv//O4L913Bs+6K6pR4s3u5SdoTYRqT0
r+M7jtVsdQN9uLQ9Dt9KoukLMWo1+DPFuX/0qnQHXAsSPReAkXgnFU0X3esEzE4EFFbUyM+2yCRO
bvoKVqXftyoZPrtk3ccRZagi8yy7mglRvWDrgdioQFgp4E5094sZ0OwunBrsjESp/dqoiyCJ2Scb
E8af5QqaqNYMghbKZ7l+F+8s1g01PKPL2ILBAFU7oDcI1nlKvACa9rZ5m9FtDzJqzgISdf6TXr5A
sc9XZi2aEfOvb1kRxVd2DO1tZAf699k16VL0YHHskv3h1cPhfX6TV7v2xfgZYAPZKxS33ZMoUsJX
6A8M8/LUTJpfnQsjwV8hChWr61ZuHqLLBvaPv8LxfUp3A4DhiqEoZgL0mUm2f1FeiLOLQ7f3oaqn
BgN46rbk0WC6j/IW3jV4vbjpnJraJp6G3/1UOw2iqqCogz3RB3q2RSEv+qpbhbBNao+UII/bNrXR
w5TVd4g5ql5KR+hfpcqBl/m9lhfM4JShUah8dhnKp5IhYtYhGGKM6LHYtBddjQRlnDAHDkxc0ZKF
gKylYKrJVGlMGsXMLSVpei5o5RtVzYpXFsjZH87K+Fv5kzTm/j6vMmKmz2NiSgqIrdDv1OCY/Dje
YmF+J4yRhy4ROEdNu9+9EUNda+TMUIcQU1Ct3kbEpCfhSOuC+KfaAo9CJmJMnzH6xTUg071gthgW
Ei5rP+hNE76IG1O3k0bayM/BGsZH9E7cZOvLcwa7oyCU0T73BUVMIfoTTmO8b3Ta+7Y3ghFH29hO
N+8SPLH9DLrvHgz7ewiwWAoP7W7o0S2nE5vVpqKsA1M3ioC8BUnNOPxdZOn3/VJ6g67c/H7Uw9pU
6OJgP4He90NBC46+xpKs5FwpiebimJHWBs7PqhMOwGyqcoC2GRFnREO+L+BkUvyZ2ZGK1E7Z7tjm
eYdUP5a2lf15eJ5zxSTa4yrR5PU+RMk5L4khxCS+ZgRZ4BBnU0UdRQBch2XSta2YAOQbxDFhN4HC
qaB2ZyGnZPh23HWcn3X7D3Pxvhb90I/2f2qjXfQqMO1ud/4Vls1SNPwuLhMh6FtYGRDiWSK2IfcP
pE3p9935W3Xo3mIuIq2Pv/F9nqR0/pYOwfQvgTUIfOL5bmzimmGpQo5Nei0WlhEzTd02Jm6Sa2yX
klFpQ+HgDffS+mzkOA81UzpIEVyAhNlvYGfEy/DpIKOdyzCMDFgbZdCk9wDQsOy6SwCbrjHEjWkw
abN7S5lVDhCXad5tNkWrVn3Vl6bIVvcxzQcZL8FflwXBIgutyg60NoSNjx6qJsRP0JQdGduw+Np/
5XDwT0xGMksFI10sMPiDXOKSyGC/AFsklQqBOiDWsZl83aLO/LV+LqyBEvg7F2aqu+xKN7d1KFel
7rHov7Q+hB8WbNDKvgoz4vQ3ePVxejcSdgigzWSv/FVsKCCtvJgFftIzjMkcJCWM96ol6orF9+o1
e/YOfPvlUIV9RvBynld/uGeHpPCX/VKJoVbg8q5Ve6WjrMZvmnZ1ZgJayDFLZZRs13/YkfTbxrRa
176oa8tm0BtMv29JeugeqAkSIrttV3E7N3L4L++7vfFRwbzOTQz6XHG5iRWxrIII5uHKeD/F8WW8
Aw9iLgo1CTDw5GVXdevDPlBeCmEW1BnA/m5b/eSsHrH6bYZkgX5PVo2hLFbVDDAUEgYZsT6LGSOl
9sf1xWshhKm9aqrLK482zG5KKuB3On6R+E9Bpo1MymaAQxtKmHBvkAhhGOzn8yIzQPtpZcMSe4h+
kmbF7xiukisAjYjHdDSZ10pDtszh6IRmyzkaDsMASEfApJJFpefbk9dZtIBlWwpsUr3JB/VhDlea
pBN5o2mnNlJMCZ5jlCmAYcObDSw8BJ+Ky+9FZYeXYpk0DA0n+oeKDZSrqFCHVdh4ex1RPh+kTyCf
8izVBIbmV+157edhNKp+0RQCNTzEHyEmv6xX+Fv6rpvYsrFfphL8M1P6tesUUOYyweYkadyJ3vhm
M2FXOlRenroi1up6LHj2x/XAW++yxi8vpwunWjpRSau4xQ/Nd0lJJ0MyVGX9UTgSjyKObKkfDXiU
1DbGqGq0T6+DYcBI5prdD1uQd3vM/jHDIPrQ8N56ke2HLvSRCX2IIlv8+4qqYPs5qSpB8aDyskxi
2xjjMGFMsMecovJXB5c++p9Ay+JhgCFK2/k30Xri7epPf22iO/FX9WtEXMJ/XPpyMd20ncw3Qd4u
RHTwAmmYl53ORO+9Q1PViKiMl5r49EpoE7DJytIp+3C5n10kj0Sf3Ensc0wSjNcEnZo/Lf83DYQc
FSRJ1PoN86aywAmaIk32X8Le4Rs4cjRknzGyOG67V74nM8H2xgdNzZmBxQUhwBEXlPrm8rtT/K3d
yhrtuoCygesWRsXe5aqo2Xcjbm1CVKEHfoimpavudeZdIimcWAJzto54nECATOLDuCIfOw/hiwUT
YaGA1xRTwKHmMuG9NOXXrwig7XWhGn5cVv/boIW/AxfXtoO9S5aH0+CDqlz2P1ogzgl9NK44wmTX
Dx4Mnpl5YTQxbSm738sBsG/87aQn06TnmdYwYKn4d+nDSWjLwN8Gpg/7T5LL6ivluwZavHRWmd3d
ld9c1liG6ZpDKr3oqLqu8fLcMCzoameLAT2VxKQ5U0h2Q7SWLiTZtTX70Poe+ZMMabQ+wbK6QXiT
1UBv+x8BvKVXrE3zOjyNUP/RXLiuGkwFFIm0POfBPCl89nG+e4Z3IA318RaUawLUhxbsDiUyA+NR
LOT8trgT9XuXYBmepfQ8DUVhIttZZq1pzelJCrYlsXMjCei0x9jqOAwyHj9faSE5s/OaiZWls4y3
Y9l8jdYyeHkoaqm3DhmTsU48avIxxD6KfHKLILtX9ts+wtM9m4LrlAZ1mFZ/UX33EcSeqaMXpTzR
GyzUkIeu2UrIXjURxIgXTAsKpT8+knyqfIisqnbkCOm8dyEixQA65PtE4Vfd8tIPDkYkQuS44SDr
lRsp24P9ciS557UysdW4g4RH0EOERtFTS5dIHu0f8gQ6z47UzwnMttVZArOVzO2uhBZZ0UR1FsVX
nAZpPdab7O+vySWtg5lRktdODMt+P1fY5ozBPR0rmTlBGkOsj2G6wpgaEYflQzG6LbzaE2saJv3j
0HyO4MC/gXU33knpM2ChNClJ+47V2HtmwyBCysXQberHa7VCaud9q3mZTTS9hHvAIhM5onFm7jvU
9Rzc2BCULQFYni/fjfGec71klO50qvj6i1FI+h6Pg+EcqmI3RTky9Fx6FEytRdnLwiy1bS8ksvSY
Qs0z4Uu+53AWVGKfxoTbg75KWqYJPxg+oshWD3XB47aWceOZSHMeV60Cl1RXkM8MP/adBqtHWsxn
xDzNkpModOJg7d/0exTYZwlcWLBjUoKk6zmqkak0db/KpJQt4rLRHFPn8BFF4CmQ/gZSQFFLbmoc
sTGEel53LlWDMBaBFSqpGIDBP7PUlk1p7BjLCoMNnsBRt7M5XLxm1Cgp0XyXDLqbbjjx9c/aqULX
SP4Comiiio96Xk/f+iuPFwPShxl/ENySRGThRLptUq0syq8wxiq0p6logoLcaRfZUgnVFAZpydcw
jwcyPOe57MQAl++XYuWj86bYtOyd09nmKxWoYNNX55qZUDgAXJYTkXHyaAYpONdy9UHkdXuTn3Tx
leHU0fEdICcrBTcfgNaLYGtY1XyXUdMORrB9mpKM9vy8NAb1BpUumjZxUFuANLF9EDVcl8AnWgzj
VGzHxDbxclk1/drd5uDJtHNjfZDUWrRNyEM5BmwbiWNVJw9FuJMjA2YwCrhrh02wBQv/xEV5TDlo
1UKB+50Myd4noi54dmhtM+FGjgYV25N+grZSZBmiHC8YqBW/3Y426z2axqmJUl48kEWqyn5k6ZhN
gYYaPe+WUKmB1P0MgXJE/8b9Ic7g1gpjyaFi5yvFwL96ok+9kq5rfC5EzGDTVfN0G0vgLANr8B9w
teO0HRX0VkfxJJ8T1AQivcvuWqPxy4V6tG0qA/KDL+RIp9JvZgRlOPyJ3hiEJSNo9RlPqCFt9Fq+
50dAL4I0PtKbRmHzvygWz8sCQXnGqJ34tSmvc3NZIhtmIbX+Mc+tA9VLfRu0zw0znK+bvr2SptPB
FWPv5eILVNP2xOhR4hHLMsgSlYfw2LZTG8YMeJHRovBmBsX6izVLh2DHmDuf+9Wz+aYNT9Gvc81D
NxIlzscBh34eMailwDDR4OIfKI4dzWePohA0BcQPkVz7Xx2SGCe7jbKOOJsxMDtNjIBkTkQ+LChP
yPiHIZGWjATaFahVSaOKsMzGjfQgy1qNdk733xRXBisHfEtWt7js3YOuQ679GJNZ1i5+PT9n47Hl
/n1zZME+RXVqF3rjQPmmuYFOWFnVXEvnahbkTnbuAuvRxkjMtxwQzhTblPpDXVCF0TfQ52weci+d
ie4WOnj+KahaC65lEH7cAc/X0sCaPIxgDaFvcZeyprP6GKpEmmX7BbavRBsSGYwLWYZr1eaMKjCS
FSpRnz8gC3mOGztHy2VMBnBxTwlzixE1ArixuYHGNOZlvk6g8XTCjDgNsE3IW9A4g4BpjPxc+EEF
tNtLWQTb+vwstcnsrRHFpwgorGuHV0CIZA9ztKjsYYRfKT82RQ1S8SkxDlU6OPDIupq26YQz8LkM
Y4ySRTwvdTpAUXpWhbTdfTKWt8j1RLGH8GJ+2SupFpo/Ek9WHiln8S83DdifUEgpejkNZvOZ8uul
1sP7j+u4JGikijio/fFuMn1/W1hUxS/TWrn2pCVQdW98mWrCc4qMcTJOp5RnTz9N8A4Ger4IGjYb
D1b4iO82Vl7mM/9XoPcRGhbHDbod4UAyBlIrwBjHDAjMCYJ65AfKboPGTUDD7KLfW9TLTZmb5LCq
J93V83giYuD5+yX77roO1x8oO7vpkpE4jhpjtHeMRcGVojB7KMQg2zFra7iiCLYbYrNqyPxTL9Bv
LVjiRSGJF854inaZXBsJLcgy4GUpBy+oNDEYK+no83wGWf2CUqIdxv811+30pk9gugLGthu9+gyK
ipCngdsHsLooeWi40IPM8HC4eVFQ3YOBKANGlGHn/Ra5GZ8uNNgo0/Rc97p8LT/iMRaFQdYm/Yin
YRjU8U06t2h48DavrWYwEF/r3dM1S/1S0HL/6BZflq0lo8Pyj+J559psv9FundGNr8J0VQXhCXmR
kCRlZ+SghakiwhKQgDHxKZnieV52BKKhm3xc4GnKtgQmXX0NIro2yyenQ9jw4JLq+i59JbiPmG8X
Dn/12sLoWhEpVUGiNWDbqgTL1B/DAn5zhSSfafiex3lpU7cCHH19tq2wJUs+rZhbqoa9Bx7giQNZ
SHtDuAoSwvkk8/f1jqvX/CVca7unWceBtqZFbwhq7GbeQw9O6/MHxGYscKFICyLh7QwT1VgjBf9G
gA+HsQ+mBdm1NpSUCx25FARnVXSRGIDJW3MgMmxkb9Slkd+ki+M/V0i7x054a9f2XHhI9tWF+hn9
7D060c82kRIHDHPB3xR04VcNCjIvIaCtfTFhQTxfvB25qFMEeW8YXkROzEvUqmGS6lBj0Ny8Ramm
6ufCPLHrKFlo/FZ4B5odKpGyLVmOvM48wwvy5N8oqDcRKCjQCftLG12NQCP2aLPZ3JWKu9TVd1JX
SrlkMAhtz99kzDIfXzIsQMBfD22Xf9tbsJuObEPOIxFUB3FG5ybIP0QZPpJIj89rZwvUyi090lLX
kBLjbIAivQUJccEZGFx+QBg4/777leMjZcb/BCUyDml9PBIifgJ3uC36bH+sVxPKPD5dcj883o2p
biBR0CSaamVa5rraigJLhNbQDc2lhCiSEM41WXow0Lxm5Ivw3weOrON5uQj3bpIxidbnxHX18Is3
R5IQAUaJm1g0ziyvBrdrBb1JdhV8xpMH5cHT2A0dLXkbUolOnfqDQ+FyApOMPEbMhL/rJUXruXc2
tSnuh69lPZPDJFdBTEPfIGU6K241njXq2wC+ZeqNP+PcFWJdspACeud/k0xB6NqkrXpdzso4FAxM
IlkrWQ88vHjs3LxHGylgdas4EctlhSjBa/o/m0jSYNbkdlIYuNd4P/9/nukhDsOb2cMsSD39Z19K
q4vTnuyY96fGr58hb8Mc17PmA+FYrbHhzIjoJiBmFvxvT5pxw1YE/3nBQkJZ/vCAFMzyWbVkUodj
wsR8xLwIylzgol+UR/vAFE4iilDW03/BN43Sd2eH43RSHfwVmIY/dKE4GIK0tl7nGfc5rclXQwKU
GsZQ1ZIFl3l9rJU4T6vLk/0i8uFsXbn7j/AQk7xbxbiYnuidt9fxIbUGIMMnULBIL6dZl/pn8LU5
BUXHz5l2F6xG/p3V9aXd7+fFchfc06+U/ZjH7UantLe9FG0EilqirgYzQ+Vcmf7W95WY6wuV5f6W
MN8OhxNLOMVfysnPklbGRZQ0qQK+DQez1R51HpVdtPnwr/J9h/KQ7xgAvrDHa2yo8cdwj3il0eXq
KU04/XL4uD+6OptcCjxT2zPpEaCFa3u+22TqS+YXFiv8/MlFRAzyxjYQgzVrp2ssxVGfwciCIrFO
pNj9BTS7kr4YKUGBbJGEhg2FhQ7GbzjeoDS6qb1mVk/euEF7SBwM9Mf9adKLLYIVRNLk2/Fqhuvt
jChedadNXrla+x5gCVf2mhEBud+UeiM2YpX8zLnoc0VnH3KaVL1NBDWoGqP43U44Top3MfaQA66f
RsicjSGNm9sh3ztUKn/onDQkFGlOBH6cUHq+9iXu+/9zkBVDwcWIoQhg/egNarqoxsUYDN6Jh4wD
RY6Tus07e6JlOzwhttZlak5VNtzH8Gd+vx14nND+2AKelwRbQsC9giAr/RP0wDalf3G6NCNInR2e
aVhsFF4k2j9IqTiNtMIP/aWtaQ2Bdv2iCGeyY8Smr4IeM8lGBZ2p40q7hBzrT1D/+5cJaYTcpKSB
lwQzBkHxdoeVy3ICU7FlCD883iRE/VPr/tu6Lc3SefdhiJ2yRx0YaN1oXjR0EQSAFLWNW5r7Nkds
Wzmm2MuFmTEi4WlbPsHw/K0mZUgcnPTHDQJC5XrFHlsEdFIEnaqM2RtRdxBXCApIpJ84zt3WW3lO
6LWVxd8wckiqnoNTSUKUAbntIwrL1UKNNrxAiI/sMSNoVmpsnjC9p49GMxY+P3zUHr7xPM+KXNbC
bObUZunlkl2RHxidbZArBpqVN+3fWVe1RtyQoaCYnsJMKOqXejHYFe32b+u3bZlli/dE7xbMPWa7
ccH0Ad0T9DcxLjeUoaemYF5xJC/CSNmmjCuc2teUpNXnlH0I86vex51VcFbo0Qb+13oigSQD8Xa+
pM9P0jZPh9Nwe8SmCE6bXn1pObE8k/XxynBiCYAZhUGdcxj/ljvgRFYFh2a1JlGgFqzblTYK36Rf
npRRLs+EWpBe1FyIO2cgOa2mztGhY93mSNYPjbSpG9el8Aags/nDSn6x89PDWn8sGpgmf/oaP187
O8KlHjCmA4L5kwpeC6ZegpjaBOGbRVs/w6lvBkDVCqh5kgJ6nwgUtdli0dM2GVSyvlJ7q3vxcahg
58nEWNqgUkgmntidhsLdVUrKTvbdw7tmUNonhzbIIL35teH5arHA9Rbn6zaS4D4H21bBxT+DPQvF
NVepnGMBAFjo0zDUePSjyv7A4mt0rM869EbEq/Bswt5Urjvjs9378Jn3zdCmB0PSt2x7eLTwqxSS
zPUdwCvlndgk04uLv8ZwEJ0nSYr9qiawmfk27xs+edH2kljxWqu58yDGUmbWnG8QmmGvcHpcV+9r
kI6sckP3/kiC2V0CU5rPjUc3ywfN/AbGxWdrSWhSo4hxx00vZ/mMzlJE8eJ16LHyQn70T1FhsQBc
TZm5bRQcLXUpCwqXi/fEZkQFedZsYIpVQqcLpWAGKamFBOKHZHkxu4RURVJ25DD/fCCZiZk5FKnM
xd/BZGIfnhuoE/eLG/4A31Ua5F+GK6rMZPBchU+hpkxWd3tchByNBC3c+eFc+UUYGt5nsvfsPUet
KFPPdLJ4f5pA4ahxsLXn1+6Dm0ufTptPvGgIvnOXmv6vBkhBKTkTYfO8+OVj/P/5CNUo+XJ/OweW
6VDudy9GqtM0Tr4oUm4CfznAHJcqDNqKqLAmEP3pPpCvpJXC+XWkylB0Ry1G0XYo768wLf5QXEwx
EpGJdPhF1WD2K+CHMVc2d8ccEKrO0kZsIAlMA9JJA4wjTZncJj87AkFYcBMG+ANH4a3Uj0ubayvf
1Exfc2ebUzQ+gEyPk1dPYUr1CuQe73VY8XwlTsJJBuFvx+agk8G6T0hevLg1Gmo9JojLqkSRLQcA
limpeXf7g5+75MyzFJ0YZ0OhCTJFSyAf6HNBojCHVPIi7Rgx50QFyXiYqz+YcEJ1RSeTGYk74lAE
NyzjCRNZddeCMSZMsBBD9OcXcuAc27z8YCRv/3Ie7QGcpEuNONq5SQNOQV/qtJsXgezsMEYPDUok
8j6FL3if72RA3zDEflLWvxg/yRCh9YR0VmfdruisbLJn4zHFK1kTjHsASPXTW3Xdgs92HmD9ojSQ
E23HePij71EvT71T1ELZilRJ1kWsK7VnQG0OFLdeE3oATgRzSyBh8TBGHpLmYRhcQbsjlId1OrOr
BR2RGVc7QoG9uwpUYSoIUUVV/hQkeTcS+38cHJn8RAFaJhnMCQOmXa+aXu+uzuL6Hewf6OQ2QXKT
eTiIY4y8EaHCzhwz0nn0aM/ueu9pnKxn5QKbCeQ3HiXChjpVGVPso/q5WSuYRlID2XvIFIZF6YAJ
q7S/goY7O5YxZwAz9C2pQpNxAKar3yiosYt1IA+nCi90OPykGmtdev5YZCIapF3ChX68w8dmDVcl
ImkByFMvHh0tld/TRpwz/D3SOV/fWJFnlBJQJS+TjfFmQBT/tNmatmHlQungSW0b14UNM3S1k9Bv
+x30ibEfkoUX6hMPWb4mRw3l4kX+oLayH9GUrp1ulZSX5Cs0V5iviM+WN9/WdC56ncPr6VIJ4bKn
20i4Mz4GqdEcXSeL2gaIlzvCPIC/2TXSGwAYPD4rUYH0NjayD25IjrgOfWBb16ZaOp6Il+UFve+J
p9F0kZBIqw961I/cXVQZMhEDd5mjABQzEI3quBZ4IaPqr4VYq6JPTASHaBdC7B5U+QK6AXSuiI7c
e7oGiiEQlq4KoM7kbAhbVy2zrJF+NZcJzwHY8KlRRtCPGAEjL3WeZ7enmU0c1bwwzRL5kHtYXoIR
vzwel9U9YJTKutvXkdcEg59s9f7XCdZS0nYfS58cNPP/vBNv6GxDwkDa9RDbRKFnx0YiCZB281mb
7DznjjUJe+WPQmL3V2RjDipZjh7VzLqBtq+X/JWk++fn+HkNFyioIP3EHQMjdt4tYgHqE/1Un/88
RA+j5XLtGbCNky+W/VDQFqN6EEihrqfXX9RmhD/ZxeIg2sHf/zKE3VfdckL4EeVxlibOun/yo24B
6ovlt4N0sD5+WccKLUu3t8T+XW9ewlhDcwyPl6YnC3eR0j+Ua9OsYgeeVEIewsIegdnUi6IHU1CP
LoW10nd2Q5t2/I5qQmffYYTO9pnqpCSPUp7/insyDGvjetNsrqpNrE2AkBZTjiJObZcKspP6/udg
+Hyiy0lga1SDbIDAu5qDPTH76MxkCWKnOuK0Wg5E9tC6dxgXlfJHNk8x0+1UYwt45TkT/+qi6uyD
+/ZJRrjM+q3zdlCZiNoOO3DXvqFcTEGa/Q3I1FBRzfSRK5NycDt46mJeya6WGD55U0lptbhUK4yt
Zo+RqCC/mXcl98NDFPQ2+W1TryEiOdKy52fQhorOkdc1uzGQUDBenBJctBJGkRE15ZpzGED075IP
wBDIZD018OAHVl9uAjqKqQJdcvwOi3+R12JE/Df8QH6QIabPPQnDd/8ZewcGKn1lSAOZNB9EiOdi
24/6VotfWJPHttpPxTQ642qrjYiETSSOPlGZF2jAPuzNYViTt9DIJb1dFPaeq0i+0mRsnb20b0Z1
qpH5N36nyGCgqmPTUhWpq0s1TgQDPdbHnd6Jx5aP+MVytg5cv8DRQOEy7preorEpkRFh0vmT3TPi
22e06H4Foeiv6sy83d0QA8HFmCdMfasIv9TKCgukSleI6+3tGRLNNpnadmH/J/d+/+2DhUNtFW0f
zhZF21wU7g9e1n+3mwOBBiY8UWuMg0/I4qkcYFl19ZdtX01U6vQGYeKOEdWddFnl8cWI5x9tpzYr
9wdawDz6J0vppAzE9GXxx3MfaipeJ1LLFhJc7qIhm21FbyGNm+svsU66DZVFqN/A/IIrisHynsaF
c/Ky6f1zxsHvtJV51WJV4su8ZQFfE3k0zJ+Omp8wsSou6zSr+Wk8Fi9RDbrj7assy5QCTckqUK8H
/qzMsCxoKp5xdRgsTUMtaGczOGSudeVWaXuuLiZbc2V9HESJnJBCVhpgWONnZSi441QsbpplQBZA
BluWsX0RHZ8AI7KoCff74LxBz5v1yf+J6T2Rde4ZT5M1MdJ+A2nM5ma36UJabqUJbwbancQQ82iI
CHSWLz29ZFvCvyG6FPy6vCFgWxsNv7ylSWS5etIPfGhRajnqTHLdWJe6Y1bGbi2kRa4dppwoPE55
IXruLMDBoUZr4Jnie0AOTC6JrmBs5iwtS2IryGHKRsLqof89V/40BczqP8tt+bgBNax91oMuKSMA
SVDmFf50/Oup/11DleNxvMSFANORvrz8DmVMeUZLybeefDt9be2Zjsq0NdV0B969vyausKd2gnTz
+j+Ht19c6ks7Fai7sPy2MMXc5K+izzodN9Jj6pnau9tJLeISayj+b0Fr2qtoW8XPy9SFx1ZTXwOI
FTL0fQIkdzT7eeKt2Fox0xSOzZ6e+5CVEAcXEs3NQpNxn+iPNaRujUs0CqHIxXgkA2HQKKpjuvyj
W2w0B49KVF6IAMp2mUGagAPNdQpPg5BRruR/VqItAH7r1Yp2zXjDx+o4+x3YqQdj0zAwQLaQ/pYS
ilVeWzqEyNn03zCBjOccqZQp4QA8VO7WXPPbjrynZ83VDe3wgTz62C0d/8Erjjiz2jFGIh3c6ytS
jng94FqGSnWtbih7yfcLojNfZI0TbNLJT3zC0CYMb+xAXZYG3zxRaDriA305uW0yR1kr+UYGlHna
mU605J0PShNtd/qPs2RVvHzFw3Zva+3jP7U4MZOjCubI0cBCDUhMH4LgdwLBtefN+AaPfc6DOjsu
ox9MCX+NP+aaIYhMOHT75tH4nRrsycdwTdSbPz4s30jVx4z3QaZj9dHMrAIEkfgGwY4JzB2WdkHv
3jekDVcMS1qZ7h+TGWvGDCiMJTX81ftOKuxbHMhSijpl+N19oQVq6l+ptxX2I28yfgdQAK6C0vXA
NkoEPIRdl2g5Spqq8icQtpiUQCeg8kd2B33fVL9yNp2JOfkGzSL+J5sujBo5jvvtdmBF/nVEUdWE
zqFZhNmgmpRLz84L8POnWHOChlSiPT84lthtF86cXZEQmq8/9wJnT5LXDc3BqP4F315vDoRl85zv
tnlqMKPvUYbrAJH60Dr7tb2f1d4O6osS+/abJdRIMQMq9pZgL3oBxjONpniDxO8mRMuD1gytGGJU
f28fcPRTDJaG519yp757mlutoEqV6Y5siN6w6/c9tTMD7y0JIg0xy8Tc5c/ZueytHa1pg0zzB4G2
U+2Bk9N6CyonJNVe3Mi3NwjHPwhJ8P74wHyZLcIxKk2dq921mgzuY7tSTZ1m+pDTUgVN975IeKPh
ppyztbjvwYHJ6TvZI9ROIpQBX16CJdWWfGwp1Nm9dr2lAqJrRmX6Z9cm9BMMCjJw4yFSNZ6v+g/b
4FKyeVXbTe5yYYIiQvC0vqgEXYRipK2yjO9Pn6uAnDLdkmlERHr2DYrHyFMJuUJllpKDVwdMB4HW
ouGr3F+FRxFyjqWixmKzSTbxs2ZWkw+mWUepqPgDBdjdciZE7obpizOMMniKonkDz8HRvJDLukrD
xnCtVzAsb3ws/jc2blw9gYRfiEysdcB1fmVxbxJbD6ICwjdbdH9+crrG1X4iuxQB5DWYVED7IKbM
xy3Q1WyNkbRo+9MMfRs4wh5MJ8vR7n9VsFUEwYAcaViq04AaUhz3M4Pypl1IaSg+IB8Nt+Fhehci
JxJBfQ5507e97X7b+j29sQyL0X33n1FQl6n3RH2EUF/H0vP/cM0hUKWIfPfKBZ5DZB9TGjMsB2oC
rASW1sWabxcAc9pCzi4Z9xXLjqU2Xnry/j80kZTBrNSqI8x/tUHt42dGi52Uop1wtfxq0zG3jKyn
hiRcLR8T9Ua7Y72hgBoseGE8zKxz9303fk/FK7A9Re7Ebt8Vc4XhkYji+ZWvdh015aahJFKh/E9u
kLUAO1wKGnk/c+lVqVUr3gtvNe9juIam4/svBeUBzg/Qw3ofcoaMqKlmOWijHrw2i2etLI0vLGTR
3mnBCePvtqXU0DZrDuio58p8L9Xm1yvGhJarRzhZwSN+QMCwtsccBC9JKXhZz3SP24O0dpPPIZke
qKtkjYUsEX8i+tZ3KFW8cKAgBZLyawxBYYHHoEBtIHWY8dUDH7gMVH6eXKf62wNrb0P7O2rziR1O
BrgvyPs6z30Jg/PaMdlv7ZP0aDS25Y0iMOSyr+BaVMRfjCqmUtepcqTz7jlWgE+qlGeLgrzdgvrw
XrZscZrG5yyWITshT9m+S1i/LaxaZU0Ob6oClYgD4X/m5ZHLm0tqk0srOQOp2t0iKVok3mIjbEb0
Wu35rLRvQYV5P1Qt0oxMBcYLr/RwyP4tV/1wAuVgPt2flvnt2snubAU7CY/3rbpUu7o41NWfRSln
zxQJlb48vd/Uusq+Dasd9gwZclQpEmE2/wIM3S4YSb1GXvgcr1J2/Wqj1hPM5kODevTDB2zAFhEd
RNAArChtXiK7o4jin+yrGwStqtICQrAYiejhnzdSOANXSpUQx/HhtUDFlFs1XCGwAGfryY0QolBE
6ccsoqiN2QttMirDA+qWEdZcAGs72I2Hp4xFNZfK76nUGnFviP1hhNtzkaHeoA++Etc8Zgzn0ORG
oRE/K9IQ9QMH8iCQk6ghE4ABBD5CPQC2pzbI6wlr0VwzwaPvT5H82rzqZl/CpeaSpxBI7q5z9MFi
N7s+KF2sQAwyy6alY8UkNDsBwjfwOkHn8IEdJ8U3bkVtRACATxf+abkXiPAIWsrK2jHl/tKBEnNB
m9REX0WRwRtoIe73OJyCnqsKJTFbMd8E+A+pb6sT6Yno29nxtUxc/ELczC8vN4YbmHf64mVx9MVY
II8U6tMc32/+GYSk6L8+eQJe1fsJmA5yLIUF93XM0kcsPj8zNCpqpNF3uDxfDaCKAa0lkaF82sU8
9Rx1gz5q4gnOl119g3wFouUjg0vxHtoOpHmofXoLFoYQd677dBwzL/VUguRK5r3lNsvpSEpDuT/W
3+eOHrBtCc07Rw+E9gf6XmikQO5JWjOwOoGLtSanuFP7UTaDNMLBis9oQVAIqqc8ERa3VT47I780
eQ3JF+nlJ75Dt2OmQVoTcU/DBhwyH/Vpu3AM/XMPFgtEb0UDwqdf6A/mBwJkJmp4abGwuXi7KN5s
MGET4W72o0Pvz3A6nwU8KGRztWCSujJQQViius+WS0uiEGKweZhj3A9+UqoPqkSuO3JttqNELPem
Kh9ZuPLxDJIXr3jP1qPPvtEqrRXuBUM/3Xia6ruQ1pkI9lVntAlbrstJ2vdESMBvo+Fxsk9+pN8j
gEl9LUxaBC6ycZ/rnYs+r50Uiusdk29+Y6+b+aSD/apbnj1gKeyctUIb00GOYIamNUhN/4POQkTB
iW5rrsUddKDuwgLflVePCO6mvF2I5PRZX249irG3M2jAj0zGSbURbEoYH4AjassY4mHEFuddF9sJ
72kPvwJndldlOJNj3JCTnzfgRUMl3fz3U9Lj+oIjqQSqxTO6D1Hr1dFHKXfreunV84yII1Bi2mdU
aw0hFTr0XtrGta7OH/CN0acJHT2zSWhu6vYO53ZtTPYAncWBOudlWACs2xmzTuaN+y+AoE8yfoIm
hxDhar7cgZvNGfN2ShDSuNpcoa6uZRWqNAs0fQBCOCWHMeuC1eHIczZDXQHIEBy2ABkZHnknLKYp
EfOzYVYa0nXf+E3fZf2K+VyaNWztM6rRS5Onxd5WbuQ1eIWwo7P+4kfIwtw9o+dSX8KlIA2rfG0g
hRqB0FOtHVmeWUjJPsxzqOkGOE+76WS1LYhbFLVJg+0N6PJmyZVuEB0cqDlnC+st91SKBzt45W+W
L7IjJuj7O7fFSlFax+6Yg1v7N2C8pfi24V5Bhk3qdXQiA+TMXHHtlBNdK7/nfNOs/S3xcMl7B00e
qzplVeZQHKTRJnp4n0Gbe+fyNp5RzrAfS8YOXDWRo9mCugiZ8bRiKkktPqOUSiRZV8tuPwkQ9mVG
fKUVM0Hpnq1ieMlnCbhumXSsdm9VuPR71flnURfyIzCrgRAPkC08vfBygPzj2RaenQRXI/w/TJxF
k7IEm98eRsSp8c5kc2UtgzIbOuEUw7s45FBeb/KJ3n3yefSFSlG793UZa7FfBkMtLXIL/lY7OudE
BpkTvkfZasIHrOUK8rwuGIwllblWYx1kCyA0ZHwWTdbJ4IEu42GC+ctmSj1HkNpr35+EE8hmW1xf
ppUhnc7MoRtPh5o2lewbUVJe/G9HgtJSK+OBLceDV7/HLqjSTif+sLY/bVz9p0wJ4s+TJyXemXO/
5oAx407yu/fLtgepokFBeyUfqo+iZGvNFxlI2rVXY4hQINF9pZQpEtOwiVJ8bG+VwhDMOrbKlMOn
i3/iOja9WjLWlaoOKbl/cv7TsKQLE2GyTC5g0Jv2S4Y3NfGyzQVBIBUm8Ej/67j2SO1pdcJC5+NW
80xDhn6795z/XZbB8Zgnp2oUqAToPsgBlsT2wvCKYxRLN19u6qFLKivf4JSyyGl7xOErRIRNLkRE
vjVBzMoWrEIndM6L026AU3N2dqr/xNEh5XbfKNfcxjP5xVG0CdAj1gMa9AA5pqL2j/kvSIuRlb2f
x2QVIpitz9lBm+UiM2ENyvTIpyy2yxvuqxGGMFkqSS3ycmOohk3BiaUtmfgXY8xLRChwF0ZGnpjY
tawkJrn99/uhELMTY/G4NNAkW704koxAC40TEENwNQoqUzQXTNNX+EQ27pc8gbPZ+XSokJEZOyhQ
+ZkmB0MjKTDRjA3yv5+SfB24Wecrevr5VA4lJ8Jb3xjp3UZfBsj+NFOXVFBFSNzCJA1PIC6lWfdT
rbmRZwM5r5sb7K6h1HF+YwJ0S+aZxitUaTI/OXD2uKuI++MgOZMMU5U1SzK1BUriLZTCKykkOTCF
QGD3EAvT5zwDiR5CzxcPQMk9fkx/tOpRCpvn5HD8br3/4Pgnm3NUItGb2jIZCZ4SX90JOJB9nYTC
y4NCYxEmj/XfqPJFcI4aOQ0tu0x/4rRV+4ZIP47X1xgmS1rZJNtACX4Sb2y35lN4KkffJn01OHT8
s2Z9pJ0FoVXKYHWD0oNMgXrH4WwmO1uOMcOKxNgWXV4UQa5b8XBVN8I30joQvd5Eff6DZaDpBJhc
/VLM/+hhdExzrRaV+UwTgtssIjLEvBaOrBaKXIjHek+y5tOgoVm93YvOmXrCrv+QCGBwHJoesiaG
dMzgH71DT6t/da4mgRnmHBasfXwgXPa/Yq0o10afYDCc+6MmYQbJ37vaAqm9LaRuLXb8ReJhkxSa
/QJSvB4VgrkC/SDrsuyMxHfCJElDhVbX9irIw/Ka5gpvy1GfvFKhCa54ZdDHw5Mv7802FXXmUi/X
eisWR5GuzNyQ6dUxXTgEQ5+ybb5mAA5VJ+O1Nwxq5GffEOApKFfA/mqWVj0ThYugVXACWVJZBTzs
M+jmg6KNDNaTeubWAPC2QCanwh3IcoD+XvAaWvZghdz90vjU5O4t92n7QrS8ULgiRm1GzisGafDn
+/ghKXRwXqXbIJWkYRa2uhjqKhkAXO/nI5/uSX/kwediVrvg5qlydJrrGigcR2+VdAHXRzXi5Pl7
M2XeZ6DwWLw0R3y7wXg9vL0+LoaOALxq442xX+OS91rEQNfkRjt0JoHbGs2pE2dVF3dC7eSBHP+/
s3aD5xh1ebsZhs+dP7TobLA+utTRZPvUfTe8MZq0X4q/L9z+yz8W8s06l0Cf7PFn5vWcWrPOAsJq
wWBIdT96808mH163xrdRcGOsCwoJ/4aidAU5SOZVdlpxgbXpiexJ/4hoTrtY3qqxyrSqh2F+Rtnj
EGc12sIwJL0kG/wXqkGMoyDErqlBTD6tE2vOJVAlSzWE5a3sQ4j4LEPwTvD7PRY3mXb0B1lYcC5y
bV5Qat18Ox4zLEHrtWEd/OfSf4LcO9e8eQ0Q0lLR4uqZhn4ruRPyJWSLwdynjMTwN0zbfJLsRaSs
4e+FXoYb7O71G6ZvQmgE8BaOFuX561IcE2LwH6e9IOW0yN6xsLTBMtCZ2U+a6DrcpHzehPKSXU36
TtSD8G0j625JTffBGBphZPywozykkSYJ6cyjawol0CmXNlKNRAWeYqR/cuSOiZsmoi/KD5ckXfzm
oc92f0cSfSgGT6zixJXyU0PqW/8AF15V9t7CiKopJA1QCO/gW95x6l+yQ47IDhJAVKibloagHEzI
aVK8rQwf3hdZYNhZYcbQO54mSNklSc5qdfPuZbEUArco13etcC8jAJ6DD+FMUgd+8O827JEc9ybb
TgXuqMLhf6CQneNRCaHJl/z7EwKCS436dekUfn76r9E7xVmkf26unLK+Q+aiCAzazdhrNvuQhZCP
vk694U/YYmP73v8vcww7INSMz3MN+F1yyDggokcxvg9h2s6Kq/qg+RR+t/cwh/UcBC6dcYL4i20C
E8BrCIAD5+UclLdeHQiYmKuHEWVRpvpvrYHL5RcEnQGCJpDnEnjHSZGO58p6NuChi2d4x518fQ3G
dBlPIsJizgMHQwoEnZBZYIeMvnJNxBXRGDKAlf8UBRM0tCXu3NAVvdy2Xj3SiIuMOoVIHyvgrksD
rGqBvis/nNSKyDFNj8i1kucTwhXaKsAFmSbPx0O2fr/Xh0Vitie5FRtcv+2D+plaiQiXpx5rpQbp
Q1HbIJ1u8W+BeLsPTKiaiWaGkdC2GCOOCrlipjzKQzkOM6MaTFj27bCzA0MhxDnuf3TJGNGo2pFT
ufhW2VF8KaZ5hG+0X7QnyDZzrworDuJLhndDyLUxImqfD7CmDHZSMhOK0L7a+FjeoPl5hzIhQQLa
LBUjia3QyeNgLWQZp3ncayvoqs4USsR6YSMzJuBzopD7kjCpHSlsvJceSsJv5ZafRJ1yQkxUqgAL
zYyVnChJvhlF5Sxs/bcOa5RZ/2NIpRqzsmQGoDHllwIuaX0SZrzxKqZpg5EEhQwU2aR7h1NuEBch
vKF3VwiYw3ZgZLWf/EXrYxkpRmeQvdsM8g0RxXBXgLqVyl6aqSRQ1dqxnPnYVJka3euQfikDWxSd
PCuUCDEbMAABGur8txnETGU4AN0E36avf8DA2SATOplPRhZM+VqOQiGgWMh7pDHQS/aA8wi9ASYR
JQFIVWYZaYfNOmdD/fNPwU7J7JqrQsFsj961Uymp2Nr63RhYF3WwQQA95y9+NrC3X0q8ILv+WUli
S2N8nIqouC5s1NoeaWzuulIkV3P/iid5LauuuzsAyaLn3pxUeiN8UiPJQTD9HEgXMS5ie6RE2T7x
od1ycAGPPuAkUTBQ4/BIUeu0R/iZnqgO+yGR5+T5jQcQBnsEJz3q7tLnG4gmJB090eMLQc9pdvzB
2DJHu+YspnCvXYlkihTa1XJvNiuMgo1xK0F5fNMppMN7qqv11Mti2h/uDHh+ohk8G9HU8nEiVSVA
mW0/RlixqnStjM7muavMSVtsVyOgjaiB2VjDtdEl2Fq31u5WZaIk6NWXLMvR8OKNNmDgowAlAMtL
tfzi7w1Eos7eQstJ8gOKWtVPSxTEyUIlSHrl97GseoPYAouUJ7RwRAxOlkTw9ew+/RbwjWwTI6f+
zQ5/xwCPSypDQADaM6qUO+Ax+vpBj9GptfW1cT7/JK1iS7PZvcIYMMO/ZoJQybIVmWAF/7eltHWw
c7g8UO3nBHpJLVKmDrx40ZcbHcAzhk8KQy/MT1BB/6tlafwGWwdQ079Q8wGWcqmpbpSltGqlza+b
tIp7XOiVcMvn9SyvHBuhM1edZ/0i7bbKf/VFzwjx8rdSD8L3lGEVGTdz2hC2CP7qFUA6wz7WOil1
zbThhfLDZ4sFP/ajOrRd4ornL9KCW7PiEJjlwV60EqV+rvLVsHqmHfMvob38R8jU1NC0ekshFdwi
HwA8pA18gk4giy2gcB+MHd2uj7tNso4YFkSbh8Ii34v2+1gRwWsa1gitbm0B2y9LmkvlWe2qeRhQ
l/Y7cNQOQaSNjftd1ChO2q4hSVYngJ3EtJyl1LT3WeQPDk5052B2eT6aTgXctPqtRcf1DknXRqsE
v8OEktBdmz0IU6PbSd6X4zT+T1R8/y+FmPjC3MAXa+kMSpkC1G2+CNN8ZqoMH7ZAtlQJDOBmxujd
fky3gPrwuWkyLV7hbI2O37ou/LkJyC8LXn9zXU3jF43WYEyVelftx+qmn9wFH+krNWljnK+o/Ed3
qIs0gmZBc90fiSEHOhSKWjc3BuqZQM/ie0KAEOBn15SyRl99yVHQDn30Mt+tNzQ/RPauS/1rXwQW
WvxC4eJS28hWwKLVPCk2LeBBqUzSkaNrK8WJ0orK9A0caqdvYynK/nSOqFDGJJFeW+Q6sWXWpD78
b0ytQot5RthkzQVligKk5mLi5Vvcwqkd1uwI4YIUrxX84a8WdY/ger4jPhB2rQMQibn1JYwbmWrd
/bJod2cA+o0VzhWtCEeJZ5u/RlV990h3TyJ5zYYuRe3kzlP+/reasxocp5wfJjBw/m1Lm783/lOU
qODPeM5epqBnVGSHZwQbdgWOJ/E4a1N3wrtRfgXzA+9OCZf11npd3+bCsljAYJzWu9HTWoBpAPq0
l/WP9jp0P61jLW3BCgfGKApdemmbUXJQcwgjRYG2QJgu/Cqo0ilHRToL52upg+y312A15UlY5btV
o3n3TTpYT2ryORI6q64+eJW97EfyXfG6n6TGytPmL8E2NOWjjf0nxqCgFz7RZjhc0uJRX8HrSdzA
i5fN77PHArHpOHL2+mf6LEeH4A68JXEC0avoZyumWBNTKv0mvQKK7LR3kzxGIbFBPun1p54UwrCF
X54URrdlkq1DGGsG1fWwFyPrnQfYhrAPAET+g/3aPtq8BYYgnYYzVl1vUoDxLJbgr+b+0o5tIRbY
4ADt5hnbl9bF1hPs7ie0Jt7IeX5nIsG980Wh+cY++FHUe+4OlE11ytFcX3cc4KefAnT1FhbePV8s
HXIspbSFoXT9P8cNc5ITFaFe+4PuRtTAr7FNuRtbyKQqLkPLx27wZ5Hk58Qe+Gs8oT01BPSiBUjv
VWFjAkwND8PKDqDuG8zs40YTEDupGbA/gcQiuLq7DFNgjnhulTmXt+z5oZ1IcH869SJrpMGu3rzj
u5cOilonph+z+iV0bmXExuBIBN7D26yuD7ggn66EzRUbDezPsrf0163Aw+1+7tAywEXBgsWEH2nT
MrQ0VK9voTO1nU2vEfJ9/DwlmEIgzXgvkFmpg5aY9uMGaGbgLC/NiI7ZxcpTjeI9BcxISzqfW6Nu
1NifRohG4uHnLCu5E63ekv2ICsKPXRSLjNGLFnY86A+yaHr99ayIwPYLnE3vUpxLzXgCZyypuwIh
H1RkWPoKLFl+Dzxq2akGNsSWWriYqbR5ApUsIS0UBnaU4/zRpHUg9mUAgl13N03WZ2R2kVdNwAaP
XK7mXjayJYpKpcEfEuT7TWD3X3iP38uDgE/wh0Udku7OCGQG6Cp4e0+TuVUdTlZNSKkSHOWv8H4M
OpDLVzh4ll1BlivLKC8Yktgq09qb3EFhVFKdL7buBDuuZwJxsARkeC/KPMlY2vm5ULzfr5ON1dYp
S9HB8Zucjjy4wFM/6SbjrBtrWi+9W+jn7abeN1MCs8YyJHF3EEwHkng92Odc0dqxm8H7Iq+hTYBF
uiRYj1VtyW64JHc10aOPwDyb1aPOt379uYmVhNEgZn3JMxnZxEVvkaco0+Mj/rg6icWkflIh/lKB
UQz79TH5xiVf46hPHqdSMsxaWWrMcszeZqYY5cOPu1joAGRLvWDSLOM9gC3LruUbGWcSyxurl02m
eBv0doziYCDtrPLaomB5ZllKW8jcd1mqTgUAgtPoAzTvse8B7eNLq29w2GNLKnhzrPos/ZNbHyRR
rwSkpc6de2yE12WyWhMYpFV01KRuWYkSEL+MpR1apIWXhzhubz/2+si6Dpnce5VqwVdGpCd+z4ys
Fv931eBpUof2xyT82v17Crhplj+n5Qix4bMtg4qNM0+fE8q42wlVlMrrcYLsmhaGjpC2d37V1soh
VxMhqz83YAfC1TzDXXAS6rpOKPKqfi6HVcho49Y8EYxzccMXb/PhUH7ezbxTjAksgrQFnSY7jSlG
BxghWlEd477R0OaijFaMQfI72PzPqO2pM0snWRQ/CuAZ+4dz+TTrrkSyQNdBxQHLx3GeJlzaWK+J
+WY5nI4MCOA8G/NmIg0FgUbNgpEdDHEU+rkKCUgZbpfFWf+w3qqPBb0lUehox6bzs+ny/210gzfg
pLIl33ry4AqS73bBQWV9+u+U4gXYjM57ikIGBEr8hmuPs0/hG9xZBAxsdxU78uxyRK6saNdTKLzf
2do5qlWWVDDA3EGsbsa5z1YO+iifdUc+B2s6CDGNy4a1BDacxCjmA3HmxgRB7rOKBp8epUbwq34M
jVgMYY/riBQsxnHgvAJ8N/jTRsQpXC9uInhiEIHN0oVdg5MfS18TFEGMQ+T0Kxw6yX4uedCRUHnA
HaQ1xb5+9tLZcamBH75S7FnNAmu6OFyXmCXUjWyqR4L2JOT9RK2ktClJXbhcIwcMjtHBVt72XcVz
zYnQ0pVRxo52nkWuEmIHuA/82NsO8qkeKOtXFhA3FCssjPzQBOb3R8SUE+PPBYvmTwoqVLAPjutY
8WNymuCrEh3+alzq+sojNqGuJX7QH2ghFwDY1nQbKEbspdq+ey2Z/whoQaSfl9Xi+Jkg5aR3JVgc
VgL+V+fr8rXQCgPaXsGYKFdDagz2MdTnX7NIcR7MF1SM+gEH7LV0s2TWKiP/5MsU+K+M5Vnakw3K
tz3j4C8mzqrkgGMomo/1QOqZvQMnkl/5IqQSP5QIMJMfAz5g0xf6GJSnP4AUg2SnKB1YV9dQjQ8x
LaW9soytydYJmc0p2k9WSSkervsnlmIRGBIrPcM4B+s1DdVMmRRfd3LOeyu01iGXGAWiC+Lkfntt
KBGrdwDDVsrhOmjoqqZgxLZdYhAdDVMbMz+74VkE3NObRHlcjGXpyXZdQSrdJqK4b8qqImX4CWbC
+I4ZretiXo8pUXIdFvDCvYn4yzpsHxl503R1mzw0CufM7luXg/SxzFljEW9cClhv1IYTLQcV9Tyc
Ma2j5iNL3ZxIpF9W6wOKsE7bkHRFdYxHBLbkb9ovRoci9FqfPf/XKsu50SXGeZUsSjhVxyqfNIGc
JC9pW702QxAvvFkpnn5LWbD62QcODLDkJhw/i3txDjxG7PkmtD++ohrxE6fmwCovzHQKuTygghho
bggRixbGmbz0FVdjnL5d18Wn7n9Hwd6fGJjF0GJlzuMBD9GhSymQF41XTmSnk4bEtCbari906HJ6
hRfaWXCdL88UYs1Sy+xkje4E+V1eDvdxu1XWUORnGiaOS3n9eSy/CTkrBHMVFF4wx8BmXTp+Fr1w
5sFYIpM1NU7De8O6+0eqMI/IeOnRr7tRVF289fHNPle5UmYha2QrntEc0aDUPtE17iZ1EBe8keDY
PjGYCqiVEl288rRWPvPZjWHZ+KCU21yhXiqYj+5jGQsGEbQ8Nm1w8nTiaXVebBX94aaJPuQ04OJt
BSjd8ymNDe/TyoB83AkWjXEh/nrOb2SYnxNm/q/yJ4mA0JPNMhSpksjOT7DirrdUDCe3Xduwisl1
d3RC29om5GISx9eYlfRTZw7hVEDIv1ylOSImAyfC1ed2XSrvTXW5vLVV2E89QzF8RIaJjA/U1b8q
MBRNZh0Yw5MJbJFSNHjnwF3FgQ3D+lUdPZ5yX9XY9T+VsZOij47KfbaIPJiBw7hKTL9e4Qv/RSuG
2Ml3onvlxYmaX04xP+kFnzz/xHYTDXNOlKgfZc3v+HMLG9IYfIAfXUQ5zDdQ11xatTNh9ua2W10l
sLswi71mqZsbauumJyC9pBzK4qDydSyrSPNi+vMDS6X8/cCOhFE2W+Pf4SZs72cNiREWuSxbEGQJ
JntmhHEItxRkiAw9TovHNAL4aKVaKpGnA6BPFhYNtqHxSlJpkn9ddstLq4NEl5Q0/skmAeqMTali
G2iiXdjYmvnebCO97oaTijy/omppoRRpER4wCwPbQOBoGsSgZbkoMSHI/Bz0cC/TLrmyvZAfJUnI
+ytsVFvUhOXTuoJe+UsjYYo3bXIIr3z5c8Rdv8KvmruPhuFhdwJddYOG14eu9L6rJtL2JSBpwzE4
OtJ/bOBt5ciTECFqaYeMfHzg+nY3wuYA3MSfeEFipPaliXYpqVpTr/quCwVvx6ssFsZoF4AogYF5
LW3Qme4pE1VYnw6f279xKf0oLfUTSAXBQHUyDpDU0QPrXLZh2R8sXUCDnYz07jhBLmLMpqqS4QHK
kmjvtgT6gmcXCghDS/tiq5zkwKAdbiRlZdY0MB/h9iJ1aHzitEYFNoS3l0B5Xdo1jKrxPaM+f6+9
LnnUPkzFIDRGqs8TVHtdPFU7Z/1h1M0bb6pStE5gVUW7TLGOulJrqWy8Lhtlyb4dnALbnIcBR3AE
XnvXJmgaMzVpFiPDmKONMmhNkihSagVw6UbKIV9wk/VFnBL7wR+WRZ91i2mso0YUgWuCAv795oT6
2e/CdHkcrxsBVp82B+TZYIOVw/cijRZQHG1/F0wpmyN7TSQUt/u5bEYZn1hdqmg2l2EPgoFuFabr
QWtHyyYJ9q//tP7d3h2O+n3Knqv0L0sH3Oto+u0wDQE1qZWGLNZzFCnkFJr58DtsnzTNiZl84tNS
kLWcISfBXbl1yJ22ChLLeD5oVWO3UcAF7aqYJuLfBg92pUafAyXmzvDV36gR27nrP0WZKHWPgDoB
hu1X2EmVb4CXYowO+6aXokOfxu7JTeDXa9Pm3UjXnCOLRGzeFv6r9KFYOa40TZjV2Yu5rn+XYthc
KwfoCznxeW5aN1qxilIosWfKlBTwoea3R+ilalKBcTbze4Wc5Hx93q4t7HnTkrWfbVFceUeef65b
ZtVKfAR7oAhVf2zFOaWCs7qJFlMBaPWy/nwVGO8jrgruvaR/Qs5ySmcgipJ4Se9DkujHQMGBxhG5
sNLUvCHnC2ZyFwsmhcIUcTba62WJ3li3jg+zZxB6IB1K2qxDOw60K+KA53f1ZbakxeoEgNW5VNtm
/z1n93IVUPOEyOG15TJEo5zm4foqWTt3I8lGro82j5Qbaw/IyajmiNFKKBKNMT/mxLIlKINSfXl0
kCXfy4kvnn2UhBSO7iL6p2fZUgq8HxDue6mLKDlAve5NiGUSUO6S1FjqKz7CWi0NiK6UAPF24E24
+gjq1s4V3JeVtpSPDSyJafAR/YPFw0DKN6uS5xUGzbvqyQ5406CLqiv3Ah9Zf+IfJeNTALKo54js
ifWsUem9plYK/BiKmJMO7BlHN8fZtislz5Gwqyek4jteWzbZDc5O6goOALypRQEQCsJUsqBOGnCp
/t1lwlZmw3og6MRhv6htSp3RSqB0wNiTO9sGipb9/uPw5H/LrJcRWku0j6n/2rSCyfF3nnuvgAnO
FasVw1VJShsJ7lWqFtu8CiApbyb/tB9oQ7y+w4jpYREB1/Cvy0V2fcBOd+rICsU8ZCSuz5SMVyMy
EU5lzVNLsjL6UNCuRc5tio8jPBUmS9+7B1i1QdL5LKAfK07JmpZtmj+r9ihQx9CYvRpIC7Ld1L3Z
WWYJlDTGECZdVAIuuIleXGdOVtJxSw+I4fMHCwwVLdycJDEJ4ym03gV0jcZfG1NoMlvxPmqNZcGh
Tj9kcsGiC1hpKjnOhfJg5YkMd8mAL/8Cxu0pi+BhsJ3+XuCCs45H1sqwwC4rtrO9F6uACpmOxAV4
L9tg9BKSrGxP8JELyd+KOH2pUBKED4H7m/CduQbKc00lh3rBThfiB2xcxIaLpGMvXhp/AoUCBm4x
PBhX4tds6eISOcf3ujSCcvyZHMG2H84QhRbg9VRCyJzDRpc4GztAx5LJIkpZMrtflUr7152XWG3Y
8PwjOCHn3mmVoOSf6wTsUEVCagUsSwlVN11xsiU7hbbg/Kij8dZfeGF2umM7FlZkPMuccxH0eSeh
NbV3w/ManN3kKe3WwWR2ReBnOlDu1HXNtlplu3cMmFX9c4Vsq9Q6yDN8hH08R7Z7Qvq4nbyoYLQl
bVxrIFv9s4r0f20+4UGf8rQaj1Em49rScrNcQJ+48onrl3/nx5BoLOe2eucr/wCSEYDinopUIjxA
Pd3oX4Vic+V2Ul1x/A4eGAlrPoD+Os/gBdCOEAijY8qdLOVcekcQhpS46Z5OarPGiAcHC47HW4Xr
DxAUBZk3ZXmnMBzhPLUQ4/S00nlWGBjdFC8SXCS8BRpPiWbyWcO3Jd5TgFpTk8NSqh8B0fW2ip2m
NirHy4E2zNwdipEAkDrAKiE5ooElaF4l85bvc33eA1YUtDkcvjUI8agKLZ9lW1eJK/bCFPgrkILn
L+pzh1q9Ix6rd8nYwt+mQaxRtduGjgCXGRzl5JaFI7AhHU5sahVBEFMM/fIDa4CuapHCZ1epuwYK
lOzMdJxRIRzhSiYR1B0DAL06/UkEkH5nDIwWncNB9PUJ9Pt51RScdDMYok0VTLroMPrMWhan73xU
AIjK7SbJ2Fp+mdoFV1x8S5jBQkh+gosN6HZkj2eYCC7ZU0EfPbnuBZZQCEPgFnHMdvSch2CqGbtC
SUzcJf40m8QDY8McnKYXczogQezaLYIcKCIvpbMH9N75hbMNgleUqppqqNere4HRo9LD5+CvjiQd
rnsBDvuSOW54jN4zC6bs4di2WJCxTrM0EFrlUsPHPaoRf4hdKzs/tR1LwGSkPnEFmjBMfZM9rfeb
4Pwi9WABX8WPxjPDUtxKvJPwS8ZJoJa/1bGzIdEL5/AJxpU69QIvvbHDhXK3IfkOzBMowTWtBMpI
BnllQGfWbdasUYs0GIfha07M2UdVZg/UNLpVlqYSC89msnY5vyW4vBGSAs8f7jlPC1Cn+WIbqbS/
FEue9gLDdyaGu7dulgxlWm4TTcsc8tGdOhmoqugV9YgZGVvz8VYvZv8LufN3/OYUlMulrhvHwHvn
IIVzpVJHXRre9660CKqo/qvsgLTZYecVpatS3JLZErngV1TFRByOK3X7KDjfHQDi71FW2kzgk5Xe
Sq16j1EKlrn8SZLuLTbyKXMW2bZtdSqnyi0j+t4n3lI2NkwnshyzbrD3BskgO9ukBZWEoVRszWOV
C0VQNp5Q5YdnJeDgMhd006XN26Goa+Tl4/QTkAhlT4ADCutKP+nl0vl57uo5jKgRe83y6HiEKcBs
p4LcfGEIIHVX2ScSeCwW1k+cZsE50ncMxfi0AVrIv9tMc0xTdBJI6RAd7RDszmEkqlUI5hZMIfp0
FosPI3/4JDcKt+cB9Eq/39PlEFhuSUu2Befm7C4WkkV7s0smH+IIqGP5OmmoDGc7Njb+yvi8+8yU
4Z+07Mh8PrfehvzoU3YOzFugUsoF2/lreQdli7fLJ6hh425y4KEatLWQ1zSOwspfp07oy36WqaYW
M4QZ00gM0LEIu23AimEJj0Rs30Zca89RozHgYsSrc5kFf3nIUw5Lbzihah5+OMWv0i8NcFfS138R
86bpeuhpMTTF25JpXOTIIkGGgPl5LP1FAJ7FvDcAXgCUD0N7nsoJUQSQvtOAG2ClP9qlNJxu29/8
gp4xZUlhzGzZJqysqcLYUK1xc4HNPUYrjnxUGvGe++ZXSnFuusUFkmZ6atLJoXS595eI/gXdjnbK
bWPwMwTQ92Sf5kS4tOzQ0xh1meMOv3akTpZhyZObZwxmis2ylzrj3bnXfTveF1jMNJybWyalOg/H
u5OW7sd0Ssk4xdcXJD/s7FynfVGR7L/h9at13TyyJYvWgt+qiESStHDgGQkBB2L4diJsPBEFKxW2
adWzYCQQIS6W40vEs0G3trfzMfMygFZTqeh5w9G23/NnXOFCvA6Wr9PmP/BuKEpzlZvSJZaI9xMh
M/V/vUTdQ6IMjZvROd3bPhKiST2F3zQJ/x2uaKkmeolxIVGnDsKmcxmb+Dd6r/Ieekh5RvRfKuOO
7J3WJJiiYOsaQWr+4ygSLYktdkmltnHudaHZ4el5FWjSGJN6cSPp+41SxHZKpc/rU+U8wlYTtjNn
oBjZBvd57+eZkAA3L8+Xbe8w+tYEVD9Rbp31OFq+41yZyE7Nk199wCG7sVd9E1bq8jIB/IENy6vb
L8Q+iWZZSm8tpxnezxSFibFbKdvy2Qyrm9DgwA9xTTgPh99CAyMmRanF5gepVplMEH9OI2zDI/5R
ERa64w/HC7+Wfa897ArCSShdV+FRSapZeD6EmyLdEya6KZAObTEJzfcC1q2rVmhVctHhnwqK6GPB
jyxV4Xy9vvcIKp1WznJEARbTKWHHYxhST9VuTG7OBY2cCk7x03FHRhgDdbfMVpLUs6v646jIi9gC
bUlOf2ggC2nmmRUTncA98JmxohJdFEvEhLCe4C9Glk1AXl65C8S5J7i1iqfZ+EXXiSmbhxn6HHLL
AQ2km3a0sikXmDywR9ywnSwmq7VT42hOWDLnV0PoPlDBeigxE4bhm4llhi/Jhz+0+h7XfDolagZq
9QKUc1cBGcIE75gtwxPpoFVMXLR39zQSijbrls9tUnmM4IQuZgmLRTaEjFX4SBQhrhhO4NXoCln6
iBYkXYCrn7aD1stJAZ2L6IbY5QSvoDxrWTywCU0S5LlpwQwBUedFW35ZA46JpIoOVy+pujayIh+1
NTLgKEwL76/qlVfNKHhb/LipejoYN/izS2aIZY4htfihy1d8DS43H9im49BkHe5Bc1YLcYSEj06A
QxQLFYb4Nwn8EuZuZCD/FIFmqi7T5oFbP21dKaifd664oXZqm0GkZMX2BCJP7GcGKQcE5ygxkNC/
eur9jk9IaWszPZfO3reo6iEyLTtVzbiZmtMvYNlYBE0xYZ/bbJy71uR4PnvGnkJLbENoAApLT1gY
KC32su2W4UrfHWObBAPmxi64JH42JgTGMuJzgqn4dyqfJv8kTchddwNsxuwqkUSXsjb9Rathhj+z
zl266cLIpxr6bi+ZnPsZptGYsm+KFt073m9bZPnbC9rJ4Vv4uDQj2CH3g4HNe7jbkqDMlIjcJabh
GRJl+kwFCTcHuKYbuiFkGJzV3k15MG2mA9k5RrKCttrHykuTxtNPS7nMtMCbgcunmymhdWTDfoz6
0Xqagx/2T8hC20Y2YmviSApfJnHrUH4xUMDpozMStyleXUaTSX1PBEDRqQ4eXf8NjstqDrNOBzb0
K/VAHF8NfgYqfcC4/m03UC6pO2UrgN4hE2Cj55WlexVF1XM4D05TrsAyCaf39IGdGYSDJj86Hq4I
3mBquaa0JI8399SouqiMUB5mOo/DvkmPcZYdanUzlVP6B644WYSQf/4PpIghrMI3PiSAkqlTYcOW
2YvfXgTg4X/74PowDMnM1wM1pmjDDGRzUXjcaiFfADbNY4pPNroE9VfallV070aHMbgbd8xPM4Qg
C258Z6MpQIke8DKGVfD7g1jYYaMEkpOrzP9Ry821NaHOIrRtjcSQ30G9ntrT9H+IUH4aOxNNOgjZ
4/2qHS/dezgVAjCcUSCIkFpQEHQsCysfHMhl/j2OAwsW/FsohMOoG+3Q27jhivYEEGWSxEUeolZi
NMZ7CmgZE0Ce7AWY2i7vM04pH32N4k+2zwZrRNVDQ2rW+8WW4YGZQyyhsEqqEXH3fqa9+dQWbVYK
Gq3EnMsx/BnrVWS+LTXz8v2UZxpFmiTey+ZyhkUcvOkhBT4WFTrCDHSy7Q6vcfYpGUln+Cy2i3KI
bHRZPRhm6VyZdsKTl9Q58Wnd2e0R421LHPMaxjp0O5FplOQ1DBOgLHlxuHkaGBBCmgsioeOL54SK
1MDpGNSZpT1naQIeopv6UR7dIe6wkJTKBuXAi5hQ39XKIlZqoe9glH/+W0YIZCMDV6gIhkxtPTnQ
8rBVrxXwuiv9BdvDW5c3liU3SGlrViTOPtdFtQGEcg2QKANY0+dqAj2K3lwSftcTLAjCeCQTDORM
aPq3DxIcZzj1PJyf4S8ovBIMTJ7vOh2wzmkv7u9sAKK5QwlIXhZAAhjplmNVqZuuPNi/dIwn0k2s
Nt7iE0pHrqysDCp6kROZYVeUvUDzf2LIUtFFhVxJlMx9MQ/qs0hZ56m2jcG471c3pwkv+RTId4x9
92PUS+t2sKmd2vQaSG5i9rxtB/jZSelx40FSWpLyCqAsPc82ZBUKanOLmozq54ST5K3/4XBdDsxB
DYXWQ8Rv9fcjCniTt+m5okvv9+VH9r4aCE48ijhMycd71tROuAiT4XHJfvj6far9rxPp4s860tjG
amCweJANUpK0HlnEeZ1dIdIWjJbzwlHZfVgHf4GZ/lF8VqCSkcurx/eMsU3RoGogMmUVsxRXrvNp
QP0oZEbfQDme9iG4Z7sYX/XGF+3cHCE49GZ7JklV7Gd5vUrQne4F+vA55CaHeXcMaPb/FrWMnjkB
KeC3Ai8YQcrlK0jSm8aj9pFNk/G+3hbX2E2Juk5b2VwJTUZlr2bFHWUImQL0VTbid9NsYR/R3xzS
snnK9cT6MsWQFr5hyEYl9p52rMEgItZkMBluicTuUPLbHeGtA155VOt5EzyNZkjoQzrqc+L70b9Z
VQUfJOvqcgAaSIIofz0qLUP5BMaWjbzmfxF7Q9KE/nt1yGHrEO1+37ENy0dASUaA8/ur+aiQ9FIl
cU0mPY244l40uOeG3BG0V+v4kEOl4maERiiffyvfUONN5uJKat8z/ecbbXwoYDsoYWb5xB05RA0N
TIENYjN7IJWuayon/zIKrdU8mg2sCzS5UZCXulYiriPZSuuBrg5V9esR/lmKLbhwzmxPEc+9ekfu
Oayn5N1aLNOlFNteWQURqk+8Tp/xog7cr3ikeBazBEi2U97lF+5Csc0odxxVAe1p0T3F8u6MMkA9
q4R0hCvJHApWBiIBPG8lW0Ojq2zFo4DizbrbxjH5S9blzhuYwI3KnKYm9ex3Kl1uYeIHbq4o/gew
CrANolwY0B1fj0y9FUZX1O/t/XbWWNhvEZHu2T2dyb6VDPud42q9YL26uHI09R5ScIJfgK6RmiQs
ceWqtmSVB/MvqV9Ryya/C4C+J8Kf+O9GGIfZXmGLmAH+9amL0AS1LBO3iHfcYv40cqsqjlPFY1jj
WdF2mCYtJAhVc7wFWlZxGlEqhNujXTbKlSUL1OI6Q0Y7TAonSfyQX0hsZ0+TyBH9Y+9VTxpIx21b
pZeGjTfm8XM1WhFEuq3bd9VMpv7YXJ+OrRPd3ToRJYjLVkUhEGYmnjrpVjM4zmkrBT4dxLr3+765
zW1I/yE+G6Kk4PZD5qriAuUYhsG/s3PJ1QAHzm9ZOBN7yhbYmwCiAN96o8Uaek0vFBaeOE4bZkLp
Ylg1A3Y03J4jgX2JWPLBSFc1X5Ve8uSP+FFFaO9737nVjj7pPqiZwyWhO3KZewMh3jGztvRY255H
EisLwaXx8LzIpMU1AZxSRsmibGEXiwySGmWerQJ/r6dyPP+QsKttyPBXPaJS6ybZW+9tFI85yFTm
CdnQw3gB6rGRRV7DoXu0166HiVaQ+fR+bWZTvTj6uScfx2CgskadeOxLkvLsPYKqHFdd4iCzsHS6
jTGtyqnPUBH+LwQWBNo0VTqKJ3HQOWFa0gl8qUIzI7kEnmuR2l7BA/47NedVQbHElRn4KVA6y7f/
EOyK7QTQMhQi2zbegCpbVQnbE99xsgt3Z2n0AxxKV4Nmy5e2verAKxvJPPDKZpyphPDsMIX6InO3
+JEtmQS5jZ0pu97IjNvcG20OvHZqD2O+ZMa/0u0MaiJc/ftwAqBTHeNqoP6+NRpz0UfMyxnPKCiZ
ALX3uALdKxiA0R6b97NCXS7k8t3aryzcE5j2Tfi+tSrrtuPxL1N+uDwuyfoqGa3+0KpPHDhpCNW2
zDQXLMHkZ4AC29mQFJlriwiERrnHosE8W8IAFXJBvHvyg6Mp7YpvB9Qm9dtu9YWu9UO9A9gnuiHA
sLHpq6Sh7s8nkl5YdA+d3eTjLaRyl5LtXY9QB6xqFqgMwWPJbPIkYqY2KoVB6WMpixzEfuHnzmzH
yFBbhUZWSaYUbEltYKzysGZz9RjKZHp9Uv7xzZ5CYB4KSHWv8WQbM3/CrBMga5gEirDIPmYbtXku
PBbUKYsawIXYey5jk/xkcdW5DOwFe1BboO5IBLZWu9mwu8PXjux8kqtFz5wXttlWwronhyDKkrN+
6/u4+xLwiDF9CI/bEp18alL0Qy8CX+JP24fj5A3GXfHl6PD1WXw+pCB3dpyiCmdzHodAok5alaZx
WumD85ejSIj0D5YBvK9JLtP5AI9Q5F4fBN1+y61SlbDUwUCKypK558V5Nt6bMszKBdFlhZeNewzZ
08doNyJ0DfJ8HN8cYifVbXa9NJ+b/QzpX+SNLSOUduX8gXHd6zvgHWY2UimfoobRmCcGsiIOW4nb
aDKplPteMozQ4VPvfAoOJ+toNR3glE5Gz91W/OoWdl1RJdvkyvq8Rd8lDimYrml2q6QYOG1f5j/n
cz3WiWP646Bd0TjwqeEGM3gT4ieAIM4a/OV1T1y7dzQVhPVX35KluaaD5qnU/pwwU5obG1a+4SpC
GINpzonUS6ID8An1vgcH+xBRHxxAn0PrSYAPVcOzu+n/76C/kKA+mDwvh9hMBM9SWRnkRWMDf+97
pGXpCgMNEYuiDs8CUqt8LIV0fe7CULlJBcHOuuJx5suqC6CvAtxCwidDPvQumpMsqBXT6CbGNDHD
348w60h91lW3rZQYFxzSA/s7fzZrbTWvFy2asez/rbSAsMjA+llWvbhnPW9DjShMXFudKWurcxah
Go4MiIp6HO2dKd8ynMEzSX5ALl13b/8s5hTnPtWhw6pNeH5VMlkdbnfjWzvIRR8SvOAt/2wXyBB0
AW3+rzvhoflXm4QtbI7aCwh52I1AY8HJwvExDlGWeaQ44SSPu4ahLleGa/MjVnkXJXmdxwQodyqD
oMQoJ1+KdW9QtM0bgAkJkCBrJQsjTqCPflokBL5f+tpMRxkvEvNaHibuzXpzDRtA+C320wOTpdec
9MyZ+qkRN4OJBpGNYRqADxbbs5W137vxWRc8IgcIwU+mKs7ld56emslQBvAgNStnen8X7gKDqP4h
TUtQtU0KyOFNAafBVADtW75pcyTtOO96dD4+pRRj9PjWPEg/zTaImHSxdGJDpZD74Y2zBzMT7fJi
1o74pD5FtQ4sg2ZZ4DXrwr9Uw1b9B1BTaWCV0Mxh0r3E0HfBCrqVJTid6WAMLl5ix39+61qfRkYp
665rcwnMvWgOr8/WzZ4B/s1y7nyAcrmWQbC+NTKD3dbJtzz2H7UuB52H+U+GYX5mgLnBkOm5zAB6
qRyHRlWp73QxWKMpZZa/RkQ/wek+ME/i+DVMyzeNjdkdP/thp7I8pzUENEqVEzyS/HPyxT6q+1j5
zw8X3GjbwasHvvPLfeea9tQN2DEBJKNIXFfNKx25PcJ/u2yM8/MYVPxpAtjpXtywAYZfcr4rO2Cs
PFWNe0oZswPqa7ITKsuIAQRF6x0/XRm643PgJ5osZpMc9zPa9rYajek9re9Ex7bHoJpOEKUmIFgh
+mvL+3wipWG0KKDKIeV42fyPmBbAtD1I47IYduxJAOnrC7VivrbfvT3OBYUDh/w+2hKH11ogdNxn
JLjQ8KvgLyuFFqRMGi3hIjxJQxMe2bnTCAalqMr+Rw8cS3iMmmWFn/F578B7kwhcS6VM7rQIlCoV
hScnFFpR3vLrJoL6xNXg7Rd43d7x/X//6pgFAs4aaExtYqT0/e+IvjfJqeYCgegmAql0/Zy0RGfB
8vbl/6/eQclTAYt7SfztqHQngo6kc5A44O3tqiSSUuq9lr71Ot9elcdsK/loy8TtLpIbbsY90Z/l
vKRSCzsWJ4jHVHPKkaY18p+JJK/SacX9FBQb44S8ZJ5YireJ1YQG7MzhmsPSdii6uPQa09JP0brB
61uMZnK7dV5lMHNQ4QDdASJfHHPvUC9Rx011AQki78rTzrIL3jGyHq6Rz2eV8qMp28Tg0IPKD29t
xAJiJsGYomWIMkC88ndfBqhJMhZu+/jlxcfKopOwu5TB0YHtkbsSV+jKW8yqOxeeRlglQo5Bd7S7
7kKu7/TqEPfue/lrKuL5iB+IN3lLi2MgquD9nDxf3CHAZkDV3CdCQqkGD55JmZ57NL21VNe4oVNi
AJx6INVYkP71lLmgxcD7KSYtWW7V8YiHqXK6CtDa5tBk77DwokhddwNmOW6v49H7yb5LM15wnM9G
F2aBmxO0nP7mQSnjBg2jY36/oHEPy/D9eQrYnx1h6tQs17vDhCa4FrKjfzKmrS7e2ivlIDG082EU
veSvQe4NC8ByKDPtWzPiQ4igtcGnLbAUpcatzzTj/SqhGQ+mvcecchBk0N7ZrHjqcDujKIpYYLPl
sGwIaikIgsPA0EN1mF+bSLItDOao2Mj43wjNrIIGgYvru6oj7RrrusOO28MKJchQWXMavuTsO3KQ
+3WKuXKRzyo3jzeF+yEiDiXKJwte5Hqf/CKbN9aZeZHJp1hfXrS6Bd1YgTryg040D4Ygp8bjxCtP
zdo9rShADKI6wYEDS1J3xoIYhYZDHZqnGnW6v9EX44Xsvohhu3X0cJyWv/tuoDVoorPBiyi30zNw
VDSJNpCi4Ush57i9l63tc2Mda7+d7VUn0Ny+xwiSzJbQAf6PGURRSglQehgGmtqhv/4jnejHdwIX
DQioWKI9OEramuQBHHNmgq6JUenaLFpkANicnmXqpoiBQvNnJ4SSnT0z+FMdm/zV+RRNgljmp6+K
OzTzQU2tVeYWHr+hXmbiT+DXmZdM3IXGzPysB02NmPXGW5QyU1rVifx1//WasiWfxec763yopl1B
dn9eQ7saSMAB3QdHNfp5RnBzMGOEjYHEtdCXhqCb/Fete05I30544hBBEFuocmIMnKiHM0KI/JNH
5jH+Ib2bs6qJL9nL6iiqxt8UzQir0ttlBDmIxkodWUEkC7SfWZabH8EURXBeRS3LqLU5hUnMCGMl
9Gq7S+5EYOE/yiTsqxFkl8LKAvVbJmwD0ypsdze4lcvk/40pbiXgmovymI9dcWm9tWO3gu/wMgI+
4jGES/jRHQcaV0dC7xylE+FU3AI7oTGoWzvdrrkJFMDfjIC2TWME0BYKCzBl5urFyNsrGNkLYQCs
oK1MYIe0SLZBZbp3WjtmCOjS460qiwSLz4zwhdChWGhQwsw8fhR+uJ70ON9HDinLmCIjZMS/aPxO
IlR6p/qCD6Vl8wbzePijS9T2MIVYkmBKLQT0ev6esftOgiQ+aju5OMMW82I/Uht8kUCezqg3UTCf
AbVLjQX5p4QBdBkSEVXEyz62wlTdTwo2MEcTJYTd6DGcZeFtJWg2ZiK3OgPhn1tNpQtIZBmCi7uR
/nqVuGzBIWNuNmrYuU4IMzTigt2FNIY8FN2EkUnv+R18eRCO4H8JH4rjHxvY9Lk5sYkqqtVwOGr+
U9AU8/U4qUSoquMF7l5liDNXaEqt4J8h0B1fqGxUtilFBLd1y/0INmuGbJCTzPswtXcA8J2Ooe3/
zvgU9mTZjjXe2mQaTn2zqCi9uWOnnXYz9VR5pHxRWWqCaKeaAxc0FQ6hZ4zD0Sv4WOV0qK0OitIa
uevbAL96KNSxSVjqBh/fB1QICiGm7EAhfw+YVZueeesdBX9xu8kt8f8LNgiJ2hdtFHWDqoUtuupC
1DXRmCZQhIrxVw602cAQUWRaErcPjYxFto/gvzTsRWBVtoJ1lxDbIlPWcm8A3K5on+AcOicuhn0v
BtGrtyAeytVHuHrcOpKIpeP3mR6xrNBQQkQtQ/zeN6iJB5ApvCSVSh4wiPvWXBZzvwNmJMS5wt4D
YiePWNyGc8CYMV0hztk7O9q5PfyIAIg3Kb5yul5Jxn7UW0dcPcpvWbiGK0AB3sw2O1k2G9bygONo
HnU+yVmt2H/j8ZAMI4AeTQEzgwna8y+EbHBrsq97LtJTHMqIzY5dapxJsJHcttWw9W9jJSNx3J3W
/qtt2Mm2/mx6MMKlXqXCVwHk2YPwxTC82RdLYn16XMepqWHpPwNXzNX/Pzt7UK2Tz4MBLOosBn1S
R55gc16EaI7ztBuqPP8bXZrmiZC2GzcOop1SXgSv2pvh5X80CoxFTZ78OzKFUyLQ/SInKGEm50OI
YMvSIMXRtYcb5rthYjqDcU0/Yuc0j9Dd5ACquAfES41759Y3wE/0Yk31enYgC/vZja8wBslXlfdz
oMBW7rrKo+u1+azK7dKXjMP1U/GJ9RZWeoixLzak1CYWc83Yfol4Bn4GxKh9rTjK/YlW6QdWGsDx
jhz8Ou4ej5WCAgHkmoxYAJ01Upwq4SDGB2rbSH0ujG2bmI6WGvTam+ULCYcFv7rCwcVa/vtsLGIT
oNbKTKm9gz4YIc5O1H1mVskTIlkQq9OzpD2NqykBRveL16+TpMLMTaJ/ZdZeErNwH3Z2d2nyx0Lj
WFIj7yhdX6mFoW4/9I8MtittudFxFq1kgOe2QhyVgT9lrCmpQXGyGNnt1WTfOmTEedD3E4UjfGeZ
5cId7uGeYPdKUuTf8Yq5gm1PGLZD/87obTO8SGkO6f0dB+d1rsz5nsjFQZARIPjs64rIpWRDsSS4
YXWg+o5n23w6FZnk7LutVtoOHmSA19HmdLYrBCnGcOUJI47eRWhszSAIwPyaqS1n3IGdhvgOsxx6
QaJY6pLw8+fYJJdCEAVot0eAQoEAsx7H0CDv8z+WSk3SdY0541YwXmrQ7ZKqE6Ppy4zMjh75EOX3
fReP/uo8zVyHWh95FuV/DZfixE8/XznLUjFchYwpTSSq2DYvXQCC64hAxAYtOKHbgCvh6Ei+8WwD
wCCuECg4a5NDKYHyNv568z4TjTvnp2mw9T9flva5vAiYyyFR/F7GYpTehZivNJ1pYlGXawXedoHf
DHkKdxg6oGctms8Bu6XrAG0UkAjqw+dj8fb3ZasBRLCaAuKZvAklISDp4h7YBuHk7F4IyTfIipxr
byp7nD393MBtDUs1PSqHyLiAZkdpARZ+f67NkJO4Atf95D0pwjJ+JTn9UJq5oYHpgE7nZVE0wrFp
1uOIKMKkaZohOdklyIf75yqfj0FGwos235WZH6wKY6uikiMwBE+ZAFol9yggHP+HU+xBSHyV+pYQ
G7U5i8OTeaqBTmYjWT6UIQCCOKiG7SvKT1abJFP6WnMxc4AfJtGRDS3NgQak3nnEkmbRMvqbYw9C
sfAXRKFamxoYchVji4Py8nPuOcvC5XbzoEJEH6RtuLMO+HyNuBzn/UKWi8lhd+fr13VIb8cGNJ2+
0c8NL+bLtETVLue1sCfs7WNZxJaU4yts0jz5OwGOb85QCgyPC/ewa1rca4165ikkWXJhiwgYsOcj
kur3puWS6xHNvrpvfqR/EgPZUKLIczxg9E2ne5ZoAzDH33iuZRPJkhKzfm5zkYTLYsNozClGocTG
GWVvOwJI0tBuh3qlYim/EYU9lMzjPJZzgrmW+e5kOJx/YFOWh4UGWcj28u3S8+voVH0Z3HleO4wX
Catk1H65a21x82Aign0+OqlBRCtfhJmAmDtGhsxqLWcBFYghHuzPahPt1MJIDcCFLKWQXitvA+dl
DwaHlLKGwu+SunKK9q3/3gV9+hPuf+UqZdudBICbw3w28jmFg0yZEKqbrsl30g4A3GHpb5vriuAa
YiFLzj1ovGCXzjKMP2Mx2jM5W7D5NQR+tXe2NlOhR6KwyMIR6bdhQMGZ9kjHbYQOA0DeEurceoay
E88+RpwoxGQS6v1ucxgnoMNUzZqyQNNepO3wIxFln2VNJzm7xyL4pgg31mZ7qab7/L5m5Yahq7n+
oydG4mk11p5f+BXT5XU98ntGcqOVRJHDJHAzAwpIJqfHfkDcZ3iDYxYqSPyNsjdzvUC6S7vScvxj
dGxjAJAIAHgBoRwl96zpnwWDspsVgXMyimpQ/v+ZABHTJch5+YOC6hwV7w8B4wzVhEfy+K6CA3vA
+m6ypIRCq+6Hm8HyswBoMXJyHuC7obPdrGr8otIX9PTWVqMnFCblWBtBBM1fhYLC2fmYq13dGOlN
6d33b3eQx16if2lhR4VowLyYygAcDEt6RlNWpGl8BjEcOoKCp1f0NslZ9rQi5AaP9MUvEeq3Vu44
c39dGmu3lWgyk4FbkRia3dLwXSvSJKAKFGFSMzOnyZzBVShcEgG2VMC5GZ/5Lw623E5N/4AaOHeU
T51r4gZdtli6XOE0Ac89b5NsN3s8KgU6RyVcs3G2ghn6sv8E6S8Qjp8Ae02C0tUa7FKwcdFtGuGN
Q4qShBw1p5HEYCKVqrQCE4h/7iFssaAcVQw6Q3AJYh5qROk97Kn2M94j3+87dRW6v2KOYlbwAfsY
sAn2j/C/AWARQsyv7Z1rQyqIjLCYN8YrWe9WgmplfZY/XfXG7A89w+XzstesXVm0031f3po7PW4g
LZ8JZs42lOdILImAbXIiryhTf6Xm10D9EJ+jgrH7VzHbxhDoYLmmTSjxOhLYVKUr7AZOx/6e0Xcu
RX5lXOGcT0DlYyJIzXScCn8VpReE5oCwreHj5Njy5vFG+p6eD+/xYnBD3NxpDahltIm0T3STxV6N
79Y7fnm/OpRtQG9KeUE225iL6GM1+sK3NQFdmHRFeiSvH5Y20sqfvTwaO3or1qsCA4Vwax4lUXQV
CCwIPXCR28E+6CvzxVRxupt0oap+iX/u9GI44HhD7QrOpvpNCjcpjhBEF5I+r5u/IBFOY/QTvKjp
4acEuqecafqmqnmmLNghQIligoOxen2No9T8EqqMGSf2gVrNCVo8tO+ofsxjxPCZj+3JQl54S1gQ
kHC8H3ZmWTZRaaaArC6Mk6au95ewRgLk9IHs/fhVIhNLNfOid19tUTyNwPNpbhr6Y8tiyT5krAUG
ED1pBAbX037zll3ZOduF4J/J50nomc5zd1SfkkE3WihIrjr6nUPlXR5J2rMFSwOPiM2/MlM38dXQ
Tv7PQ3P0aavp1qS1sn7awRbqaIpD8oPZ+LhCGqjGE+3E4fse9LEYk1xVFO6b5cF90AyhClFG6oxx
4o3N9c564c+wfdVzGu7tzjhRqSHKTskxg+nQdvjmyEQrJnPQ9JWnn33yED53sZ9/BMk+LiVLyVts
YJ/MAYIJjoZoNCpw4pdy8MAaVl5rMV+XyOccsCMNbOxdKy1MMwSWPLCzsVfAB9mi3/qDBD73unWb
JZi7d/gEgAQOADPWsvGvij/zDIwRbLlnE3FOXyV2cLv0ZjZoHtc+qgWrPfU97pW+l+MdsXhPBptN
NP6Vbosbn1UzAQZYf1Jskn+bLXNUKwbXLviFAB+op3g+6zyJIkMUP/WpCKVBdSnDxEXl8eegBlM7
X7ghbKGmTZEEj+XKE+lk+pF6GRRn3EnTtOcAXWEfH+LsHzK9pYxJ2ZUVjqb0Tmrlz5V8MJ1kKd1H
T2pUZaT1BEvhfvq43Tfce6tMQzqHyuo4PzlozGvd1wiAu2kBFfyPJjIUMhKg/FzbIS61qjqH6HAo
nTxSafqKXM1jVAKXvxtfU1dkukgJVWR/rLHL3RToZpanRD0dMjT0Q4X9oNZjBdVgmMS1rANLoh0r
2T06ZTN+nBqlgx53JCix/U6KiH+LgyBcuw47+PaiBHRWQTNnYJTcBHEzGSPGjui8iuZflhNBhkd3
zScEnDu8KKBKjgIexK4MTqdqrViI9O1/ZpLw0M8R8kJykcpyzsac1YpQduBQNkCs0ON9+P+Qw+hN
C1xnwOk6BVJ3T4HcFST9E6Bok8Y4poUnJ4pw6o/i9K+q8Ets7BDi0TlPO1HyPTniMcwA565BB9D/
Ci4EAL2Ofg59U/r5zBrU7zQKMJIWgALPAxeYMlxZZCNYGlcn56kwCNGo1usysPRZlkQlP2lXlMUH
YDsn8BCPckGgwZyCiEswVyYL0TKUUWp1xvGH395+2FOxOT0nbZMJ2Io0OzclADoIIzEO17blLSZS
iNU8Hyw8WPVyu1HeGfp/VBhuiVMdZsbdLJAmohEYczBZc8PBdwmV51R6vVMwfWrALLdN4OxOiHB0
OhfnVSkLAr8gWfGwpfL+Cy5zm95IzgQtzt6cFGHQG1qXWw516i/eOrelYvIJ5BgCRwX9NiVHWtHU
fhQhvIkoZXEF8XwCCExJ0z/jJyVYWf/SkaZlaFI9WOPN5l2GdGG8TboGV/xT/MBFJIn3IRYT61uF
HCdWlcutXU1K0XyB7UmVMRdCwkgVxhZKtYMIgjrSGjRMkA9Nwy8QlEJiaGftN/LiL9Nqh4DXjPML
Z/q70TU4DyNjCEjQ2lsE8bczQFwqFs3F9uSS5VDsZCCyKmOPhLVNrdVHxC94C2gPJeEKsVfNjvSC
jA2vEURyKEbJzTAgvE5uvH060mjuBU8nK9iidMnB8R3MKjQFUww8TvYJeIPNZUIjRwRU6VSEOl3e
2gMDoPn0cN/+CGzHqIsc5lxX2oCdc1Hd+z+E7hoZhV4HjWzCPqEMXX8Kx+gUx9vnRhEUK6FwLq0V
dAhcvsTqzJ3MW8DXw6hUpvzJCo6fEtMbaYHRAU/1B9FF6dGfTfaFLcR33ZghFwQSyzf9/ClGM7+j
dgKT7a/a8G2QJXFYn+rqauozoTRjI9uvS+1qDrGaCWb8sZ+Djl/RVjdS/6m92TYuhyvuJtpBmyPq
EK0Ljbchna/MBFBmDA9tViN662ENK1aYss6RRsLeQyAwbdONIpSF+pQnL/EwPGkUT9TNCxR3gt4a
JUuP355Cut0FZHwjCrQE89LMJxhV0QnYpEKjHDuDQL7eO6+kHrFPLQKg9ib4+LsXtWaP4oEx1Wm6
UqpjvKp75c+diG18TidsDitjTEZcEgSdUiwchKSUQl1+QVd1GG3M2XMC5/w77T1ct61/H1AvmA4Q
duxP3ImVXubn4g3MMKVQRsA649g4OUO0OJyfxX0wVQWHdc8aX7yvW4Qfu6oDqvbwcCobt3HJix6c
VimvghyJQOTvEVTHFb8KzyeiM++JTVaBeYId02BsluGjfDv4/3z8w0ABpnQSJ4/zNqLqhz/aUvQI
SIrBGTDbBGh8EWJkE3YbgQzYoYSIPHpIHTdxjlxVne8iT4+tLGRRK+JbEWxZcReSe3AEvDOAk7LD
EnylxA/3V6ZPBwDqqPV1oVDI/x0/lBBJ1OB/yHBQv6lL2APoxQEaLQvpzua2+oBd2u2utUGc0hQK
ICaMkjiKyWH/dbh0qH+rTCrUDVXFTT8Oi6alVxhSHFiU5evRYaoAodDr3TJVxKMVK8klCgeuS3I8
kuBMrhKrCxSSH2PuvI0JRkZdi9NupMvH+IsnIQkWU7dNoqsmZsypiTYWpaPR3/23AtioHsTliPEu
i5QV1nC1zUnuQj63A0im9vH82hNBuQKzFyJxkRHsftBBfa5Z2ezy9iGJD0cccXUw9RCClAZZaQSw
9DklXIOv18NXots2b7xlGj8IzTgBrYHIALj4uUSLl6F6JNy3blS5P+TkyiFDlwaAkCO5Rvn18TJ0
wrRj29mGvz6WLh2BlWQ/Tsq9TwlmE7fckBe2qtiBpSVBmBNnrGBLv1SW3IBUhTpamwx7rhoOJQpA
Vy+WuRdLMrPgEO3EXnbeUCbWGdT4DfJWSIckD/HhwxLuR/a+ANeAZApQ+7U0t8cfhNoaKZdZ7ZNX
iOxJZbeCILzw1I/UfAC9OwGGrHG6Z5mHAH+QsBtE3mb/IaNTXUQIW3lJ41IEMxW1YYXbrCXSRCLb
pe3IHAnki8DXpJ+5N6Nx6dsUXlsrjTXpVswOMjXUk+JJY66ny01W8OcE0fWIJMohm7VqFOFy5N8f
DpIHvFQXgDwWANDn01nvT7f+Hg1UFSeceYeVCQmPFOrwXfHMc++3230ABma4b5pYB+Ni5XvgiIgf
MMh39tmP4/WUmkVDoR4F+ikiLv5S9qj3iw7d2iakfDFWgGSSOX/iXMEhxwZ4iPxSro4ogXXnFWGz
9EHC5TCy4Li4sfQkMN+eYduEiGebyQUhGYG1kuoSA1yw/41Xg92RZ22AILxtZsPD1G9M1W9lnpi2
pl+qFeujGZmJMxAHfBxPnZyO9uPjfndBkUPyLSgs64TslhoITKbMjrKJWjCOwMl/prVHjtMVNv0v
mD2qVXz14Isj3fZXbR/KCzkee0UQcrlCyzVf3tC2e2lSUk1Ra4fdnI7VdrgEdvouXK/TToXeO6gi
SPzHKWmh4Lezo5dQSZsEBtS9e6VHfezc+aPfmF6qaOdo8YLrVm1O0faxDqRTICuOnh/cRtWhR8rE
A9Yj5zoAZ22zY/9iJXGdcRA+HK+j04B3uRNvFoALxTyjuDbbYdyc5taRpoyaPbvvkPt4FcWuyZz6
LuzCOyV2Ivf0xQqSesilCV2BTDD29YR/irClBUEuA4eyY7QXQQpF/AvjJjfGTnlyUKfAK01s5DTf
F6VrSvh2Py6IcHoOpOLltcaZ/ZZl0sThi5PzhR0d0jz6F3yW9oK93KCXVvdVQgteqQVU5L3AOyKx
Po3LVGmkYV/2uxBW6c99WYYm1ak+Gj+p1FiM0DJ/QX6s4qmVtUWgS8ayhO35RAcca2t6+xWU+R+k
vgN/GP4w4oSAFMHtGFEP/iL+X6xSPBWq3Ae+tVhvYmxgPZ83RgXacQZAGTj3+olJmR3sp2FDSpWB
7eafLwWkQoYw0cvlxP2LSb9+X6WmhJYIpRSnj98MJgxmbahnpW190xeo5s/1gUreN64wMzMfZjE5
bfFhuCNOyuhDd1jmJPkexviHV+hLM1CWSwsMz4IdHbaDuzicg2nMHrakNRN3T/Jltn+cGQss5Ppw
S5Wx4vVjd/PAIDklVlQW4Ztu7voSDjFizM9oSKH3a+BjMjq9SAIsTm2BCjHM3GhXtAlUyO1LW+20
0ah+v2o5PT16NFwg2uSku7KAsJzD93hTa9/itQpqnoybEXmq5C9VRhK6n4/11GCZd/L4xj0wfwGo
v1x3h3q132Y/mkoDBvBcccLlXcdDTuznD3c98uvRBneaW5krPgsMMi+7bkreKEe7/8bxHbiYYJnU
8oLgw3CcUl4FqAC/Ngp1CNoV94b36WK2NfVvC2ueyG8LRTb7bx+0iuz7WUa16Fj4jaGCEwySDG3E
dGr/CDU5EzP1nSanopeJzjeEn+xgvWww6eTkOzodQrOVQ77gKt+t8dEbTsIV/0tQ32xNcUS6LLOU
fH0YpezXw2DfbNrPBOb4fT6cNvCdbEl3izTAN2RpYKLp2WssJ8p4YrH6Ki/Tr/xJwmu6W/fJ31i0
48QEoNXolAy4uW67166dJd3weqkGeE04q5+4323NISqCtHFDFdZz//9fmKsoGKxnu3UAbaTK9re+
oTNp7rZ/IuMwrS6QbOPIENOO42r+VL/v5AIFWFsgxe+A2WvohBAHG7pdpTqW/NKnu0A0VJDre2mz
m3rN2x/7HYyG57UOKUgf1YJlLAj55pWDji+Oml4PAl4HGFtGK2vmHYrIkohVZZBXQeHomGIF0QAU
xRrB0IZAZSa+O396YQBYO2nx0T0CoiMZ9Rgp1JxtXtFsYN5VoRDdYujkN4Pk5RqQRd0AHDG8gD1h
zyvonAm9iMui3DGU1QEb1HKEjIAkEkk2S8GB91kIlCvd0ncI7NtigCNlUdI4+Ovnwe5/WecXJ6eZ
UuUuy96P7YsgQwa85XP5O8R2+djQLIGhoKBJH8q2ibyoatY9JGPIy76bcOZ8UjfQYQBv6fp6Gqrz
cgMWfwtnSJArPgzsc6JHFSxdxJJbPaRc73s+piRFb5wg6BvaObQAkBwYdO1gtWfCXLjgE/rY/ApX
9+dMlmVH80TkyX9nexGl9grLRYxzwEELQx14jy2FLL/zRQoXimF2WFvD3g6EErmkc83ihQ0bqyhJ
5b/1UVlL4wawSCbTbD+NdUPeMlwUGjAVE9vq2sTcLJMU7C/cOkw/V6Ur8IqDOdMnTYBIPEP/AoxM
ajDZchzxuU7YlhvVZ4PJlSqYvSWg1lK7yzWeXCfv7RIAO6rvAKhtFAnfYd0gyp3uGmPoXNdH9xFi
ApyKsFcvxipNYMnEMKv+sHNRNTPmVAfWna1+nI+9ez6K0tX20zH8eTYfFfc1lVNKC7/K2L0le9yI
x9qiQXxmT+Y5OLGnEkseX4Lmia79/vCh4RmKSpE32jI28wft7ltTSRgja/x2xJXh/g7jompCjSAX
it0co0dfN7gV3fP2jC3P3SogfpwEypYp+oex8UmF/f5DOM5ScgFpV0Fh4xyN0ClkWq+HELVnJj7H
WifV6p5wBIvK5lfJ5s5s5dvf1vlnH5NUF/GyqH2lENmqnQMi6nshWszyYNTGhZ2Vkt/lJzKV2RXu
aIYnMh9Akl+His4Cr3sbx1v8INgfaoMogmla4fzqhef0XmuBrcQHC0+2XSQE6I5m27s1oERjQI06
MUVsBPrrWhdRZxzIn12IwGgMsXPkPmnk9PCi2F8c85R2VjNFjG5XHkD12y9QG9MXhCAyXqoXlIXL
bxCNYzg75o6FzifVn1R92HXKspybLi6NNdYNrx2yVJ5mvI4Odl89Qg5Qj2k/rwQliXqOAQhEE90p
ow+4gJyl3p1gLghl6nVy51gX0N/ScLU0Q+MMkE+Z5G9yJWrbM54vBJwKG51VQkvIZQ9O1YONzBA/
834AehUB8QD/z3zok90GZKoCcCNb9+n2Hcx5X3iYUfqgue/8tsu9FXvleaCs7zplvsYFnx9CRuJV
lzVsMCbT2oID608Tn9rSQgiEljz0sp1w6DE+Vy0ffmCDxZ8rULKJ/2PDTUrV6HDvxUEKYvcd9bHE
6Zk1Aa2dPt0Zw2iaWOsV9snfj1ATfHrAB0goUxFtzCUqNJGWTmT0BpM9I6l4bx/W5ObJOovpa0h7
T3TI9FSD6hhSGC1JTMvBwsd5US9SvqBxxdYhFfTK59GS5vcT0aozzbNH20stzKonKuAaKr8eABKy
AD3oeon6BSE9cT8XBrusLc0wqHmGJkqeh64XIkZWJFwUFHY7Sk/uy8UiTMAX5op/Gi6TKa1q+4XM
3aldtP3Vv9r3XBqcHe8+ffKo2xYpkUN3PhUPRmG3VM8ggmklJB9N7O1ORfe5QUIOZ7dHibM8OuSK
fnrVRlFslwBMNv3UJs+IXSH3xRIgOEdv6+U38xuTEsYzGCR4KpWrx4wyy3KCqArEi/Fwn/x5ez0W
2p9Vt9b/PnkE16ql6bvxlgypwxgSrJSQk1cLRwQ5iuJNyfHBymS01o85NDkgrgnWyGh5RXs/CiCC
U+O7Or5t7gY5gyQ0ZViaKR5JsW2WQfdBG2ABpkAB8c/dRg3ZPhXuohzhqZhSHmVsT63och5nKsHR
IHkxuMjD9HDnzICX3gXkLr0UVMOvkmYpKLUfvtuAN2LlOrwkai5f/zaukItvY5nsX+i+UfxvDk7l
cuRb8zd81SeOjw+Mmr2RpY+VBJwBLsDGlwlO8CPP10gMDj7DUbj0gkLZfbHku20fgqfi+PKZTIHb
tq7le/CuOxsufcpQnsMxrGxyijJJHYRz3weDsv7Ll+kD2xuVnlx5J4jCcYPBwC8R86t5pWg3u12U
CtNxxAZIMv6sAAOF1nBP5mHe4x41kCLOMNW9EpE9N0HdAy7Rg46WFjnngUERKxq8S6Fs64GrFvZO
mm0H6xdsNkx7tG02uVcZurau6+TGo9MQNHJrpTZoXym1GibtNh9rDFJFQr5EIwXYkZwMO/5y6miz
SNNqcpeAbWOh6PN0UhKgrW9aVH/pzuO5SmPRBKkNMCoutHQoqNSriayk/DUEDpX67p6wQY7Eqm0q
DF74hYA3WJnMBvNtPcGQCPnOFppTVQPLSL5+vEoEeConjaons3hCUaChtxkn+m8CCiKl1ao+RgTk
6Vwla9+HoIQfjuClV28KEjpXoFG4ppD3ZkYJyadB04/0VxqikJ7DZYq4PlN92V16e2Uk24SqJPFQ
SEx+DPbNTI27vq3AbcOuVsudD3c1NbCE4MqCSLN8n00MHJAUL5vlaDIMllzc0dPtNmYabv77J1K4
Zje+fao83yJS/uqw59+q/D3xxtRS0r++c9E3zZIVNAsk/+J58RyzJHslvXNwsPaNGn15RZHhVr5C
jNFrFNQ1FnB29u/w8FKclNSrVu3pdvUJzkRLvfIT9QfkjhK21W3ZZiZ+T2we1Uvao2SYotiKeX8y
F2mVvlKXU3ydat4OP/mfNzxNBi6oqGujbIGRMdoN4ZJ2KC1eeVlyn4+xPEa1gFnUDSc1Qcp5Gya+
j+eIZNE1XDgxuJ1qhrWbh2szv4lqbm1TM9WCvkta8AdT0vWsudGQ+I8lBQtbzkHbs+7VASUbxInJ
wzV34FOFqWjtUrGYYtGYjxgWlKhy6uR3RzvZoyt9UiYnvX5pnDxqDYtDBMTD5Nal3okWpcYvl2ef
4GHh1g4W6tdb1ujJY7yCklnt3Gh6yMW0IGkOafw8tzkdswXtZdIzAaak3d3Ji/Rmw6ApIaX6acds
wgnYdmd00WqbtvFyKUFqQ76k6Oll6Vfcjdnxc+8DJy6hf+rgRbMcQQkS5DOFuQOENOGYfVZ5QwIK
59nnHxKSkN/jjhKsvBtBdGIXlrgejxC0lLsT3QwZ6+x1OidneiZswh62SP85KZNh/OyIfhaV9WVt
Vy0Bt9jk8EEvSSz2fZPuRU4K9uDFsajw80lBiX/13Uko4ep6/RcKSYEU7Rv7aHrUnX2zjnmFPrl4
HOwJgpZByFumClfDtwmkZvg5RLNivOpomqj9GRq/1IT3eXUFm3SBTeNCxnTBsVUZTSIIijIzjdc5
tL5WIeiPL23MXAmFJbBTQuT83vQ6LZMNj4iyn6AvFTM9HyDHXhzmL/Syszft26aQyNPfbtXnKaRm
Vof/yDymVuKtA6bb679qIow/uZs+FBt8nvv4detgVAj5Nj+Po8XDWJl/4fQcTpKDhHQu2ADftA4h
sxX73KtZI5spVE7mC7wqOHjKvGG/vmJnnGa1Qx9iO5mbT6v3WZmAWdiOyfrw3OrKUPAFs97RgGzp
VbjrY5uyHtEIih1vtanOJCs/CVCXQ4wj8//G+ozOKfbWX8BWBx80bxWpF77AH9/Ntb9RxrXBPCHn
TOoVPMoXBAqz03Q2mg/2Lf0I4Ifmqr2Jai3dtEihy7xxUbk2E0MwHu7sGM3k+vOWfoByboPBolwE
xD7E1972Fj79Qa6OfsE/7j0DrQU1qtAkEXqbD7Ko28miqTPdkm9y7np3dr3PQAQgivWzwkAfffTn
kTZKu6UjpEX9xT0ftFv6I8RUezjj4Kt2NDuOa8eQKkpoB3ylBwUpRQRgw5fLJqy23eIYBzMYqtjp
q0xjNtv5iRjMBJPNoQMA+Z3refq6gsaScHF8rIRki0zbjGQ3ECKlHiJ2PYscuZZ/Za5638DI/Xih
6aI+8herQhRV+XrNAX1Br7eWEntOF/ivQ82ShcBhs3RkhYqHWKSLhOiGB0VpwE9yKj3ApRpGns4w
yt5rXaxErS9OjorY5xDwAvmtF/fVOT/hWh8SAEIv867vDZPzjJMX5Nbyaz0899Z7vCIYfMo+k1U7
BQVS7sFMB3aJvAd86y4Xff7noJ1g3mkxCw6QFsqglDAfYhJjG/jHI+OqWODC1thxHWLYy4R9klGO
jc5rYa2WU0kexRYGw1B6luvQpAxSJ93xX+cSty7jZ6HaVZoRSLyZHxZsOPOG2c3cIaa7IDPyVhEk
qkC8RP7U54qGGx+5LmAzyaUwaB9GOwSs9hxYgY5TPAwuXAJkkI9CjO04iwqOk5nCtnxMA8yUH/ye
GCH0lP5wcmaoNdfRJrqS8vbjT56Qkvs7+Itu/Oxv1Ti54wU4K2MOdFYqpDgNRvqRxRadaOqED8SL
rsCkr+HoEbjS2bp/1b9KQtDfwvc67pD4bU4InEJODfGi6VhEiooXHkz3EEZgEqLq/L8jmoyMKvy1
ItkQ1OYB4x7vyfpLg9apnZThREQEzVwSlzu75qkyw89KIs7485oKdtSr+cIHvQa4iSubBy6C12xA
wf9jRiPG8v7JodwJ/vE062TrwlP/nrtXBUCLpGfcNHEmUaYTahjvmo1Z0zqGwsXV0ZEvYuogBFg9
Jox65kplf5Kyi2nsj+BRNwFVZKcmA6QtVvYJPcKU8UPd+I8qWsuNN6J/m4UWkcb+3j7HXcAO3fa4
JLTiAdj+IIBRYBF5M4xxXz2wDtF5y0wpSB6najC7RSojgpAk7Blzwbhq9G7fMW0deT1NDzAaSB65
XV06MSYgYv017lW54gx1GGOaxiN14dg6f7HpSNRPFRlbDvxLvX8x5XZ48tjJpX44csPzavWuKtak
XIw7aw3Lp98yV3STA3SREizM9zXOl0V9RybzZZflOiruC4XwYMKW60hqB24lvt6WYgAFVqlMzrf5
MKbJl5ykx5Mf78HdDWcqu8ynTderiWem+JQE+4dFBKo3v2TBJEMKzH9SKbwNkjpSPvI2pdsdtpGJ
UHaD11Pw4jFHUhuQAVO0vw/Ylr7Rt2wMcDfSE4pt27XSVtoMEVMpkShh2XBxiSvU396RrGDDQzD6
1K38Y4dPbH9VRL8egSmud/gY6kM1eziPDf6OjElvkMDm3txD4Iv7bp5j9gLhJ/Vq9eRQHec3d8V3
v561Wpm/OMK/VXAzCSeFnhL8KBeB6ofLHgzMwWpgO7CFzMBIo7IXckB1B3t58gzhQ7nX8esHBj6x
InUTLOch7ALXnnCyTDfwkaG+gbUIuegll7Jm5eReBjI1YI4SClU5xj2BlT4Hgt0qQPUGGJuF+NCK
NvWQqKPcGMl/CCWMjnA0MqUv9sBbSHwFZYZTbUbp0WPt80hE/c2h1Bqf01X3Fd8Xowa2VciNDszg
QvNv6x9fF7HcKhfr68pPrfc/lRiBDRQQbmD62YgMC3FCfmNXHjEgLZDGVuaSEfub8YuTy2M3oYGW
0UhSGdMGxS2SzQ4OAoJqKs551PZ00teDuv5AG6rdtGayAZ62jeYT4h8y2SWftPQn+Iff4D5I8Uw2
tRQ0xz425qnZgucJkw5RQDmwg+PsslKPZhPfybA3XaqXEkQkG+QDYfqd3e5i2l52Qyi598T5lA6M
L+n29scdDChqk4yNHCJJ6rEsoO8tkOBTa/mdHOXxy5glxkSQjeakSlyB2qyGA+dgG5TO54MjxRlk
nXTys3XxFvhZqr78HhZ5PtzoEnGddzxq4JuF7MewOwqMJ6AsBs7R+mG7QLmcajCnC1L4Z0SXeK+O
sPmN4LfYFzOGbbX51ZzX9uZ7Qgql5PdUQNF+qOPAWdG8YWdBCZirGsH178vN7yOh1Z0VLnW0rEvK
kdt4dzpqYNgWcsaEr/UGQNEXMAvgqpdnaZ0JEWQIGJL09WwHLZmVcLTyiL9sYCXIUD/hwCX1Le6Z
eoIqq85zOoMpYi1SP4JILgMBAjZKs0eZE7bwbXO/S4QiExQ2QgCN2TFd7oVp8J6oAMql5aJdYiaL
AueXHNBxm0HoGt650DcuELp8ovNJKwZnSMHdnol0yalYZXvi9Hie1Se7/PlKDA7Zw/09qgXmXnzr
B6lk2sOexFAQAUjHo5RXlm3tD4W6qFzS4YxQOwho6q/JEJ4wmYuVFlZlh+xbeMMIRAuivn88dAlB
kea/jldcG0iS/DUau8W7ITjyJKJlL3dqopVuMkvL2PjPf5aG3hGAKB7j5LrEmhy0T218beIYzIvB
tCWqUBy+bKOo+QqGpViIVGC/rZUhwoGjQgu+ApKvL5BC5kR4j4WYFBYhfWQuq/x4XLXOjozB+MjK
o1bxoyjmvaVckPRabNX03r0LhVbleLLRtVlDlWql+aTsnVShAaepHSJdtALXZnV+a7leLhe4DjvH
YVXFEK8wyK1QeX79c0F4mJYq3U5VFo7ZaPHv5230Pm24EDz4HHw/+bwjsPhamLAVHFxBNtJ61mx9
YNvv3PjIME5vpi1bTKoXolUOJNbhmwIPu+/lV1xVT4NVRDv4Mhfn94B+wRvudeFiDvd1QcEApeRu
hRYAdNYI7UxGFJDTL61B+3oTcu29SlTWsDKYSlZWBACdVwr3CjRASPTS+aByTgjnrhgkRzR0Swek
SsieIe7sWJPhSi5zSocEhj7tfX4GNs85X+/KNQa4KlIG0bX/Krm5+4h7LpQ2L4j8nvVoP5E8SAO9
NjznvQY/JhF37I+It77PHqCLgCT4PTxcDNx/W2nOPOaAwtFyLz7ETMeM0ETZWqtMg/WBU3oqF8+f
Cd8PJq0g4ATPzuwE4mZ2/0sf+pCwJQE+sRJkdur4iyeQ7IEP0q6Akb2A2pI2KNN7XbEZCnB7OSQc
UCiKErowC+Jrdb/R3J9XcjjmXUAvP+ZruOBfP84pv2TB4Pdlfb0Aw0tzqCna0085m9L+6RKhwvON
3jR9QmyEtyNwPjmnY0c7IaryLnMqTghWEc22b5XUF7xXLe9AAy+iqHL7FB8+0GBm6SVxifVeRxgl
gdgaqJyu1cfbaCf3qQXJGwMKa42a2NZALi+v8Dkuz238KC3ripnhewGiLL53ffDNL1QEnkbBBqfN
KgmSayprhl+0iIp3KjtJQQXdN1TOqosxBm6NwzyuInAGXseWCnMC3qgFIYd8Fbcbyuj0Z99EYqzj
jZbv7pJwRFxT6QbBF4jHo6Jj80r0B4nXBiDJRhlFx4Zq2O2Dh+Apfea2ph3SihgR0EtjV/DRYcdT
mAZ+yaylcNvvn0tPUbdzTK5dAxgh2doM/ncSuj35cPuUGw5RyscPXXvQ5Lef0Z9smtrkLaQH3iTE
exE0PSfLKnxdk12bLBEjgQe8Y06kxe9GGS0w+9hCVCDjD31LEvD/btIfMX2fR5tlv8b13bzE9Wkk
orguM+83lf23Fh492TxAMvdXWyl7e1/g6oZOgPabQCt5CSz26hfPdN/oEXjpnlnBG/u/Wni8Z+w+
rDs6aCWNCU/uzlu8Fsl7Cc78Fymj3YzQGOFVBDxrvP9ZMsZWDi5EPx9wXcZSl2OexNC6gnDSUudT
WT9u+fj7TK6DW2s/N13Ak2Uz7tzxYYzqgdeu23nse2H8fQl2m13DNDocJVbK/jBaUH2F1waG1K7O
v3EbmqLwsHO/x3FiJCArsfCyTmjuwhwX2DxknoIITEquIYRDWqgu1rAl/Jj0kiIldkBXA3eNo5MX
XE6TwmuETOcpwXMDAGxVGrKxPysbXHzrAxxugjnz2Z9TQuSWd308tDiHIvzN75vxvF6i0I2r4zin
YfP93xlM75C9l3CbJu5mjNC41ZQ48C3iA4TYSJB1Hq89vEtlmEBFJXjibm1ZXz4c9niM1+BALYc3
Qv7CbWj8o40Z9CeVR/IYQFDuz/9ePj1/tzJ/Z6ry49bsNpAAaXRgXJmj7nrv8fLnuzzr9g299fuU
It74jK3HHEP5ddfqNy1gyBVW4BKz1GfpT0BvjspKv1vkSs+y/yt4A0J7p7Fd5PfctbO92pOJVgBc
w4/ZQe9KCWbdAYiSgUxXNdi0bOZOpqQh4tQw1FNeNeYB9OYElQ1dWKSaDK9fZ6Q0nbbHkccWhvGv
uAtusvejWpDXnIULKTuw5Fc8x8A9Eea9V2hhhrZwNrMAe+1KxI4IhvSsFU2rEsGRknO3RbpBejd2
w7HcD0eKyOPcVf8l5moSh26BkyD3slXEKFGWB4z14xBjZRyAH5INbj9psdSn09dtQkH1Pa/IbeRK
fs/wkCVz2BvvI62e4rMwUYWsMtwcWb8gzMXM6sM/udLD1cHhcil37DVFjOwmhy7CBFUciPpnKDN6
4EMLxHTDqkd2KuqsoLxiwLiDi9cJH1Lv5wP3E2aVdqP0dW4tzzDu4DMKJFXDGKRaUzxKUi3LagQm
hNct79DHA4XwXXPG9/U/tpw2PH1xpnnhWJ/uL3u4VkuPXA64+ShIYn1tUy82NvKc1R67+yg67Ssk
1UKZgMRbWmZgbkWBTXlSZkN3H5tF+tZGZK6G8lRz7gjTsNWn5F9QgCvBPn1ZuFQN6hOo5RfUpREF
9MV08IM8KbNCQmE5zwK3K93unV+wMxxDddbRUpyNU0V5lVWNiWMfVhsMYd2x8pg5LCNP28omPb5s
exRGP4hl+RmDBE7rGXteGG2MWJKW+ZsNLGi4snEXcVgC1fIPBODLsWmRPP5XUzOYhYTfxnKWfnut
DrFVoZ+IKyCvaDFs3gXeH81hL7FEPJSkuQxsaTl7nNoKkhonwA7eni6uTQGBfjZCZKnkOo/zpDmM
UVpnQVoozPJDKIzzCnWEiXdGq3hlLfFbNd54xZ5ZBm4IkaV3fFtxFtxacTg7DD+7TgF4o1U3B+2G
QWr0b81sAObChhoSYtn9y8a9m+QouRZe8uBUEIstRyEcrilsRWiZR4buBxxJt8xajFCT60MEMjzW
NxQLfcGDPqRPz3qA4056mvWPVyMiqL3baNG/LbbnbiokgezQ7U3IvIDeiH79qt7FsQXnsxMh+TKH
c8/3D1VG87cojZht2GvQyuZNqFisb6kjr2QfgxcoqQn0D507RbBktYwts0/hiHViu7IJo95Vdj4c
Dalj0CH+6RzFtlYtcStU/7SeEK1BgZNDlvlI05RPprcPnh9EARRIcijkwB9ly2KuAFaTLTcU4Jp6
m0kwh2x2o40eJ2pTHA0v6TTFGjs0YWBzhe9vC0kkKFQ6b/Yk3BlMwmLl/czb7qKA1gEF8zYWuSV0
NXloArhPWkH6FUHvfLpxoIRLyYUBqr2Wsktu9AKtFZ6aqYx5xiOUwjBPSNgrjCLcnnSsYajpxJF+
SF450ifMUQ43oCqqSaYy/6Ilji0AGxXdOd2WO1vwsxUeGu4yPXTTinwscxJul7xutYwCNnezeLGL
UUgapcTQvx2AnPpCkVrgWZqRal5N2e1pyJhWs/4kVzUDi/i2mUSy+fS84Esdgmb9QId/7xK3jreb
gvCP3rCTWPgJp90OiYJCiKatjEuIiBK5USAOS05l2+ZyFB/OMPtLAfgR8T3JN/4Jt+2h/QbsxH2I
LVLpyYDM4gPNw9tLpn4RZc7Gf5VaAnF3wYrXhGPvxG23OF5CsPtd1i/4GTuWKSfefu3H9Wpup/pm
Fs5OAHiOl1D21tPI+OWfDjXywSd6Cr+m3hpI+Lb4KxepvgEX4Agna1Z7Ysktr+Qw6h+/V3l3pv5s
u9EikOX52JyjyDB5L3jdopgVY7fDi6DnvOqDPVGkUiNIyj7QWNUvgQjGwrZiyhKLRbZ+725OmMqp
pCz2ipw1w7+dduysaIrN2+42NbKgVEETd8EESGLUoh7XbZxKWsnSejjswmZtTPrLeavPKCsnQ2X3
s/kHm1ixybIAWGCKtYw9TTXNGDCn4kAf4FJj+m+7fRinDzomwxBuAc9467HjnD/lQtkLVczjZPoa
8cDeCRhbemNxTPtPtSs1D1BS+2tBVUHwBb2g3nOtaf8Mo1fnBqeWbbsZWvvhYsdCxU7LCbzQnjBJ
1eRW6GQdCX9L/fw9MvHgpNDzNrsdkeuflacsm3PumgtiyVn0WQTeVK97Q/rqoRFJNFhvrYWAigY0
31RtY2onkao7PnyJelY0kkKtAu0Y7XX6xhR+v+ji4NFGcTx3esxRoZbZkpirwoE8UiixYahHAFK5
0nlXP/cZYwWwa4jctlONy0GekEw6/sRvdQw6ryX461mSDET3t5mo/FUY+2yAvZU90Q3LNEucLVZ0
OdKYMemn71tMcta76QoiNK+Lrs43hNiJmb+EcPFXjP0Zpemn6cFATUE8u9NclgcDKM4Z9NQSD2lm
qS/dGOHGu/ANxxWf2kwYxnxaTtzyFCB6QmyU3K6slLirOTVUHlYTYenlwF2e9h4QGJsB+ZiGIFsF
ZbNO04QCG8nCWCrIk6y8FMDHYW8z5hA7x4iwKBm+XPTip618quGQh2VxREW7gLNqdMkJaGIC6fHC
yQ5EFWyKB7PwPSJ1gJTygHw8aGb3rWYMhX3CdRDlPu8rZfolrKkJAi1wLluw5GbfS3RWejFyCGqw
1mnHTS30vQsRTbrfFsuelGVDdylZCvorucmpK8yZ4gzhv/Y+ZijVf2nJNcfJ9v6K+l9a7zxk6CEo
8QPuB7wzFHQJ2J3eFVd/zfThYwe4i4HajOJ72r0zMj68gOOrbr5arYaOgfzN9Gwx6ke9a1cA+edq
/XAm7IQKIBf+TZrg+RtZ65qoYjs3/pR5wypjGZmL5pEJexQfGE5Q0XIgNQjRpoUPo9SCtRjLxoHY
suerX34GRVT/wqVTN5eW61UktI0H8VSQs9/+BxmHwrT9xfxpTAuTmkPUA+M0rKVHFl7jloKpDKme
no3Zks/6eMajfi2JmsIyzy0RroHz9OmnXcP8+c+N3tBUMuqnEIMsHApfwdWkcRlrYONVeh0NTBAK
fvmPZIsLmn2RGjPg2hBUWJ4+LdznGYOwm0q2d0V98ePHaTuq+H+7P99NAFrjulWG4Ghf5A6jBGbb
OGRJuWtulHHk9Z5pfNrspBtATrhcvQfBgJMJyAGLDKcXXgsHyW9tLKV1VUJcicecO4xxF3FWOVqL
ASO384Pp5rZ2Tv9/qHp+qaTUV5AugT8qBxxYpc6CpErHYEwC+YWweyhx6b9UkRGxt+BKRU6Q+Uto
r5zV65Y3y+K57dABr5AHz9Cp6FG29+kyea2qGin22DgckikfP60straUcKXueW48KSoblUf0HVll
BPXxUPcPMFRi2CwGkg0Tc5TFCh++i7JaORfzubVaOVAzyPYhMqJyJi+0WMoZV9UofYD0JlaVQMJB
RNXUbY1myh6toYvUs9c7wUk48DDQPmrN9Vavl0E9U4ksAxFfR1Xl+j8pBfQaM/JAEgp1jZb4N+nP
7a95iTQDD3y5bLPjAbNtDher7L8z+Fhu5jfjDQiA59DgFUYwQrT4vLbACu5hwpCXr6IFwI7PRv8X
pXxlbT1CNUOXj1VkpkHRfusjFf+ao6XFfgjn1579PCSgfXi8HQYVfRXBnCFoE8a7CD9Duz3iyogH
UT/uGfy3bMUhJ0ImeAZCGKE+qbszMjxK5ATK4dAhdlesYlhvMi/4fiptdB4rlwmffCSS63+kCHNm
1NnmLdZQUS7Ss0WKJ+pZcyn9SCvErPpdgHaVTsm9uwX1TWirbYNlr8KZVPihcHIZTC74tR7eEAR0
8IsHoCHbILDErOlQrnd3EDl07gT/G2TeJ+LdqzM9kBwDMoatomZTGW2dDv/ixSKyXv+jmcbUgBe8
WLALBZ/zpq3j3vLzXy4wIe3IrqqkhC0AzXuUqf1fre8A4ALO0ARysZXMlH/Chaj8Cs8ewqEtXugK
eTpQtX0ovY9bAVoP+uPdiCCK5IQl15F8iTM8UgGNsMtX2sbP95RTKtElh1QbdUv4b2US1pCxgsQ/
Pez34I2PaFh46nZCWJ0a2cH96BnT+mkPR1Tmzr//lf1/q6yB7KUEiWt27hSZOfAFu/0nBR1ZRxbh
JQotV8/nn+riVfMs0GXhfNIuWmM1A6vgzTNL6rEWE+tv7n/3HzbI1AsEfqTbUIRMBgdtwHLSpzXx
jQbs1Idynk/KbsfX+7axGVnQJvXcJhSZEuNXN3A4Ji+OoKzbU5ZZ3Lqe0llPPtpbFVjuvU7j5Qvk
ICpP0RYdhhuF+uT14tsRZN3a9sWmjhrJ2lekFVSUrDi261uwcUC4/YFNLEVfEhGyGj2AVtY/148h
GjsFmJjPJq2V57vQZJrqJYgOT8FRPHWCLCKW+ohS9Tayb7CetrLqTT7uxlbbT5j6cDltklrQ+O2k
eQYtd/vS6SeYjI5LsBvzYEYZ/uA0kIpmGwLlplHL9MSlAFEhQ2StH9ecaITBF7vYio84W7dCV1Gw
Bu0PYYQN3rTJAFiinYTEJ6PAiTblDl787ncMaSeiCVMGU+8Eh32bCu7G+NPHfuZuECcGVbdbWvTK
+U2v588Fk+F6dyBZQkIJmT/gmGj3BoeN1wRMSZyvXDKCckQdPZdbKZ6IEgejfN7faT8mVnqObrIp
8CADiyAzO2yxdgshLAZf3hG2my2cYtLdgYdGrevrfoEewT/tuB1075TU3YA7z/8nYOG0flQaZNKg
NdvX6aLitazsNkrG0lmdVMWGbmz6yWqHTEs1al1BybWgkV1opsOQf8y3ejtIoLI6QPzrtdRWj/jO
CefRQYsuAnW6SZsbwA29V57fN4J50M0UiDklfQPatGcfzaIMTHvrhjT1gHQmBshMAcBER+1jPZMh
LfaR6qaBKN79ivxZf7wHreCDxDQmj4Epo8qTKyC4IKbnHtJppIT6TA4+eC5ZEekcCKg9Mpgt+D8B
eYpGDPLFtahyGozuM5NUN4ijWiZV+1Gc7oDhhZXRnQ8ENUOQKuVsT6dskAvQMFSla+RnyqWLbzng
xN2VPLMti/zND1h3JgSKVBg3IHHuU/RpSCrr+DciwFDi4BWYIwZJPD/dljKbxHidPE41WlHnOl0E
qcQoSsryzN2jD78m0rWAjoI/mVotP8tTOugy4pSs8WV+ub5QGCVQSPw1dRM54MMmGVHTDLyYMUVB
lL2wgFC9KF8MedWtG8Gi7o8lXzyOzlDldQv4r5Izn6VGDs2qv7mwAP5VjES5jtn8+rToXGgSLMWY
+uguv9nYN6wSR4i6PGnh3RguWv9VS3fdeyuARoaUtxroA0yamb+6VODxA3LmRlvqibH7HjPzKSQj
eoR137/clxs8oNIC0F5tNRIrbuQxUxhsCIQYjBFF94/1MMd52xl3gx3ZA5oNAR7O+ab2LrFjNNGv
24j9RXvdrO0GAV46DKqsUtLF+rEyB8iP5mhD5jReKGn0tqiZeoN0StAlVHv32/Bo0Ney6XfIY3wD
YUFnI2vOekkoAlbBgjdWwWWkkvQkyiNPjkp271IMzOGgx5iS/kUeWgXx3ESMAA+1GeSM1TDEAUK7
JOhpHkDsSEz2cZ7qgkeW/EDe3zKpmdPt5fqkS4LPUQ05INTk2nVVnOG08064MIV5a9BpKvHgT3cw
a0z8mBVovKAXIqdXoy9sSkr7gh02eTzSibYBzYAwt8S6RTpBpW+RVcp+IHNdscWCbo1HH2SYK+g7
5O3yAbpHIU4lTU6UWF66Chcc0EUwUfFYcf/8CnliYEDBcWUDN5XdM/Pwz6XKqiEnGs8CU4MBGrL9
G/JHBrS3+eZKBmC3WwyqHoetiPgTgqdqU+oPLZzZkrkSGBnB2dCQR2TaMsLCcnr0v2TQhl34w87J
MZh9sTtuVbfsVDtrArHL96T4zARL1JU2nFBiGJsN+GQh3e4b3Rof052gPfoNsitpJmqz0t5qYspM
OO50HetT+UUYDEjQpBXo60j1Ku6hznXb6WUejYPV/qNy8BSr5qr4zpqx/FoI2yoV7e5SQK+xaBfj
j+o3EQNuQvgniqUR7v3P/8ESJKCQDSgSTnh/ucPeI6TSvvKj8ZgWvs0C7IIk8v3LkROItXGOvUnz
htQsrvqw2zRiaub3GfOusVyI4amoR3sQdUPbCOw76/wjaU8VLRaAOnLzMnXOJaroGRBalmo6+Ju4
jZP5WRM9vNDcmBkw8WDD6S9M9pd25ZY3xzOefpN4FTuJshrx0KDktRfyCDWM1y7obbimUAGL16d2
kMuiS+yan/1sB0HmlvPxiRLoLDGT/FFNkNhvi6foP7rCLhx/6A07bNxkqerDj9cEKeuaCd2p8mcT
I4/kabDXgmFEbJZYC6VQc83pdtOlnAFUqEqcdH3+wtAyvIFdBPH8RM5emIb55sVuhmQ3cn2QM2RV
DSuI9O6c26q/eQPnzMxARiuM7YK5reGmxWotQrvqvlgRzoUYPedmJYYFiJv8CNqsYQXeTjCD2MBP
a60EfqmXVbTtE7/yP0DUZrrQpeRaaENYBXYdr0nwOHgx6GJhQ0VtH67eqrQn4QIbqTJKZv459yap
1FTCB8PYnoNqnfKim//Qo3YcOPCiQeH3biDWamXwyVwISUHGQiqHmFbE0YpQiR/ez64vgG388II6
F2iL6SxF9TMX6/zei6U3510SEd08js0mX4NTS40xuQ+98/NqraVvpmjVOXjm9HdtmwLS/MvjPjrA
0g4CLBtBY+JsCo/Y0sg1DIVZCLNl+ePKuCtmzOuDZ3nNvgEdvyPa1yTwPJrgO5pbkgLBO3Fhu/jK
YsvTZ869vM4j7KZzPnjelc+gAl0ks0kQ7e3B30mRusuom6colKMPJ1TxS4UjDkmBilHq/YHAP+YR
BLWfxtvirUr37F2XxrgLR28RP4rhbSO2am81yeNZx6gHOjm3cApSZO1MhHO5eJ9243H4O/fvYtur
1Cg+AZLop9L+GuYzqckx67KKFZoCMdyEsjxjKkPI2zFOFwbS2OB1uc2lXMWWsEHaeFc+5Ea9n7wf
JxZH/sml7/w/Ue8yWx8LUPpYe1nsTlwFPPWG+MLubQHGhC/BOsPUeudDyRQo2pGtqhRwgU8q8jfI
K8/CvxavFuUkb4p8A79VEmJBOiDnpLOxCCTG5cRsSELghMq8jq8kJVO1gLI/LsBv+ceWTr2m0mZ7
fCdWKGjLPD2WQoHqFv2UUP1XzPqDLg6gq0WaPVToZjHgIe1/a2P1JlV7hzJLU7RPRQsC0m209rjP
I0r+uBv+vkdME/zG7OHy0B0go1SH2nqZTiMZLmhtq5wNVLx2QuthP7CndCIsN7+0X38mFBnnK0ZO
/Ku+gfvj/00BGr4SmD7t7IXXpOXrEUIZhTmyVSIyKjjARR2rxXNi+3iUiour9mX8raqTi2gIoml3
DRVd1guB8SIF60G8my9/GIbFuZf59iRcKMjr+WSyUJCs5h8Bm2v++uM/P7KfZK7a/+H+jbgJc9go
BqBSwodC4h9OB7oBeONlt7lPI3AfkzMxXJRWl69Fkrc9bxURBi3OoFEX5k2eZ7CNKSNO7ajHGtaG
iaKH8x4ziAF9fO3rNUWHaRVassiLy1dG1hEnYYSf6to2MIUPDzhimOvtKJievc3lsByM5dp1DrkD
3JaMVElxQUD33pKq8dn9/eb9naYdDTSb4Me5pE3MZLUHDw/qG2oNovtgfohaSNqz8Pa1bP9+PAJD
Z2A2mQbKTQGp0zBZuWniv/JmpDm/vqTjkLKA9S5sy+BDk/7weZ7MspRaeBZ9KuIjHaOagcmmJFRC
wYJcRr5bVYp43NKld5d9kGLXaKu861QGo7K+NydjkPY4vM984N+kJTndEn0orYgg8+wXotK2X+i8
WiY4Y+kCarLYTvcgymowjV9S3HTdIvLKij4oaCJKs06dnbUUu7rycJA9N2lxCsitrfP6/akk6Ggq
Owgbq3/U8Ezyyb7sQBTGx8i5f3qUuSI3X/tq0pgGDiXk8f93j/71v3Vv5b2ztuo+TAX4WmoYff2Y
VD7UEuB3mGZ9JJnojhmNiWnOMq/GOHN8D3dzNZRLxbCpi4ahBhLQ6o1hpYvLZWUT+ADlnY7dPJLx
s1npCqY18DGpmrIRYSWBF4B8eucUzlRhXPBj1Xq8jdlRieZnwRkX+ezrFwmcN0ikjrOHNUotWhOV
V4fk2QIhG/ybDXh9WQGsGyJXh5V2+NIgb73m+cnbZSy0rAwWjX8q1MzWLuNTI7I3Mu7jpwhHDGvx
nqK1MKddzZOekC1lsi/H+QmJdZI6V8n2ObkcQuzCMy/12A3P5oTJHHESPDjvh9IZb+lFyEkwTehQ
+hEaEP/KWq746KSxEv0HwLwDS0SEx8gWP95Ea9uH7Mg17LPVmcWrCxhFkEM0XaVQMDFNXaiDbS/H
7fuvE/viZ5ea/2r6q3s4MLVE3YOoTxnxJRhMLrNb1wrFoVORYn1YeD1lFRYH6rlUoWBxsDag/2Rp
VYeYRcRftv+BAze7+MDL2voVT4glNsVZOdznzpUiTTGapsqch2KF2GcLanTvdMqo4Pn9k7n0jDKx
pXXkVUIaeliTie5pcE5rpidkA2sIS+o093lrobcHAhAtMEI8IrhSO/s2nGfTSv073lEjhtzhUoIe
w53J/q8uwbi2Yw0A/xvyrKCrmK1zB2l451h+it369GuPmAvlUTeuJ/dcU4EGlP6C5rqxcuF3UjQp
zdpArgyB/HrgJr+xkz06WBBfZBMzZm0ovbwMcHwZxcJzeUnkumSRFg468e5KDLVk5RmgNitAEgbF
lzibkajGY+bRbE8cLLSjV6LYeo/Dn9DlMKELOhqCDVKWSh6Qup64x9+Zc8/u4RfNBYcJaswmUfim
WZmYvX1cSOHvo2TtWY64zo7A9dpUXEP6w3yK14yvchlK+eq/cQZXyb0j9sA9cra00KWjGSKmCaTp
qDj0d9cofI91w31rUqDPfZ4ppNvC5iaYpe0MFNI5yoDEvEekZvfOdOvVPI/MEpbs/IB1AtYFCJH0
urhBjtM8VoGaVnCjWl7JGHV3Ixa6tGroCjAF+N/Cc/oc/4PBxJAI3fNpTtEJlJF3r3Rv0ZPTVXBy
ADLWlGLT3igcTIPSRxtWFO50YaE9v6IjpMK+n3HqkgpqWtfFy6BeEYanuzVe/C68dxL0jamifLzg
m+8uvUFQeXjnLXkkrO0c0cXJHwy5MiCZNZpGW7g2PEwBKmSlJNqqyC1zI7RacAXrcmKvxvnOxkem
XdTS7xSs79AJVOBMeLNbHlKRb1lFDS9XWmjWaOJkCdXcc61iR05PjCPUnz/yu8JLxy9Jaf1qSEdA
TWx9iUJZpcEbHdBPMvGHq4AnRffF7zj8Pg23KSEf0YmaT7XB3sZlKSztAPHmi/QfTV1QyTWjfAI3
jup88OAjOKb9B8DEbuG7BCYZ+QH3HLTMEF1mfgrAiUEqk2JHY8NbDzx1M1XxK5GtrAIxHKSUYqKL
i+gBsDwZS0iudxHtqDFG0IbDv1lt2jdC/pseXVDsBoSaDAqVyrEZyqJMqH5d2718GdNfQ15n9oUl
meRgz25fi8qf3aExZoZMygNg6H3eJbEKUMuM3g4igD+ALCS3BinPXEosjRQbmntBmqx6ClquzGyP
imWW9e0rer7Sn/dYwYBnd33e5VV8AkfJzqcUk3dYfvTGs28kjNdyQtMKoc8y5xqRlEmh+dNVjdeh
DG+EQTxRAUo3Yzuo2fp6C+ncjQmABEIX8ttnbG5i8PEVyHpeVwBMbEDnOvPvYxS/IAGfXZ0m3BLE
WSuxC8VonB8M6ojQQCyIFFj02uvsUfMEdIqRZLzUe/qcEVw3PJ99mq+sdtgyDcn20JWlXFx0Lhn8
0f9+MwWSaDPmZTLKHEQhJbvMpWnlOGDm+iPkbLIfyFkvMz6vIZN7miCmkrG+iMenSkoCBCQB5kyF
OXp4zUqSvwIsSCxJbt2zn7wP/u+Qtklk08igUq0LdvNFBbvk7J6rC+jOTlxaoBSjBS+XcPM8/W0I
AC35cvRcOiqfBBHMaLvUsBeHap88RanD7s8/3iazroyWMUSFwDZxSAR3ZgcH728pp1RdHVmCXOT4
TV4q86jUMh7fa1dPK1k+8f7Xf754FTtmCW4Ga11u1RsLYUJnqCGZ85+TaRc8jpIv/SOGiBk/0MPP
bdcE1Of1/ahaypC78TM+V3niVY/p/SMNI9qK3rn2cu+uxkzA4Xagb1GAXovo5Yxg1aqnhy7lxU3x
QeWW5Cdvye1lTIB9XfmlM6FddH4PkxBqOGU4z8pMGI6VSKjZcf2ZGoabEg3Ltqq+tGebiPvZnLZR
nC8TujbXS6KhMMcukVOnTAGCOaBSoP1419HaIgMFn8ADb3XCPNYBAteUDxrFIxKzqGbEF3tqikvq
6vn2WhPOUUxMt2OAI5CnuNzg+YDHk3wySlwifsylhILLYTN+2Wm2Jqx2QtCTEw2r9UfZHoTikelr
B7NRmT/vkNpi1P2Z5vvPiv2uoYNOODTVou1ngsx9m2w3kGj5L0roK87agYPNw0vnOSQuwELkpW+m
qDmi9Fi0uLb2L+GYZCmNsViPWCDg1AjXLvZZOwKmaqcIbdjjJ4cPvhZGKYIE+F2QYkG8PbC96Fqt
QS6zPJXNiTOlcdqaxNL7mYUcr2hczK35GP3uS/4SE+I8+gbJPK9vzh6NAdqlvGwOeKGg5k5Lf9XP
N2G27Ykc1y3PqD9bhAI487r9AD20GyaaAzf2TfnvGSIRxbWa5jibZ7XSeqtFKsm4llJSmbk+QiTm
PkwAox35lYDSp3ldSlKzVY5AVaa3qo7cRUv9bUaPNSmz5ZqpoGQ31ZSi0KjpUlQzNHNm0m+VXvc2
tadWD+9LkJ/UacgDs89OAPZJ4h3ENcmxyKEufLxCfBTrdOQY4F0KlO2AjGC0+5Yqi3tWJzTSxO5/
Q4SySKG+RMTLX45VfDmPF8K3K1iTq6HVLk/OwZvvRAeop1/shyntDVvsuUxFcLAxEsUi2Hy0ctQc
E480CQxVGZsm57x/k8ndEySJt4Pz6CE3l2U/gHcWA3ydS3u9LUIOqmSDAEYRQoevO13Clt2KJc6I
jSlLvzaSnZVeFiRbZ4eSQEbDet0S6FMx1TTIVUphlhmWIKe5SJBrs8r6LX870qG/Huq5muOwSgmc
+lZH9VvkxB+HhjxZbRWA/4N30E7fxCPXo7XR21eOfKEo0SW1Kz4RBw6XFz6u1Vs/tYHPjjvUvplD
I+QrjIw15/czgwS5U/Frzx5FzZYP6KWudt0niPufi9smSWzGYhhco/b8H/77IvP9adnHZvWnQWpv
OJrswKW/g50E7cXLG2SgBj/i8JK+ehHNmvfsfli7kc9qRrm/hRcBQVu0tW4GWS2cdrvbkWB8i0iO
6sEfMSNVHwA3YtMb/ub+P+A8AH8HNoHIsO6GTCrD8sVnfSZbwdKua4uSEE7NZppvp91kqCdU8bOl
GiZZmERab/xHQBcUlRuJfYuwJtFBZer8oFPt8YIJBnKO4rrnXRQhgMBz0kHLqkm5jeFkztoPq6Uy
KF7wrx1DJgcU7RrTBf5ncySLYCqvL4gDeP17UrTnNvcg9s4r+sm4UQm8YoAlX+dDu9CoPNZs+QJH
Kp9mrDUm+1M4VnEaFxihLkZFnIleiK1D2ds+jbw9jOiOnwd5xLdaWurAXe8LVa4gFyU5n50OeCFV
tTNX5FsgrY+pNGje9A+3CE737YspWRhZrLiEMhcKjbg87Y8sHNGmynkDWVqCibNZz2t3eLall46M
hiofu8G3G1QyPZDTBGV/c0TEGzWx/Us4mihzTKUO8rzbFGT7o/j57iykSzrmKdERFl7MMoCQ6cJX
7tTIh803WgWK7iODR89WpuvNEemRlNoBp9DXv6GiYew+PsxJeW798IyfhS4T5w9vdLf9HsyhvEWD
jobaTNvlUZfa/yDmu4mBXXdULNyvYV6SmUBhkDkT8Gqx27OQLcP7I+vg2lKMMy5h4CzEQkqruPZu
FdJlc8MTg4AQPuAZ4uQxQCdL+i+BxrG0iAkzLIf7T9MPTrsHoIXeWCOJiTZ4IMDBJfoGXmZE7yg3
MBgGnH5ZWSoWvAErT8eoB4QlqKV/FtGQsqPXVzbExWbRKqQUfMRWF38xMCj/OUjxqqmwwddc5Q8r
r0EC3cKL4R5VXbn8iRqWlOn3GuAJIG+S+f/YNsvLq8EaXtSagD1idL12kOFb4w8zSvfOVLxaLgDD
Z+8+V9bIXO3SyLTQlzVkqrrlmb6eOF7Z+/mYXvXYHllDMGorPrsUwN61RVaFFJJozNYouKeuVUpz
XCjd8sBrIVs40LG53GwU9nSSEe9hT1RMOMh+PGuEOyEZIjr/qiqaESP9gxIS7d7KHcK3RkJdYCCY
OOWjlbMUZ7nzNls92Di9+pYDgpWwSrQA86pwH2q2qbtYjtmLv45g0koD1ooCJpKtfOvCK2fCLzb9
T1nfKj3udskea2EZFjlz0LSpNwJzvSVyJryt4LX6E0EFvSREJCoNbn7aYQXxJTQjtTuhI3hCeUCo
9hTeuBEvoT6xvzpxJr+oRmNb8Xmi9Wi84ysj52oyxoYjWmy5XLrnHkmlG6s/NRFBDSqXX3RSnVZv
3hs8LyQVVUWjZ6C3Q8gHd1SqAEvhb7oUMQRA/OHX2+7eAkY3s/PN0CIQCNAtiskCcg9AyGeEljdN
z9/tyEYmFeoHjjZkjnZEp9BYVOlFfK/UYF4QMYg4hBfyfy5TnWfAmHj4+SSsTvfRFu0FXhrXJAog
eCpZ7s4ef0HkU8AzV7lBMAsoM32mCK2PjdgasV3HBr4PHjLlzirzHz78PIMZNRa9OLJouNUloLLr
KTiKUVnSrkgKKidVER+tRz4gkQZvVVRdnHMBZgzp7sYvaaphNgU+QuqP8OxPYH9ImXnT10Vk9Fdb
s1qbp2EHmJqnbEYSaKI5P9xd7FnW/GKpaaiIqJTMijmr+rJQSSJ6e1UX7Bm75lxHuJyRV4Ec5SoY
IHZXLyVGv79JIRS2RFiy2XiSfO9MDcH1yjV8VV85IQzq1eB+1QsHhIqgR70kUOh0ZRysdZCVgBZe
JAHz4Jl1hgJqv7pY3OkU4VgILRfuV0cVeh1GcPnYQXT4GuQOKkPcAsvaqRdexM/FLNs6UmwXQjfg
31/GR1fBcwFg4jb/Q9CPj1eEIdqihfl+5LnEFKkjcUghdtPu1fsrsLzZRod1GkCRSXEkiMeJP0lD
fl7FKFMXjinfSh+Ahvwr+4I0LamUYP/GsMihhpx13uEHcUbNuqvfLqb4MpRgQs9RU2gTYgGxsSHU
/xXo6hCGlWmzTiP2wqqPtTcdq0iGAfQKCShLHHXaEVQ2mXQgEsj7jHZf1bwSK0Zb/1XQQRix1v17
C0J2PzMpB1gMyl70ZKtRMVkjz/FrFUX5hpOJGs7+G9rnwDXIFEVTB0cKoukJtixkr5YYR1C+Qg2B
ECvzsxi2xnRefh/JjxcgLHYejA7nXjTAgz8JAkN9IegNgeNQXUlWLA2QpBbYg+jn25fO7JY7klLl
ZUYSU1U/TqBDJmv24GJnNDkut8o7v0bsHJ0Ak12+CRb09szqtgQZaKYUlppV0JgZApM0Q6Os3PDX
qifXH03CXDNiQAtZMVZ2E2BeUhzdLquK1RMQ0klqqT4lJVC+mqR/YCvuT0ht6R0R488Jn1LKm2No
v8AIzHGK60jbIlFVppzU9PO0w3AtbNJ4AoeXdMe124zfaAy8GOwM9t2seq4wW0Ma4kYvutqDuqxV
QBxwbF9qRvscG2oJ8iEvO2FFYbPvNMFZg5OCD9HqCmI3HTE48/45KdfpI6uFSVc8nUWgtF5ie9zx
feQfYXeoSbHV/mMyhW/PH435aZcqg3j2TBPD/dkatgj0WsZNR2OGE3LQ0vhAwIreN4kXX/+0Yovi
IvZSrTlxFUXvze0KlK5ODXJ4WjisvRJC3MYo5nClYEYcUCPh0hA/l4kekrUtoMzCGbrzocCwnPWw
UvP7vDvngoP6kAEmAK3kfY9GMMV137bc28fWqMPUs3vgLZm5q7OttDalbSFX6CuRLLyPadCwQCQU
nvXcbg5cN81f4OATh+n0UrxMFph4pIL5I05wEBAUNCGY2XNJ3jRere6Vbvge4WsnBHx89wnnz+dK
ytubesc2Ccs25+DzdtAp9QF39YAfMdF87cGHdwKkbA4SF7j2azRjcxAt9huOjT+s5NkHSTP1cGkE
yWOF4ZOt5V81ijVnCmIYJKa8v8K2HFGllT7FB0Aw4rVj0rIIhCEX70BHVZ26o/Oi4Rgeo0Otter6
Vx7hFCZzWcsHt37sC6P5iWxV/AZO8eAwDiSodeBR4PoIyemOjc6k7hRNUwhcIKx9aYms1P9n76CH
5fC4ODgqwJdC+Ay3k2DctO2UJ9s9ajLMc2GaJTYPnS4kv10LC4KIvwnrSI2jByLNavM/Ts8rPg0U
PXkHGP5G0kGhTnoNqlAIwQ9gm3Xb/l6iyT7rqTyARy6WCssfWzcKTuwFFAp45890hX3mwPmy/d+5
dqJ8NXXMlzUtudo36ey9Q+yExjssIAuNWc7E9+UiffLA+H/HO9VSbhZUCeYW4/plLeZVVFMKN1tL
3XgX5zDAZV8DHyhMmpFe4fN5kb7eCnqB6EUkRIfQf8o3lRd+RtT1Ts4UVYCEEabTXwzuAS2ZPkGW
TQepLi+SxR4OPjh5lvtK9XsL7+++SgmUqlVLWi19mks6wepIMcyNIbE6gxWGE1+K0SUnvzi24LKR
vH9TfFMECrYRFHzwthw4O2l94aNZwDgHUV3HHdEcFs7tk42KuDAjoA7OUX+GL2PMjwcAFQKT9zG4
dH0+Iz9lO8wituUZr3lAm5ycvuYyC1fu/U8odO2+XC8hg4tsq5ckdCR1D39ZYqGb6P7T0q16LOXh
wxYv4xtDtWCa8CDlvsrOPt8vdZ1Gm9WwylvTMt1tnELBeG+X9ZQDFI6rT8dqAq8Kqztj6D9TtCwb
EZtFRCaUjqp60vTV66D9NoquN4++KljRvRNH2v1R+VJzbs/qxIRDGmfCW44U4F1Ap3Yiy8pqaWuX
KJ6vetdUXVDZ2PtHN4Uksz3m+8RKx0/SJaEOPoBObqltvlpnTc16VsrV0uc2H2k6drbhOHv6AJN3
7ArA40/dyk1es/4hm3wQoIaDAYTXhunXkq4x8/ZdkuizPZZ42FZopmpBTSwigsDpKhKX9xZwepWn
KqUZSOF+Q2zZNfoWNQo2sJ+/K9whcZC2U0/KZt3HPjUqtpBuozKt/GlrFiOBHvGIeJooGzm+j82F
SN4ZP07Q63m7P/9JD+1Sc9ieIAc4j9Xyzam+FN5MBQOQ/nPFZf8MNdS6l/JqwJV7/GfauaPRGeuM
IK771yYbVJUEriCeTTzege4Cb1K+WJ7ZBgNuoeOjxOTEMd9Xoc4er1qxLOJfTi3ZrkTpKVljvt3H
xuiJpJr7AhJfZlZKvayY6+n4+fH+SXiP5KXbvFtHyoIZCzLp6/LftFXQhDWOXGAfiXMnX273HiOa
AttmtmavJ7z/dUKdRPQTt29LzdPxTzpDt4Jfi4jG5W2RqP7ze+sFYwlivKRgGue9vVia52mUCPa2
qiksWVwgNzSzr4NHAZ9aGfu5H2QBSfRehysztiPyPHDXYnrlusrQ6OfyocN9dhAfWtwglmslMHE8
CU20+THPZ359r3n3MSMZlBJ6X5WEIyicsBO3kMelRLoYDdJs9OBzYT1/jXpJjeHCABM+C1siFV2z
vSvD4HvF8zx/rb3I3wcBJk/1uGWPZoTUTep9eV54neF8hDuYW7vjc3lVT0QWV51hKZKSwJ5vTYox
FUO69wmsm5fYJ5peryG6ll8elfmOVDOYTU22Vlpd8k0l2FUHhx8Hg2WqDeRLxbwH7V7H0OfWuG+8
SN0Ndtzsb7f+PJJlBYlJNYtbx1jbLULe+IudUYb/+GIS6OsJR5neV0zm+nwX4pj2QtbeeMgTGXnK
ep03PUn1FtbLNRX9n8vfdqeXJPy8rcFMZFovuE+qxJalTrPoa/mJz6sj/R7mR82aiMmMqJm56W+h
xp5oEgD4NUAoAL8i+3sjMX1fpuMpl+didnpRJPJknsAeGoZSLL3fW99zzgGm762ASYIvJcoNK8Yd
1MShuZ9C+m1Xa71iJlWloTGFvq+PHmqB5+fbTZsTEDVXoJB3G5ykQYRBHgI3x8jY9GBBaXKfFZLD
Ess2nDtAXPhkFJLo46PwMcd8RQsySpI+Qsg9xOShGl6PF1ZHveE8pQ1Z+sBhONsTMzUa2ht90CHr
rEdxTgGSDD42tcTd4zAaLBRWkY/N1+qhG4JS3svhQlNLynf3XJWD5g82a3RQ9xz/Ljl5dH9/GbjR
FwP4sywW4QVHHeXb99T9T7AN+wx7X3hm0HodW7KpR2BmIFbFCPbb0bPseCGu0XotY505+UZyuo+V
WM744A6KM/BN4Y9NWElM5ZHyiO/PcS84XYgfyqOHhePA0yG/j2vVBy9CASchNCDbxizkzMvVLwHd
pTVytRAioNlxPZQRLqASB5ieN963GyjP8R0/7sqjPgGHh9zOUuC/mqXmeThIyRA6NvhAeHWiRXwL
Wipny3q/I0itQc+j02/cpDm62dPafZkjMWl6/bRXQX1fcNBkNRklQT5mXc8a8eYwaG8h/26uzsas
ar2IfLpM+0aMiwj4ulHuDoqx27m1+rFLT+Pn9x/uRB+WmHyvP7h/AxbCO9e+9iijZejEm9Q0N4zQ
mghMv8WFSTfiiOJKYOzkwmT1QzikqjjQqV/guQdUtQlk63BY0XYgPEAytP4ZFPybHI6WtfgeItFh
igfmjtW1PCfpJCNueSCmzHkt+t96tb/R7yE++kEcnaHew3WhWFYj4gDN6Kl4c4SFXE828OHICvl4
aahq61pcvg99y2PgawHvEgDLNFBarMIfs8EKT5gH5prMMAXUeognZX2OrPl9b7+HTGcezx0ER416
4e3HdOFDYHkgDSfhxb63wyCbQws2jx2V/Q+akm6Hkxoej3SFxOKvKUrZyQ5x37ZoCSHt+f2LtyRE
KUvvrZjiplsucLHcvs7qITKxCAy1+m/B0/+vPb5Vw5cazL89dnQUamOjRioBKhsGBSL19dNzPlhy
dlykaLp5NtJBr4rB4ALTZ+pYztOLp4Nti5ssTexn4K2Bbxk39gLiwSYICQcogZdgErwuA8LdfIVv
UjAl/Md3vo+dikdijYrc5AwL6ja66/53ZHW4m1mMMLTreXtvCMLf3F64NB0iiivfPPjZH74nTPMf
C8vSb5oMrTlXMHB99xfRUceefOo5/YEH8LwwXgZzpGvR4k3x2+0O9ylJ6fApm/ZQqG4sleyR9DNY
wzp0iT37UszoLCKhrAg9zcZmF/FFvCTIJEVlN7WjR+9WEwOnARNulfO80imco4hb/wZS8w1LJy3P
HbvJHkCz8b8e+RfqizRwFMRmXssz0S9sQ1t6gkYUnmAZHmy9J1Bz+5M07j0RAy7np/pPWIdxI1dD
qpZlRnUo4l9BugkY0YvjnIFyP4oY6+TJPw4oA6YEqZ7qAngJbrpIt+IseqTWVl42hWB/Ht50lglZ
bvLxH8USTKhu66+0DoKMvLlaL0YGVJ0XGQRK+cK2/VZqJk3VPQvU9+rvxk1tNOdsmoYc1pxrAS45
ngIqL8dD2hGcexI20K7Vb8iEpBsUzO8rPuL7wkLnA+MXdzCoeCULs64XAgid1hlACsuvRrgctYdL
TfnOz/LhmPkaabkvULtkfszIwHkCWwkXDWbEuZAa/j0B8S0gVsoDL206mjCG3uVROjsZq6BVwSb7
CZr+TSSMhSXnMvtTfycDhkCli4nTp9CZRSjOFMf3qId1bUEEXb86yCB0mtlKUtd76+B9YrF14HPZ
ncktYKHWq8vmmTSCYRgEy1U8idiIknjIn9A8QUqUlRa5EKdB13FeWbYq6a3PK92H/NaturBYE5/3
eh8WLH2E7IaS5KQQ5HXTOjnVc8q64JrJZYuG9sKzQOhiZrjXCWyouR9cQvgLubeznHtlF/skuaFO
BfE5rhMxwhJWMKWEpgzgygCegeuqXYIebljyeFegbnrH6rjOwMpDh+xa4kEEagYa8Be7lR/PeiAw
LR4a4IB1dbGcRVTelkHc+AH9nZ8jkMNS22/BuAbO9885orF8ZfmVj89KXo8YbxJ5RrfvaS5GsFGI
HoeiSq1NVtqiq9J4Avb1G7xUOp6SZJQIoqXyqrhFJ5piesbVsttPK5cz6Hap+1Jj9JdUN5v5pVeN
SKcIBjy0PLxrwzmL14btyO5j0HMAV04R403+TV7xe19gO1x7SyuWZDw2v9dcqpmXeDeDqMWc6HLb
28kN5sLcgT3UyepN970rSAuDpYl4qlStc3NQgPto6y2CkRY1fCAyXZNGAxse1pZAHPZkSRkISpbl
aP6Gn83DOx10MrDimyvEJ2+36Rgf04oEnTvIhRWZLdQ/g6/gxfUtaZ9QnqMpWbMi6n6cwBy6RXtw
WkJo31I2B7JzMGEB+J1kYnQKbaukiby1qGj7ydMI70s8XaAlyYjdL7M/JCZU+FBcMZo16z435DB9
XyXMb9ZJPIAiaATjlT3sRrBMMKQkWrpYgrgQ7MX2xhKO0vTW3cLOKHLfEjJ/bCSyUp8qYASzWo7N
TUdOQ/1Q7GgLrpKzhvel3Lw0pyWJytmnfogziwaJ2uhwUgBqqwS5/+ZxBqkUznHukXm85ltdKi6F
qjx9xCGm/qJ8HUGwUT3e+WC2LTFleZ4x147B0plx8RDm/Rli9p34JjkO6qkgmcOawZds4VMJfocM
f+huGD/oIG5LgnX2olCvtcjZED9ttEck/gyyPCGJjHfL9XjPTXPHR0GU7ExC/ciO+58UchxH6IkP
t2PEI5jj7Rk7p/Ck7bDc8cNJZm73qhbTvnbFbGMuZ502dMsNpb6W6nkdncPvSdevotuvdpDU1Ics
wpRAKPU4N3OJadkU0n9tRX/LB44Jwezq50+oSXlDEijkbsjmD+9X6NudqnujfI5/ayk6oUTejbIK
eJSgmjawENjmFVly7U9Vh8rmOXGni2FJPlwG2BQLv/CKqCFGzrgW5Sb3IJ1G3iGAnDZbXwvNt8oM
TeLpNHK/MCopZJofktzNO1kpqFipZJOvZKx6Rj1Fk6WMTbH0ywDx38ment4fXolVj4qmBRewbVDZ
5b+H6Ipp0G8h/mYbhsCUzE+RL/LJG83Ad6+0wJQ5ZimqPEzya+uBrWkF56VwMxTbAX2g+Uxv0uza
MBOpwwh3x60ers8efpzC5cZjnYdQa3dfKne05lxucF0cPYkP8RKKIFbVb2aufTwSuyV1VAGKBOW5
S5RKTH3iOOUbib7bp44wsNctNGgpaXgBUmqr8bOe7H+0RsvIVmujDqZXMyuY7ggFkK64P5AqHln7
k9RnzDDLniUrf2MnwB7BxjHNGir/hPfbOFzeyGPD3E4Alfh9WGxrrI+RRYdmreDx4dXKVG1D80Bo
H3KuhP+ZTKoMqP7hThS+HsDGNNL3+t6fNX41DOfor96JoePH0YTSd28ehh5TqwjtGs9/kb1nlXxO
zDxaHY7g1MwOd8xCUBLqzaMrbsfgx1t07DjM14AcfquVSOYZfBzcsTfWRy9Pm1LVQDZfaNFNUeC0
CyCVMigRVZf/NH+pBUR/wL5VRK9tS7Nax900kyeSicry8z7G4NAkrGp3/zyZpqTyg7bd/Ze+oaTG
0305EizKz2gEjQILO5nIMdoMPM3dOrXDs0ehFj1mKp8oeTlzX9iLYlMmb2u26gF4Rv0glASBK6uZ
f7cOs06wDXueMgZrbMq/glb2JANpnMt9HKKAKvCA1F2RmPRyzc2VgL1noWr64dBKUjvnB7xxfjcp
eXrBM42GtQfRSgYv3PhWLzNbVKygotk9NeZrQdliZwr0mV2wqcX7rIg1bT7lmmKJD0gN6eEOLk4Y
Qo3khCIVR4kYNTYsk+6P14eq4u1lVgp4bjJxfOhc1rmWV6KOVKMPt4RbUHC8a2t6J5XHZp36NQP9
lLqg4CUrqrbQDAnLkta5B5ZxpTSqIe3FyHK48jb1kE0aDEnkywbiC9VAwxV7bntvqAm3gQCdK9tK
zOggN26iCNIxwU/634XUd33+dWxG0Y0ihMKIJ8/NV6//prj9amEBDkSbmpI88eC7kweHYero38Yx
8RKmVQBfzS2hu5biLw/OU6SZ0cA4+17vpmV1wmuUf9kbVLbKdZBTGiAwPzg451n0Tk7m8E3KjPaV
pZBHTnDHOJiGQSSZ4hmy6MrMQXvalcWumVfehaU+ynrj8cjlumFcYSzCmcaRBZa8BMWDERpNV3yd
DU8PHO08ui+k7azzIyCG6uckrLhtejd7FilfVBlxCy5A9mDTFOLskGbl+gZxYuLRdNHf5qBTPVh/
hTaHIFh4A1uG4g7Iy1kjj1oJI9F52gYqwExRvczmgEQMKmDkpFoLQdBskg0LnmxDA1mki5xuS6dI
2gzE58jHkDPVM144T8fqlgtHZQ+ShveqeC+QvPAkIDXs53DmEj2PyYIvVWB4MKZ+zoY3RJvyGfaS
gDyxwRvPZLZpYvAoHZDF080od6aedcukLWVznqvfL3GTOOrX0hWg8UMQoo7p8qMrxr7OK5ygqTMz
o9y7fqlIzWG2AbfbNo1sK9a3uTe5uVi+5ixhtAFVSZeZXH0prWF7ynhDRt0w/8LFmH+Llx1TN/WI
3ZKoXC9Df7Uc5MfnuP7EeVshFcGuRzArLxcqZg+eUPUoB67BCLECsF0A5oGTUNQn+sMFdmTc+ujd
YBFdmRbeJ+QZCtMO5voGkcjZ9YXvjjsCpHnD2Cdki4YZfN3Z90kHC2LYooySi16HUFDwjXab9G+r
TzdJZys8eCVjht4sUDzr4zjY8YeRCSRZjg/tfgfvmPk96KFye7eeHGw9wPyiJHxs550Oigljt5PD
H+vvKSR/13qZ+0N/3bs70rnLXTfeBgyckYWBXQrfVw/T/DmGTcY07wA6hi0gNpHSQ3pmIOs44oHq
Rtujxxis99j1oHq4iQvPEfJI7HHQPkubWQz/cim2Gj4/XMg60ooqH9QJejO+UweoChkc1uFEH37K
OvCllCCdbFcQaevgdo/xOflEIVWjhceyVFfc1/6O5Pbt54ZS7R536rGi3pJyUJ0NbTktXVIHsnF9
HCeCdpp4R4O78FfiIQlDi3hwodRWTU7/hWWSyd+r1ahWdGR/fJvcjMKQR/HXAdRTApA65abgvk6y
C8KAWcg5/ZaNO8IOpw7peli3kCDNMmfu1l1eKHcSSIJwuUM61P8DzgDLkWtiMLjvZncNJaZB2zwo
0++mG5RsisXTFhCqJ2gj1Whv4tjcwO5aMKScY3DXAQaY2G3mVaAH4Kb3DLUdcPRtHSCJUoFchLIH
FAsTsn5fcWgJY+FtqfgfXeNfPvVOrAE4Xsb7qzBgRodsbzoEGBu4/3BYgCWEJFc3cUB4qrB0Y8B1
61yDiBfOfKxrmF9RTaBw66ubL5I5kKjMZxN+tNcX0QB4RjqkykCicIrdRxFhMv2pnuwWynpxkRdj
Ki+avPP1x33FhJXjyI4sXR5+cE8JmzlHE5q1Hwf2paolqKNDmfb4zy1ZhOugNpL2qmixNwKLhgLr
Lb0Ev58xXVDbl0vx7REMj6+UvsKFff5GRxRC844d1L0kYkO2effRHqOObyLDYvi95BYQRdUkViMK
M05cvQS7Mp+0I7hmMyqUdHnfpWieCXIhmZZKcl6jZ24+EfAg6RNuRjGaKyc0kjj0NjCZjKxRKe8l
ue7SPSt/lkPTVe8WNkYxJHBU2xCImaoFodI1kHsJD1+vecOKGtD6oYfOL68FiptA6Psr6ixEsk1k
c+Y2xbC7n5LYw+7N1i1xUSLaXYeaTeuqWckkFpzw1J6UN96K3kxddmA5IMWBC0RB3orXFeUbNEtn
IC/F8eMn3pId99sYRSPmxoXFO0XZ6m1MbIk/lq6gdCSXigyoTFmDUt1zBhMEvMbKVhEwgPFDlTbO
ZFsvUFprbl9wVZbmn/Xjyjgq8q14FKhpB53iMUVPkNQYU1cdxdy3X3Z+kn8Po0tXR9rz94ZZGhum
7flhF4XKf76w086U8V7Cina4uBmrLtZ1oE5lBguu/q2waW8WgaIxi1txWJNB1fINyS73G+xyWSZx
l5WoJnur/xpunULG8vGKfmdOqiRomnknLg/FjoxYU+X/bo9Wk4mykLwvJQJX08n9bpmwt4S4Ha60
fRNpJnlQ8FPft6DzncuSbacqCH09YsCZiWY5ih8zI2NbIhkL4IOyGb3kIKeRsnNx0KEo1nX9pow0
4WsEgBBQganNsZ4UAh/Qaaz7VXIOZFZW5S61x4deSe2TkBv2qLnNhvpMfsvjmu8hjhDCmPK7A3h7
/4bBW7KhrVQ0dLWCS45p4QRMCykTKNKVvlr/THvRUUI1Bt7G0JS7axky2YKl1h0BYsuhIYZ0FILC
tvUnX1jVtB9T0rtacrM1skWQ2u8lk5qgrMogUR7QjUppXtkKwxs4k5ODw6yH0+9nV/K84ayYuM8x
ULNUFdlpE++NzW+GHIu8nQ24zHnXUAxhnHtSBkhmOvStS8Wr/F2oBCDOnM1WinPHEYLcezVpfzI3
r2we3R43+a/5Aw4OoUGNTA+IVBCKZ7it/rBg3tDj+LvhqagGmvxTOQid6obQ6+WM5OurHiOnVUmW
Z8PK6MDd780YED/GS2klA8YJQ6CaSDLX1Pr0Vj6h3VSHXT7+hwXCwRfHcFoi9haO6271f7P85A3U
kYMsJKrS6NqP/Fe7d2L7cPutliCZJWxIWp4UAA6qJ+vasSbJkwIE+cvtRRyHgxOZLLnL6pRqJru8
LJ7BtIJzyOFs2l8HhTImX4GFHcKie8V5mM/vCQS+XexXj1+jDOxTEhHwPB5s0/leGkCbrxBdFgjD
AmJ/9kL2u/9PShXp7MJegjdw0HmvyYdrKZ/YeLFdi3kcfbL+WhGGpZ5H5NMZdvcUdCBijgXqTCXU
z5vSqCW4Z5WZCJNeIieyZwOhOqxWip0BThOYXqcyrcnPRiqU6MaOsgPc0bODJPSMlYGPdJG6Gt6+
YLZIBk92XbN1fUBmJ9Fk0A6OE5gVj44hoigoFp6kTXAnl6lbyUIpoMh79fHoer3Z1PvavmnbZCTI
zvdS/onMVMZwr5VMa7Vk/Q/JHGr/ilepYyGbwZvMIiHPFoLguEohByCcxlBOKLeQVEeew5FOGijP
8J2n2zd1y/OWTnzuEQ/2TkWvKMU2XPQ8bZo06cixrI8ZJrbHlN/1jGZhyiBWOe6Qp1+jLoeayAK+
qGsBq+nybRSYIC9zMx+0RxbB36oQ7414I6Cr04Wl9+Ytkbaw+2F4ASmvOt6qkfLKI+1We1sSoDhd
AOSXxjoGi4B8uX2mGsYuN6iR0p9drq18xPw83crRjr7jPSPfGIGtONYYcKnaXb8p/qfZH/eAjHa9
NL0YEC/sRbADHLfq3QJkPHYlXMvP+7cxDp7YpQxFuG/SLv04eGtZoEj2ycAu+s3warhwASMCaWkR
00qBcklPzT+Jld0MaZ5v7euhsns1f/px9HH1RQdn0xgf/Ks3AW0Sid7An5b7ozr60xsczMb0ylc+
VZwv0T/88MzWWhYCWX7/RBZ2cYY51fk41Khy3tMTQeMEkF4AA2WnvvqqEIXZQwj+aZEm6qnNQ73A
8Bdc4YPDugoJ15Bhiil3e9vit+gG80t0AJRtZuqZ7mExeucSXN0q277kC8SUl3XSIKexyBJMZPyG
MfghleMKJqOThK3MpXsjxTFTFQYYzKbTFTFqhadBAMg9+5NHSaRL3TQ1M8fErYckynQuS1UmF+6R
uTqliAR7Bt95aQC9GCo5asPzIym38bhWaysmoxsAjTHfhP4PANNHyoS6qedk0VUHaxRz5z6eGz+j
4zdnUvvyjashLDqs3gZRjbtWLOMW3Itdq3ZWxY562oOjdWzcDgvdNK9oeZrsCTr+Dg98XwQKmzv5
eel3fyNMZbuIvwfH7j6MQfWaabk8PGuumQU8cv9u62gweFO5wAZ8m/ffJ8rKiRqsUHYg3GWkbX3G
jFA3/uaiXEFTnOCv2t7Zj98IaFblCl0izqHULMsFAeuuN+KVolj96kfe9rZTiLIHoR5QMddzHSgI
r6ag8M3AVRlaGHJnSgGFCiHeVkf9+EJGA7fPFdx+yMQhbNvwKE+XFojCERyZEiee5mlQbhvKQYv5
QSD1nnxX8VS1C++AiuUVNtm0aLu6oB6516ynOSExTHPiiqJdzeXjDj5XbuEdY7/DCJ9qUCA4r3Yt
SfNt/VgN62zffJ2d4IHroDbwX/djnh8do9jOJ3BHcuqGSruE3TAETc28Ky4Rc8aSFyt9UrdNvuHX
YMk6a5gMzUSWSJQuKyCrBjpfWAuaSuZGv1DHWMyiyM0QckkRqIUF7vuZi6Pghgmfaj1zGWtDEJJ+
XWDDIGfwKYtcB/wC0klpV7UAd4+vyxnuMJze+tmSZc4ehU2fQlxQwhtRBYuNxMmgBtPQ7qil4Owt
uSzRGSSDsmoPAbYN9urnCC5FA6ubq0cMj5EwDIpQCfgxemPwmySidJSN9/nl0CqpPtA/iFkJvn28
m3WkXEy2IMVPDM0J5vN6QnPV0zjphNDjlXwkC6IUR1U7ISSdgernPnce8A3Dwlhfz+WX4zydOESU
8FHekzy3snRn/Krsfr1c1opY8t3iswejGi0QTlOlpeotUFITf+6VccdmFxk62wij8lwFwQ5eeTTf
06FXEelz5I8or78q4VMPsQkBANzrSqdwbPNPyHQ/E06zXqer0YvVMPUlckKtkxuuVZ7kHmpGPQpv
J1vEMTJlhRQDsAeoRv40hB4qtKmEfeKZ9moT471RXmdqNMg++INDpNnPMCiAtMvmniriULtdHbe4
MxME2sUP46LHWxmr/fcTYpVseixtp8xjI4PoHQFDYLLOoEnI3bco/cQc7v2TB/3KaiBZRliR/P3N
XuytIyoPxuI1qLUVH4wNEU687hzstUlfZMBAIGvcQYEXE6IowqCyKnlZU8/P6pcTBEf0CmozGwMx
l1mRPNcU01lumtov94cjZjc+qrpncJ7Pp5ipo5T2dUEyakwCdsEuVHXdrRll6O01aTPcp0lQYIUS
CdqiCdKB1nv8cdSFNxgf6W9s/MeUMVjr+spt3TAG44V/amWpd/6K5tT8jgfnrgcsX3jXSYIqM0vQ
R5AJYuVqhUqMjFhnyeQ4ZOF8V/F9dP6X24duCJwZah6tro3YPc/Das1ze3MiKQ8dnmHhUxoVaav7
x7zzdRoFh4DdFSEA7LxaLih057TCMqOCDn9w8tLn/8jF5n9PPuLLadkUCC8vr7d4/9DMK0O6+Xoi
agfKcPDQeqkKTPGnB7n4v4xk4rT5ri0huedKpFJrVYaIq6hhCNkHyBDuAzIvH0q2VCK/mP9KjPNH
eY7ddwSMiEWMqGf1VOHy2LfhqpgflE3Ogq/hru5XZvl29/pHlgkv6yAxoLJC/o+dZIBp9Hu53E/c
tMOTBtjNwAGhdriKdmF1HHgCqVApCypRzQidPwHiP+NL2l8exnWe8OBgFJljHj6uMOB2dPT9sPvq
ijAtXyaNWYtdn0gngIkplSddEowqT+9E7GZAlPN+LOIiyHWhg+Q848EfnwqESQ3Uq1dSrK5VKTnL
M3Szbs6AHz0b1lsnRfx7jnQaBkuvpp6ES2IGX4P/tdx3lEWi+eXYJsJ/8pR+uMgpWtwPeVWx2Weg
JK8TmOKgw5rVW6X8Sp7QPuMIfTW/mInAq/ZNfb97dN0biGFer5jtoJwzdcAiSYJyiBwpDObUXjeq
zCr/ks9iBndaZurTV+qdRGAQVPXq8s0VCUZN9WqiGcTvMHp8cLJ+dElejeHe+94F7Ddut5x1qlUC
x3Ox1MQItN3VLKfR8B2XkwHVRIEzzw6ryEOwK3NZsFxO8By2Ot8uPWCBlBAQZMxufbUDut5lJvlA
NFKhXULSlo4cjME00SPvbrTDyxLaqo5rkndY7FLJoySLrdQey7ClgETOsM02Cl4vP8uR4UMhyaIW
Fo4Np8xupWaO/80CDdwIzjTeQ7X5Qz5T9/QUnFTZ/j1cw93iDoN4ArFDuCZeHCCE1NYA7yHEdaYn
Z3HC60m0GU6LkOg97QLMuHNGfd0Y5aZ9M+7MU5R1zMI/andXFZtVnFpD5RxvB3htojEV0XTnPZ2j
cM/rrt8yfhbIlzrMzcDZopjlWsymQy5ZQgipgWKhy1g+6nNk0JgCKxW9Q24fDpC1MOWFgLbUhITB
F2BqfmRsk+x73vfpHfzEZoj3Hln4NPa8ixVMl2O1e0jeNOXX3u5gL1IiukMJ9YKUU76nMKhS3BN2
7URAOpYHpwHSA6ssLCMS1aOHJS8pdFJAqX/Yfm772T0T74BdDGwHTMsT2kQJUt1EuYvFBj5dRwGE
OuNtEfpP0SI3BLfrgQhOdxRDh0OpPZiYHfR1fSgwLWVaeQ5/+Q4gXOhtIgpHl+qHl0LkAjfCr0vo
wRRIPoJlUTOhAUhGfdTe8ssObrnUuksHmMaRyNJR8baIeoaPtQrzsjgrOge3KS2EKPdbQT16K7sg
HwIuUlt0mBzNHkqPMOxOKWhhLMkK3iitEPaDVrXhJm+lJ8/rbMyJZ07v4B/uo0fuf6EoRDmiTRln
hEnmHUnt3itgZohhTsHFPJWuxPnD2FJemj8o9fS0/gRmPwKejrJ0TnmR6HdZDCpUIzG/Al1HtC16
oSVyWnDxQBOlGPMDU2IbV2q1eAYBhLyPjYirpPrKWyr8ADnWj7Re+afRPRiuzmtOm0NMP/a9CUDF
U05V0gLShvso7WVd6WQDcOUOmZqSK0Q7Z7dwbnNUF4YQtYVwoQeCvSgwGKhpC5VDr+U4pTgpLOQX
nnp2OJ4XP6WBYogcHxhkkKMzDIP5J0sWGxC31uahVJtn+bLsxtJQyeKcEPC3aLBAztD053QgFqcx
ArmvKHT475zoz9dgHcrcPjlEJpjWyAFJMmKYtXGPjZTEusaUNA3FckXjA7iCRPu+rIz82qAITlAk
5ZmbuoQEI4C4CpWN6H9AdQnBf+iKnFQ2bYMyYf96JLgAZ0m3KPSKavlAsoJfICfOj3jrgP2T0yDQ
hkHu5IEoRNEUJULAPGE8/4ZPpKSZNSvdHHj2MBsreR/+gbWt5Hz0DDPQ7VsrQmoaFrStP5PpNJMb
0n6gE408ng5MhogLz6RuGUg667e5RHOdo76+Qg1wg4JE0qOWUP8twtf55y3UnGNZ/WUs1O/Zb98V
GQPieh74hV/tbsteymbE7TWtyF1JqbjKVvCkro5+/WqeW4hhXuUKLrlZppMH+TtoxgdrdyBqUhQu
S6fBJtV93KtTNMDselscxoh0y0Iwa+exdAin3IneYVCj1YMg/bOJJVQxPxxLEvByNrKfO9scvQmU
1B+8FwC25vDy2zKarRb0VUs9Z7OhyRKm0Q14QWonjPtfb6Jolqd1c5hF4g7U5aKH5gj8eihr+Jm1
IBqBJJwT9seGi9CyuXHDIdNRwwZjMCoFoaDVj/RYW16OGSVFYLxnzlHElgFnpZKvXRiGwfan8eno
jaX1ZIpzw4PbrACugew0XyHZkPvyf+B2W5iJUbL6M63Vj36EjPJheF4VwoZscLDbDTCnSWAmM8gg
MsBJ7jeC+rU81HXhq4feQNb2qgO9F2hFXeQ2Lek4IJvTWjSUhYx93vBHWVNKDOcOAlLeE5GrsJx7
8E50SJQ13ipbm8kDGPwaYegmx8MjQKNhRDvjuPpil8+cl80F3xLVorMKdCmA9owTQfp2X9SmIjtH
iICXxET/CcbWa6w4/24b7hkCelYXtmpaacCY/bxjP23Sn62v36vF5fsfNOs8A+2J2JY+6rzq7Wva
ClZ1pMNQRROuP0LcA6YHWfOGKzlMX0rTqPF90aZUHZwbUhFuHfl5Zv9/tl84DAMXPKl4k0IqJUFf
JBnUwldtJOgFXcA/sNVp4bpspBs2rVGkrsupRstfiszXBH2Atdwq73erQHHHD9bwXwmlgdabrrlv
n9ErfxebpFF2Iq1PuNFI6qHxpLm3wmjeWiym7lNTkUGq2pwfaZM/XyaT/fOx3sgxGrusiYHdbFS9
TIAyAdhO9/ZpJgUhle5ffprJY8MYiKtNSedxUAhh2WB4L+lBQCgrie9+DIGSYEzA6DeXkB2xaPXY
h8Ur+O5fLMsJpQv/GBaXpvFnM9aduTbmbRnD7iVc5jdSMD41qbVQ2/S5b540Yknhp826Jk/yoOKF
i1nIBTQa7qjL0vJ2Vn2X0vMl+4Tw+0fi3jHTJWb/vpOS4RhxEVj5Ec0UUncyCyet6MfbKy65GW4I
ET7/+etI1WJmW9rcKUpqivQeKxo+nrROQcaRB/q+ztHch4vdP3ev/lSQKrANP3pxHQ4SkQOJUeZ9
+gjawUiy/o38n62Z1/S/Gs9R9K6jTMLAe7ZOpJ9ERnQiTQ7WqLedmqUH0iqGocIIPqatqL9nCxf/
SnFDhB7lgPGWtz83ryWL0BrfYHSn9Ob7NYiREC+gnfufACu1q8gYelcnBftAQwxPRUodgWOJ42s7
rqKcOqJF9wLJNpMg2VG6JTgRvnWYuoN1vDE6FD1zOKD2M+ankTmr+8usOhbhEbPkHJT9JKkE36fW
FGj0eJd41KT0z+Hx+Ro20nb+hYZw+rAMxETiFrvfrrKzvmA3vFGS8a72fwLFDrXOeALLS074LU7M
eqnE63T4MmT1efSnSod40pNZDLK7YhpUPKvsy0bpkspzZ6g9EStiN2OyzLhFTLiRwXIQhVwP8hxc
ajujqPwvb6+SL1f25DtaXuBvZS4mTVAqsC72VfHOUZbqBqvN5YZpzYJpyJcg5ZXghVwgUwih05Su
P6+pd/CIvjUn23FO9PzWfI+I/M7ahY6Ox/zW8pW8TI5C2FxF0atgEEtcn8gmPbwfbHXB9extFHEL
MoZYGte17oJl1g3o7UZMLv8F7EgpFoICgNTeNGJrFUMNxm/QERjwMdFVw/UDoljLVX8+MjIX88Xs
ZoNX8D+pnPynubh4qKyPhZgl89wEABSyQyDVh25UsvFCOsqls7c/PSV+U4ChPOVAiesomVgKWcGN
+eii7sGkRzNpNMarD6SRzOXyHToD+gHsXsXadfHbiltRnZHX3EBnq3iGobWXeS53iLp+8Dh1PcVz
UzyunvioG8lnAPFdzORDOxS8hExVLCcb8AGLfhinQBI8xsWXcXqlA/hvbUmPrXYok2EHOrCzj1cN
IV7bBECg59LlNiOWBtWqunK4M7zfVoIQcNcoRRM5JLljjaHpU0CEqobKs5xxx6wuZ1pCFpJlKINh
3Khegs3gjVElbohAgnVTnuYX3CXQCzUyoeiwA02dc4Ugb15J8gVxPOFrQRB5JaKfQLXzis7NU2iW
BDnF0NrXmhZpSpg5L9wrTpiy3LIkHztEOUL/ZXYQ36D5EMfJcwbKSs2Irc31jNshewKQIMMNi/UV
lj9jYEgEOoSjIq25LsVUCXWHErFQhSQJBfD4hHLBhvG/eTuKeU0tAS4g8WrQ3mWiY7SG48/eweo3
GVWRVDg0XIrgV8q5gY01hk3LFbhiOk5QQzGqSeCNLPptZEQMpyBOsYZEnNfJCUb/RMfPr1EeZG82
AiGGtXjyw5nA/WK1NaDecvLuNxJ1J2ss3VXbVm0iyxeLRZYsRY+wkHVPLNqfhPrem5XXrCxgnbQH
GzCfYXNSNTqk3onWSBSdRIyq9Oy2Fy9ygAgD1LDweukRTCfLRcFp6n3nG+ZNMvtc2Xkcz8QX+yFO
dgghEPfk781Oe3IoNwgPko5Bn6lyIHjaOmd83n62POIZ9JspGEJxaUxAmc5vLKCyWWHIrco0WvgN
5ziWM0k7LZqiIaqHgeNp9g0PfhZsPs6VZu76CvFa1SdKPK9tj2yOenT7KI5MusyPkC37N360hYxi
nNTI8y2u4oFTXE+39/UJffYIlcozJKK+erRmy0gAPfaOv3Sl3co+2EIjLA0wh2Y/E3c5kXhsfGcF
NV3TTYk3KUbvzNSgkyFLzOcAAZniQi/DYvAV8r7P6CWUiK4hOrZZCyGbNG6I9ae7hfoT1Yl9dLIQ
b1jpylo6fJ64Ik2TIihxSEpkmwH+XCJMvcX80K60Ak/5JxFp6bBJakoglGHWs0QIGttMlHlOGTXN
hU6tUNQ+oKRoEBPcHs6OUhgKc+vju0BALVAVOvTDA30HjxScKAcvUNAYrbgcDp7Hy1lj7sF4eFVN
wv3IiKCFZAKEr1deidoGGvDBCNT/SQy89hRU3aiHV3Z/hhUtvAOtbUhJSDiTcc5N5tLus0Rq8/6V
zr7APKU6+Y0l/W+TkubwBJ0rI4YoRT9SBdplYiZ+4bDHrSzi+4EgXbNygL9YMraqraRMh2niQ3i4
pWu4fjaWlFSfyugGaD1NEn9jJkia9V/j2ToqKjlQpUuA3afDOCn28/BOfUkCi53RTQ9coUV9Ny8L
5Wf4AeTHlzZLQpyhSVXfUjiJvxcmng6jOn0Ww5Eu0yZZ4c7FetIcOkRvFQvK0SY+n58+9mYjKVbC
0lQq9hF1IxBjd/8jIFXABJ21hBPCJfHvx/1Tcj+u5sGZN48xry2Q0yXcqkNEzeo7MlU2X8P8zsfs
TH1FqrrvDGVHhnfGkAUfROkhEDVInZUCnLWfj29OmAfxSM+ac/dMB6oqaiO5gkLRokZmf1Ej1LCk
Vqzd+p7C1rm5wqMWWxIQkD7KLqnd2p2MlbHQEOQJwi3R/1MgKAZXIKWQ8XMomjbi0bvPg0fv+cvK
MD8VJ7/xLYaaTDRg22+mtQ9joNDlG7877DUr9hkLJI/vFPkByCVdx6iTU/dicFgRhOSs/Q5AEu5B
ctc3b0Jmw/sHvAwQ5xUew2W7pXU/upT766EOQFNeCthkzeE+rG8sPII1Kzff/NObqhgcfB8iDbsW
HLaKY1j3EEHnj4p3AolMGc8sH+raCnBwTX74Ai8jTD42wABLs3XOwPsLyOHj8kdBLzDkr4WK3IVb
xUwjaPm+6MmjbJTpHHZqtGAKYrrCpzm9dAVraNp/4tCVQnb/aGjXZb0PAGu1RRUxtthVzMlRdEja
f8Wf0lDWmsEgcUGWJJURIJzum1U5Gu97SYBxX/rfFpK+LBr7n3TJlvbPPp1fGKrfC6b9K/Zl4YV9
p1sfgYLQlM3J+Yaf+dfgzORWX1iOndiydY7DG+DMt+mTtUQnJb5lhNEKYdLXEO07Fbvtff2kD5jT
urDYoDdSjZM4o/hmiF56O6BECQppYo0+zKvnJy1kXXoO4x3bDNLzykVhJEU97HdxHzHWZFkOy2Cx
dS50xnWwbARHwjkaRPu0axROLBwTrxiq6HLPYi74KtkI0kwDxOrFpZ1yibCcKtfiMQ0Gn9Ar2RVA
fw2m2cEoOCa/nXsrCtO5iUtUBU/FSdXkWJLB0eZL6M1Ootx4qIm3Vj7YCX8bbvIGeC0oS9EJIseE
WJLQzRO+6pFz1umEd49VXYkDaQCLt7IAw7r7Vp4cTL/ENi2UnlpWxye6yHksbVS+D0Pc/v5tEjkq
c8bPEcSsSDHTm7e5+wdWL/Dp5LkULQygybdykRLApSKg0j3lx+xmvX3KjtftTStjtxjPInN6ziAH
AMGxkH4lLi1Phlia+YWe7qeknUYes9+B2YjkkJKy5z8ModMueRrQMmOdteDlax7vVn4cAvvaQNC+
ETnDk69M44zekTQ+KvmhTJOPW+g7JerDL1PY8HjNPKazxDdhdwBnhecyeShUc00qMqahgidpH5mj
QhQrc+YIc/9kk2Sl1xJ/Pn/7bmEraOn4ohLdvWh80Vc3FcQzBnF4CLt+j0rADxINbQD/wtL+YM+d
aBLCd6VdhfNlMeZnYgRDXqqmUBngOMMgLTYKf2jrRBTFxvJ1VFyx3X9EtAxSyJ9EZUDQCZ5CF4SL
DwaRknt7wchHbpAOjSOAVd/E7gfyn/p7ZHbdeXuqLzlzm0A1tUvytUrY6yPggdfzQtSJ/RvDa1xa
TSGMRbe5HcLa0gLUcWZMBahVwzRwYFeFvbrNJg7vxwdeXr3HgwsMWRivwbkdT4S4cOEj2VIsHFxU
nQwwp+ZPjHzduWpjjYu3Lfw37ZzRPVUHzLM4E0e4z0mySdxk07k7RfAHL/PzJ8pQ+9SJ98+AuQ4d
mMzFie8vRQ/lycDkHNm90WdVjA1I0xv0yhRvzSdZ20GNyHji7lUegezatbROHA2Iadt3dvF7sXK0
tvlqF8VOyGk/bhLvSw2RDEr7t0SNwKzJZhvcEp3FSY8CjpAdI1+RCncsmbrENEQWwQBMiIQsJSfC
//ZFmzPfL5vHFtfVSQ+N5FhEEomj4HFrTDRPSIhSFhcAB/gyXGYUFkaNTIgWS15vFsuTCfZcRHBI
zIsy2pd0OUKxVocL70HW+QEnvNgZlQrWgwDFvynO9z50Ejpk96BQH0ZEbGwmZFhrDUCcBh0Qs+bd
MlvkeA5kAFMUoHAr5TmNYlbJKai39vPGGFlFZGeiv1QpWNT7+y6HX79huai4rsHiRqDRGpHZRTMj
6bbVGMhh/MWAKrwIFU8PVQEDCJ36u9yittgc8IBhfyZfMbmAVN7ZbYOwyABTfXaZWE9tcyG18Fwy
ZqJzxdkrdlSVjxxqIJ0Y1zFIF1jb0hATte5bfCiL+d9wmxuVleS7oLyCQZqMm0lt68l3s0aD+r78
KiH0dvheQsh4kmUSZnAmeqU9K9QWxAFDYnexOB2h/hT1365SLT1ZDeiKO2C1QJOzSGFLmmkLyN8G
9Bona0gUpB12NEKtbkBEYuZ7rETXqlKzo0wSqCE3nHDb0bQKPNJ1A5d1bOTzF3WBsLi6n5tfJ2PF
CknnRW0Hb0K+31YNZBMBQgLhPGqRhdg285UEDNX1UHHe4ZDio5Bm96hfte1+2DAhWSvNjhzsj+M9
njoyXW0npB/jm4ZVW1oVpHvhnRRfQl5eVIFFJHxMCl58mGfLbwyfGoWwFNsCg9LBTl5pi+yuBS3H
XauzG1xwvmOyjF5H3Qq06ncpTHXqyx9P56WOQEqWC+bfeWEKcp7rqaQDdKz0XTEzer2lTW31MSjs
nixSGqHQHu5qWKd7roL9B6GYFd9oe6pX0QBXD0OcrqtMvHySJHtiliEDHkvruNoDdR18gwkoy8iG
R7X8J7zwtbmjRZSQ6QaO+J6hVl7LCp83xZKr3Tey9n7uFVJ4f0g8LmhEuma+jGpJ9hljcT1cMG6o
3TVUlHkJIvvNtfN1xr+k43+g0b9xcMy1B9qgtdXO+vaBK5cemKaiGL66gsBYAqNMV408zLO6/Qxc
NBYw0OBiSogX8kgnySMxmFHn2hMcpcRG1c0QZnlUXkzb978lYKWzjXMo9Ui9mzcEDUI4YZRTVwnl
rUjVtPSIF26WxiONL4P+PJsAk+ee3bBVYjAFfHwyqw/qzm3Ar2QucDcQ6Mkok+u9GTpqD4OzIet+
9C2VcihoLEpqQKbD9mdvhClXrYLaV6IMrpKMOBPha8unnXFM10Qey+SXaOxn4WSyirl1BJmNzhu/
OtMyIe4VzByYuU0whg/F73lkGrRCfaoo7SrMnQw+vG4PGzq3AbWu9EQVXopJb2/cvsrBJRo0fqkz
WtYYdrqRiWOFo+fFVp0JR653IhQLNlNyBcf2/8j5FkMzVfIXS5zdmLL3gPNJoLs71KkLEFDT14IJ
dQrzvs5NYpKQaI1o6nvT0qizoPFoC8CH/355DrInnBtjP/hE67m4jXanCVul1NwqkGC99nwelonu
kEsdruWR4+421HWU/TjBUfhl5FjSj2AoVfy4ihb5aQiPNJ7I3eumkMMhxjtM7Z10z9UXpsSK60lC
7QSgzaQV2mwVcZN5IDmvsaKvsNIXGeupwADxr3s7ZONf7NKESTxxwfBrZhDpRHXqWSGdfpwFQwkU
Tsi+deBgGLHD9aG5DxiQIla/anATQVkgonPMJUSNsx7A8d3nSktLj/1He9gWLxlfWuJNwzIsCU0/
lbR5dJKd0fd32UrMMx/5j96TuifLChi/H/7l1ldCMGutBpiULrlgIHIsyTWenVZS+oFKNursOLYT
mJpH6qkuH8yWscKZE4Urd+5tbkja4rFeCoU6EE8RKDOfuqBxNaQRBh5WslZMQXZ730DpFr9RuNO+
6We+dpcdhQ4caYb7CWj57lpdyor+IW/8EzMXhE6vbMSLhUqEO+OZmYovnaorS6nMuQLfmiwex3ht
6DzvuYgRnRCsAH3qirEWId1nP8GLskziRn8/Z53h3LfMhxqg5f4XeY/mi4UAiBeEOdEgTr2z25kD
NVodk7qGYxStFkj9lk8Uuw6QU6XmDJrZexZDJmwuy4ia7JfcRW+V2SL+h9Pg8ImllHwffUoaLwLp
ZcSrBUNo1pwUfmKeh/vACsGTEitnColQuevaPmscgq7X5QJF3bOXpRIgF03U5u4suk/ymTzLVmcJ
1/f6ptTDwoybeDUW1ekuzGOzGMQgKtzw792j/XbWcg/lFwsYZNK3kCJ0SmA1zn3MfzCJrLs+bsYN
EcrH1OTKlRoukCg6k1LKxp23nQ3ecKj36ymWJ79aXi4LCbfMBUSclboGMzlNtbHqcSUQVDZVwKEA
LmgcqDoM6OcQDFnjJelVjTtVBw93XeTkzqlT64jqM4BZp3HqhJH9QFGz4b9HtgunDQYJJP3rU2Go
benKpk+64YpAfqQm05qCn+qUFkDLr1J2fHnTqMD/TI+Opr0SpUOMwlKXwWGc+vpVBgpa5wFlO+mM
8pUrKGrD9eV+eOZxuVVICjlE3l3sw2cSXGXYInJ7ryThRZ0iBnvAptCuEI/0G/uaJem+7+1tUntt
k7qw5DeD4KryA4xXz9lR46VGPjBDzQvkqixLinfJjsPgjE4GcW0ghBAoKdodtjgtrjkpQEOU8y6k
byCVLzPB14gOkFzsirKv3bJ1SZGOjUS6cSEi0PDpWjOFsRsRfwVRujg1eDrYrhaQWjV+ZXv+cDkL
9tZapB5k7AbMHFKWZgSIHGDLeMlNyCIhLLwuxhwzQ8o/IYLiEIAGIYGWzqnBrSG7vHfCm3DzsJQz
K8Lzhd7irXh9MtDJjPYc+mVA3OfU6TZZsAktVx0G2rnz7QGtaDd1v0wr96osdGra1iwgkNIk45Ln
3zdT1jp0lmA6qkiIkgwa8fq1Kt5mgf2cW7AsLNFwqcSxxV7a/V6PgaEyYYNt8eQdFt3WUDwWE3m8
G2ZiKGG1JcFItuShfYxuenxBKvuQdgr6FmhTOu996lvqXPTn2Vhp1udY5pVzOQE8eMsbQDq8F2f4
HN6Z+RKAaCoNOR7w7UVZUjSKiY/1QRhuWBFk7Kje8dWwUdndMhmHl6e9bC67mgikVzmNze5q4zwq
ddb4I+w2OVUtO+AlTNuJbxgdA1AtJNwyWpkn5H0DLWgPceHBqngK4o64d75yDkR+sZgzBitkGPSh
SrRHoG7mOV3gZpappablcX9lBilk91TW/4dHvNefJ2/KQatNeFyaC4Hw6L2lqIQF4WFrLzdPEy2Q
GQ6eq/xhHMO3DhHismiiMA/S6SfbGBu2t9cyURlGrFJIR1Yn/JYdRqNh6pFoazJrVVxNZK0F8gGF
gBT2d/fCs0Un8GbQmBVoV8fIwAUdtwTuGkXXp9y+GC1RRFTvDjM2RlMfXx+F/34w8DFCHbW8JxPA
tl1HJ418HThzqZk3o053xnhHZQlnVivXHZ9lxGC377GUJjIq2URjWfeKn/tQ30/DsmP4uc9lfZ5S
x0zuOyYp2duM3nDqplbKCSolHDPunRzMfz1AxMoAZKVKqML9rU8+vL7PHHsAJqk14dmjgdFNFSTe
vtA317MoLVFPNult/iQag510hLhWAP62NChO8C1wlPW6PYCW+rZzxZpLztiA53APkihyeknR5eJz
kdqRIBce3T1NblVZHRu2WGB+QGoxikhTESpt25TeqnOH/LCUS11nnEiKdzqAqwdBEmnb7Lq6XMjT
cwoWyBk3Tzh2fRUIytjeU/22OBp7LSXCxHvBh42xQoQm2vAKFgwmCSsAQDZkUUKATnz5X42pxCKt
VyU836FVGTH0l7prDoinWnOJz8ZF5sUzNiyjN7g1H2e+yhWSak7vNIxaJIATiPhU2Rb9AM+5ebEh
LzsRFXv6i82DAZks9NkN9Tq0buUiK2GXTTV/s45k3/Mp/BEMfIdilpMX2kFvSwPkc3Ttud2l2ic0
iL5RTNwKrwMKRjejK7scPvj/jkAoOH/JAbe2lj/wB26vkqbV8hBEqL/j2K2cR/EC5LLNK3UP9ogu
6sQqFmz9WBZJAh+pSNPKpdvHOHrresjors2EBV8PZOQzgBTq5JdLMSKWCmy4eTvF7ydiFX+3ZJDw
mkeyPf3Voar0R58YtYvmyPoxV4kUD/pePJYt+7tBw/ZkCEmiK8YF4kuFDGvp8NapM8O3RCX/rBIV
mscp6sagQwYFv7RUdmrgIakVOguir9Nud3hO53JukK6AHr/ILm+CBhp3C2815W3++QUlkeEnVESC
QGprAaTiFi+cwtFAhWPI3OCUFrA8oF9SxLxCZefX5DGl6YlLqjvwsQWOYJa7Ir3w0ufqaudeI3MK
oa5LureSOx0yimLepVk2VNuQF6mxH6J4/GDsFVV6KH1Cns71aaqksI2Lcf/S0D5cUQt0QYhLg5Z9
dV23LSsI1gxm/GNMUWtlLFp1KZosK5huPchammRmFvHVCK/MAFVYzSrUDqT1VixHpzShhTQ/sCOo
HbBVk6mZit4useFYM+VYJcKOBpYsJdGY2PfRHS/RuoIb98N+EqKGk1f10rJBuYyk+tn2kZftB18C
HZpO0jRpStftaQnLHvDTjb3X3zo3R0xfZsBuwUBVPRpvX20oKK7fpsbZ4QINr0aBY7RSVsU5uLJS
gcccesG4e9RMR4lF3Y1sXb1X/155KMggxgx/slKknuxS758TKVb5odL91YFOGunC3IKUMN36G5kP
4mL8BWF+qC1BirtBajs7IwcnEco7spBHmQ1cH4VWzPiIi+W2/ivAkXr/CvXqc8f0cq3D8wXkqY7g
jpQ/OdZFj0+ivAArGWV4IMUYOUVl4J7s0G90bekuNHY7WVgVa91q3o3ODc7clCdJzXD+R9ByxjJE
YI/2grDmslm7cIfbi2+U23bz0jaBS8qerrfLkPQaQO8ES+H36KdQUw4PNyhpgZHsb9UFrcpWKlE7
6Tn37BzSE9rBhKwfnl320dpCFQOGEtBNQSoPQ50Y1Jyj4OLZLQ5eV9+Xp2OPNnFkIjKnZhX3cnfj
yJehbMdW8oRI9VwlEMk9Vvg822HHOOEIw+6ivUCffz2vZL0ezf/iRQ9Wc+7oyYNnibk/RgIc3usG
uVIwB4radu2bfUKE45xldY9Td/hjU3lwSln6+Lphe3IA5qqb0sH++Nw7/ipJniR+GciIpKhWKf4T
IxXmAGRDsACFtrU0z/5xbse5NsPhxNbhVuVR76FM1rpWaQJX4MfEe7STHaSonuqo0loXV2IoLwIB
yUFlk0MNwC/45CHRncCSmbzgPUrXn4NEn5W/QnnccOM+gE6LOdMMITFEUOSjyksXy7BR/aCRlxW4
5uN3THYjtVV3OuiJ0fxbbPOqPesfbJlJduf1JysapF5R/QhcjNRS3BRK5CdlRsbf6YqxnHSzQpuR
1ktu3uDfCF8ccKja09GUyR9sEeAxs0A9FlYVYkiDsjHNvusc42yA5otYfMe9sxKFhzi8NpLPMedN
HL+k9ttgVrJAM2Wu32S0ju5o5xt8/QdWwUShgV8wF7nmPYaEbLwFOlfngfHlap7A2aX88r00MAHB
iOV4od3oSvRTkN0jUFI+ZksxqjSGYxkme7UrWhFJvA9chLuWGAm82SPJ4oe7k+yfVcsuc1lIigHx
cDaCRyjCzVYpkVkPGWu7TuaVNG91Vt7GmOs+VTbx+B5iIk45OdO3jTDYf95dEwLyLC3CDLXUTkkl
D4k/ePcjGLRwfQ+0SqNJij2T8SNdoH+ypwpuAJVOyofutyCV/fHkSChSpNqo5ZXeOD99PPJHj/Bp
f4oXSMCVPW9Ezmo/L3/qIZVn34a0//h16NxjoOX5y1tgqioUdIw02NIL8nKyk7tFPWYfKR/czaFV
AMuwUb3/IPQRrQQHZBjH1F9ZIxpNneEeb35+wlAM/QxUQwDfO6MJ5xQkKAiJ0u+4Pdt3BwlGbCC+
9qDMlx9Hr0wzwYqDH1hoxpf96NTmF5aYm8GZYSPEk/oDZn5r0nj2L8XKHj2goilVO2SIz6XyDPwF
AW82DLIPg2ER1+sp9snYiA+zIHJodanYYJEgNgqqgvduJW4wdZeYD4PJ30c31MgVs3dWHV8PGp00
TyrdXgdiGr5aRsxDD2YnltGWfFswCUheTIxuToOJfsRKsrPwQokLJNVra9PRkQ73m6dG0xIIQTAc
VCZ5cUmLvCVSNykWgWaOr6g/sfCeQkW3P8ZbVqTLk8sHnyi0XF+FDgQvRyF7AOafUDWyJBquYhKy
n1QzYlvwhDMNg2aLFVr48eTVh4rkuY9JtDMl6+qYUHZO/vOTZnoPATsM7cUT2QvqgrKwmMbhAby2
KxNi0mup/ALIwnJYvHJSJgacJL12B5MreI7EqjMP4yxYESSr3RLM2TUw6OrwFsZfwXlb9+ZCyYSG
QFaHku619AYy5u0AV3yGsLgO1W4sI+8PXwsowPZ3dJo7b2c1IeRA1JLt0uoaSiWJCtacC43oHRsb
reN/gig520+Lcg6mtgFY4YxwXdxPGKPyzNMw7BpeHV2gmVXAA7tgD8HVDe1DMBMT6SCZYAc3Z6dK
/az8BuKuA3dDjSIJFPFK+qwfzWb7APLyjqWTJHhpRtmhhXMPADFFWjITiVz5QtsqeWlIsvGpzRR2
cq54cku4+gRLgDCR9+6URAgkvaHpZ9ujS61qz9CKimzWReJW8MLYUgI08bxsDklCYbJvlVd3ozct
4Cs+RD2G+aySa0BwfERCIogL1gIAMTT2GZtCC/3lQnlDBDFoDf0GUj27UJKRsoc9OKlsjNG7GyfQ
o5OCNMg7CZda0Sq9nJjpE9DA3MrzFXxy2Cb4F/4DsCAdMdwyGcZYXBNB/rb3mN9iNHMWkasGSUVz
gN7aIhdgusB5iytPqP7JG98uswawTcHQsIqmb3e5VjmJ8afgppiKPJt9utZDgQPB0+AJjgjo9mFM
Be9BJr6IM8F7dDylx3SxRKJSJtxHUKbn6TWCuZL9Jpc+1T+8QFHutGC3D+hnzlgtycICiNXvOVpp
GdPAsaNWWZEv7bT+PZLVdsj2D5sn3t/yY49moRRRjMLEB/wL4E3hos34FBVxxPw2TzF6GCe6zqM1
62f7KZ4O9HFPEgdKPS5cKIj0ifPgSzrzqEQQrMCRtYt0iDbODtsNW54CRi+ErtgeUpd9/V2b2I98
r0bM3THBZPj2hWZ4BjsqeinGazgaxwwbybKtgJms1NZkHLsohlSiTeouOem1QUBN8Q4p7ChCYb2F
o/V2snyvzIYPrpHaT8QCxCRKxyg6jXiRtbTVHVS2EqjepyF/ufeuPZMmbYqQ5v42mdfSNAhqkj2i
+1dKX6xdubyslaNLDvb/BuwE4/jb8bEWbLxoQ9tkx4ywpYm3dLmKFAgVahcB1CHZnm2AMKc1J8ay
7LjrAlWSsKxL0StgFApPjKoUyPPoiobffUXkYmBrLfg8tkzi58SbNYP/nVYKS6RtmBtryXsT8ytA
VBWbNeMs/TQDX0XBs+puQz7GLJxYlnLrSTox1a/4iHd0S5cOP60mKDXan8mMRGY/jL1xArDmqUt2
7E6t2j7sEVBil8YMsFIg2k5+bilv212lmOpywGXsZNDCPPALU+Ags+YQX78BexuApeKb898LMS46
qeYmmLsSPeqyZoLvZ0knO56psHamDoXCV5b9XxVV0HTQy8QT70o7zaeY44aCq/YqiZX+qN7c+PdQ
0dGKYesb57vSrLPJ4CdcW+scpzULxJojegqcEoRBiEP7ULIuyPhgTw6j6jaC6naZrCCjBm69qzBm
/8JJsCNaz1JoOWXsoJRI7ijFrjr7J6SLA1tfjsRKTAyLruz+WxuqLsxJ0iJcspxzuXmmQEmKpL7M
tssfc/FEs09ZV9sF2j5NIdvRpdmWIjKCzOF+2rdexEv6DnwfnS8FwXk4xhukJOKIoW5ReWbD3kTd
0YTEIWVWDZbIVP773mQq6llqM3HA+xgj5Ifvy40qifbcYRr+R8tZFgMuXoO/vTbZd0tGwer4Y8Wt
2ECC8BdmZWLrsAzFd6N4H8kqdP241NNIKHfyoWGOXWHtQSE30KedWVePc65vy8EKIFVDrZIUcvyK
pW/e+yoo9hnsBBoW8nMMNfkJTSEGvxj2FIFhfZ+YBDmRkyKkh2w6w43LBEKhT25xNRokoEPvTVIj
TRFpiCfcy0fGBoW8WSiM/4xbdIwRtCwukhg+9x/D30ZGOblgwwCoJhG+GvYOyUBa53UT3XowosIY
O5VzuNk2Ju57yBuz6/0If0uFuUwSLBorW3PyqR0kzuv/r17ynUS3JP5HfqCdAdx1TF26gKnJ0s4d
qoFB8dSNaFO6dA7xRq9fsbOtOS3eciU8BdUbuQ3A9VS3nwsrCs/iOxHPSwXV6jN4iuV77Cycukp9
OcOtYD0+qNbbdX6aZt4z7XpkHdUjQiGDRBJJsgHS9hJyKD6fwQKmvn09PiHxEov27rf3bHd++to1
BaVZckCmK9JWJkGpEyf8fubEdOrO+CpVVzxiB2PshHe6JbQSoSNOHmWp/jNuo8kvHNfLfo9zrXXL
AgOseacYW7o45jTWcf/OCNCu03tcgZGQkAgqZSLLt439yBiDLKJlriM2WcN2jOOo5cahMrXoPif9
HPRcPeAQEhbmnDPwnESKn6PZ3qjqqVOWcul0IfBbBJVJcHwQKRMp5uTOaz6uqcSW6M2SHvuRCxqg
Y/IqF30lpHAm+KS2R8LM0E9Z+y1QKyX9+nc9f4mh4O9FNeDZC1yGxhRHcE509kcr1L884IA9AHuD
Wrj+BlcS46gkvypKPxISkLaPFZXNF38i3hmuHD3AFrrk0W1ds8LWv2i/h3mSPy7lsuqtAJbaEHlr
OUw/vurAjrJeGyEA4XebpVU5xnlJWckIwEpzqG3CXS/fh4LA59Kwpwv/+RiD2NdgMvzLUuvml7z0
FTJyZf8FbkMHdSgYEhuJyUkrIonpGZW9o5ubHiLYHKzAtgkv8lw/wcYwsipZTtvOuyapJZiCBX71
AZRvbu86VVnLGbEB9o9MHiS/A6/u35yraIBHOctoftGOYTd5CuTejvBkazwTqIoB0NxfAnBnWZ0n
tn70Knp7gOpmndubb8Y1xgJh9F5IZEpUnlf5KtrjLZANAkDze/CZrwlaiO2G2uIas8zfYnDn8R4C
oljnQdKh3U34fjpxTNIWWYXqQRR4unzNT5D8eeRqwyE9NMWG3l/XcVTHGdGD9eKhk+7NVDmJ/qNi
iz9m1kvGOQI8QwqStYZmCDEQaHaM4t5Y4uZRmFneV+izlb2RU4d5bqMZMVldsLEu2BDkIKPjkYX8
RxQJx5jyMcuaJ2TnnCdTrLVjO4bMF5C2RhUtrMq+iQmsMy6XWixa0CGBb61bFuifIG8xp0I+2PLH
WPqVfK38ZgsG8EfUk0KkXgftEhzyVgllVvNUARj+WXyNgDJ9N19uPG1BQOUBRggmNIlndffBG9ho
2aDDFVxO5BWWOU1B6cY93/IMaFskV8iu8vyg2hW73Ks08+KifD9qH9ff6S4NUtOLgX28D7Rdw0j2
APZiIYXT2QHZj4GH/5pHJ0r2GeFXOlrh/Ulq5DdEg3OrhDPDTLAfXBHT8R/8venDIQ+c8XHFyWhF
eMN5UfG/3b5ZI4iPoXhB3QZFhpHlALL1ZNKiD/9rHdgZBYPmYpw7GWEW8yWSOOsqFOpskqDrciF9
M0ARyEVs7v82OQs5/qeKa8+nBRWquhOliVAL+ecY08QwKGMxkkEIur/Nf1Hf/wVmgVTsN4LcOJGG
/LaueAgdvaGxquAn1O13qyjRWB+O12e+fg2iHNSLv1p/k+K0rAkfiTqDLi5qrdI752wnt7dKFZfL
1UeJZBpAiPrGiytYNLkQxEJnnP4FNK89rkuYgYOnEdPIx8h4/sWo5YnyPnsOeVSZUMvdOrfO7kYS
v+kdMppCbmdd3mVjto0/s1erXcqRKNrparn22tlG6YyaX1Vr80/rd65Rky0xEY4vI4OH8L/G6VcG
nf7ptAeblld2YIQ326H48EZvdlss1Y3VO8Ucprxtp94QjGgWTBbEFDIXEunywWy7s8wb2JwxIhjS
YkBo47bwC0IdIbPHUra/BAEXOqDDRz6ndILlGBxz3o4HuIYNZVB3Y+CB+e9AvxGtdZWvwJ5KM+Bd
LtG0h5ajq+dyEKYJ7rwDhMt/JGXiwSgMFsR5ALOQ2Joa4/SbyaMPgxl9+TZcaQhdoAzdDOIiD/HZ
YT9pVpJ93ZqGzo7X/b3S18tMW2Q6S5TIzRVp4ZrwX/mQybq+FdOobSo18emzQXYb9i2KLJLSEC+w
egBdnlgTS35EkN22LtkgRruFcotBwHTW+Gdrqd9zsevnZ8JCMsNNlaPzlqlvJQ+YUjYFrb/DUT7l
lWsKW3V6KjtxyomPbiMNkGIyTF4io0EpQ+A6OUhLjr47fUIibzQKgeb2lLKP+GJXwozFaPgCNseV
3h3k7meMEpdi4p1P9uGQM6RmorMDw0cj4c6SaCudGig/YcqOu0/SDGHv6Hs2oC1tFw3J1QV+nWB7
nYVzx7R7DCJMde5Q6vmHjxkXaYIqO8UYbLxivLbtOsWe/Gr1mIG+i0myrM2GkQ+ZFUUZ9q/cDVhF
HbwC316Te4MBdEUVwSW8v37aaebkvTv/g6Bkk/2KdgeLnR/0rt4Fm0w2f3V4qNmCELWT5QklfTk9
NnF7M92eXTEj6/Y33saysYptxb3kGDRzKoQidxEdlAX3stymL86xA7z2PoRS01X6bLMGCIspRjtu
TvX91V3rLEWJ5McLQnzaZuil60BEenpR3w8ipl8kcyOcFagWRZapSUwOD7BnYU0CYhvbAcmjog51
KZZLWWiDU4Njt2HhvxOHN42TZYQjR0XXXvIjDuu6dSpV+EslQMnEfFPIVY6tyQjR0A09B2Lu2lYm
fSUX5mgPTsit8yLvrWXXqaHP1GaPCrbVAugmdG78B+5nX1itosDTiYN1eQYhzF15s7AzxyMK27tS
3Xf+vqMuaQUSLve2PVatJMOhL846kRFzqJ7d+/lH/nuij1j7xJcqyUKK4YVdZm+cOnSDZDDUS3Vf
UbFPhGpIG7PXMKeiQx7cgwmKrpG0aUrC2ttWr0LxlSFlAcQaHdrcZptbtDc7lVbrtqA/wBwg4X6p
+4NVD0XZhG5IUuGaCL+3KcJRfZQ7Xgs8TSWh5q9yE6R1Fs0oKWXI/DyrOUUcbbMG8B2esOZoMVkB
eLhF1oJMrmXkFntIft6umuaWm8EtqYft0cPEQR+iyu52ScixSCO9NyRCZKgXoB1c1sqd26RxrkH+
SkB68ZVhnjh3Svcdbhqt5yXjeQEGeXeJUleKfUXsYimAhSMXvH13Avv2p27c4GwbD0Rtxff1UnRP
nGJoLauYeB13Lnj9jg6xSAGUdk5aX7TWXhYM+BwABhez8bXLSSl9gdJcrlyCtpUmfMGmql8T1Hh0
V6usBUqev5p57W3CP5ob0ihHtycm6o22ZEXlX5yy2TJR7QBnYCHpkyT0RC1m7SQrpHglEk3hHEU2
kSQEggIAFOX6H32VEsVUpDRNWRgKG5mWFQhMXPYR9qhBiaCBhsueEdS/8/tGhWfwE5VsFT1DF2bV
zjrAYSpJtafqUkSivy2dq/dNKeUIHsyfTiTIARDzIMI6vTkLHrf1GEqujjHcYz6FHKFqkR+C3TXN
uZpTUTq1hFDRZtjSy78k6ijEtKhpMaBiajoVaTiZr8IfJ3q8ckDHJ45TaVZ2f/8LS2vNLc/p7ZIA
IVzwkYX/wTiSRy54/x42Dhmi71pDrQiZYH8qX9de2tIe1G/b37XSoHeqWkXsRhxm6x7xK4nJfOK0
YUjKfW0WAK+WJwsbuxCsms03ThMCNbTxeVAMzfK+DlxC9UtQM63l5hrFdwZ3hjMBQTo5l5mDH6bi
ZQiQZJMNbRMlL0btrgBUG/ObYJz5hST1pzlOa66gHrGlV0KJgyvsmlqwWLfHGxR4T7aOYhfAGJXC
8fm0YRRopAFy2k8UcCaNVtC3HFHAeBAbX6kaYNAGmkB990p3YDmzinoX2YtjId1a7MRABHRPAFlU
YVjss0kebIJrw91gSSjp79cJixSNekypQmU+xrrcQ7FUH3hYO5l4bxcqfP+D+LnMHFAxs33cql/O
zBdaL+ILFi4fRg3vhnpBLPM8RY/RK0S1GTT6befUOi+EAso+ZuHLfFUIZQqEuLmBJTHJlAoADOgt
8ekhtbe37jMPiFGOIQZpW5PHq1LldnD6Vh+lQkShYr6HL1c3Xqli+cvyjqnK6EDgAPDByo4CxZsK
sHaOiX2nr+PdGwLuHfV6YdZjafjO0yqrOOjo1jZDsSoj5Zcl+dd+8UUb+sO70deuxd6+dH/qn7SP
axZ7kIoT+/5S0cdJ0G79B1rBhrBdhB8EmAJH2g50nIBPZNWjtpyxsCDuw+aMS9tlN2dwAXWyyaP6
QtQgOv2lFf0OiVbzEZ6qNycU8ilszyX8QxU1mshRPJXBOqlI4Po+bye6IooUpN4NixC7k9MH7Pq2
bx9Fy5hN+rSfWsB7fT+Gl6p5HQl/XiR7FbFUDthr2cjvgX9E+VVh2BriMfkNzVuW6Eq1GbF+mpJ+
xMeBbYwob920KDZbVup0GY9ZapRISCkbGQXP0S6v4+AaZYZLMtlE5LR3Tand3GmDbh54WdJAVsD8
Q1BX7r2MXGDXS90J8h62VdJOaDd0g2jfXQTCdUwlWwo/BiJhQFvk659Iwi+SainqPQlc176FrZxu
fO8OPS4zWZ8J47jCZ1/oAg9oI0mcCn6h8Nn/fB7nwBB3EhRVXo04faJO3XUKsW4mikTciUsJrClg
P6bPU9ZSc1LKIF6UYagFiDUHsTN8s4kfed3zZoM8iiarvMBWZzbqozPrOAefFLM1EF/4dWvQjkBf
dZdDPoUOcHzY7eEoiC7dSJx4NbVINfk5qGj9uvzYrwMBM+ZmmOyoOphyiIeCbH3Cfi/WVuvjVEaS
qT+GocFGvg45WygKHerfmNEAYuYOVHujufqCdepNcXfI5lxz3UKx+ifIcJqurZ9YwmhJTUWw1M0Y
m3u72l+unaYx9zDEgygl1bJ444bQ3NTNcE/0UcDzHo7hA0vVHKTtmRxtrUVHvcrmV4PT1NQaaWCv
pPCYtMqFpEKoPFNpF7RW2MsRoxgMInKX0ckSeWRaCWh3shxn2SSPliHFhpUu2/nE3zUeBReBlVXb
+5rI4sACQgf6CPoTGo2l0v10wcLSBhzi+eTvCZsFi6yKeInWo1JsHf3oDGEPZzFcMmjhNIP5x9s0
ASQSA6/f33ZTfyNZox26ne7KEk1ovV4AZ6Ytrp/aJytrvPCi0tm051E6rpCPHRvv81Nv0BIP78Xq
RRoKT2TbgqwSPAtpe323+Ij1egfxkT6u/MgEpsAWJaiNmvaKnvOO+FJtm8UknhK7vZgiGO//HjuI
mhfXyiufNETQS4MOuLKlQohjcTE8I3Qr8mm3x6rOXop4BBTJGDPjtDuxd2N+Um1RwP0AHAo5RQTU
Bj+djkRJz58YxVPpAPRc6B+ls2v8bzVMJ7EZ7g1mX5OsUVpNGG5MHAdfNzgst6/tJddNYfuVNyo/
iOKZrewMaINR44f5NeltuwlgmZzywzWUMMUHb2jHOmfiPl9yP055UZnM42kMSxCxNXzaDnRxKdzv
LMPTJu+ypC3a/dHsES4oM3i4wE3mKhNGWGZafYJM0y2K6ZJ185ZKBBkee4xa8OHGVICCbsi0KAI+
OgDPwU/ABaFeQMnlRtHaEJT79XBGxrtLkRHQARba1+0JjQhFj9tam+7GYvu0dlPWy/xUPxwNPV30
h+J08T1QXTgbKBez4Uki4BAQke5JqUIUhIcZP+jNQ4D/+6JuimDI3+7ZnZExUyaQ0r3tzqw9V5mC
MYOoTMnp25Ye8C2zMeIOs0yyeCSE7sdDK4eedHzttLFaIEMwsiNc+BBbp2ksmXOhs08N2gU4X5xJ
w1JQi/4EY2YDqw3+wpWuFytoPZPVNRjSjktE9q6/N5w/tEAw+sd/7U5dsfU3+zWYFczr6XBMO+ye
jApXbiiYqnhfjf/ltXdxF3AHwmjiCuA6A1YFLrsPWPvS8wp35Ct6NgMKF9QTOPdMyK0ymg6zp1He
pP+QZzdtSu15VvgQfN89WcIJkF0EWTfsoj12ObN5appC1KYc6Ym+y33WXqINt/a0Ap6TNTy0n833
LEXD01/MlOELO+tdW9Ne17PXA+kYJMsEAUHmbQkyirI2d2kePq1SI0K2r36z3EbUaMcVRWkbNkXl
NLj1e82idro5f3UhUoS0X9KAveD9F0+59y7r+YqugqnihxU1eyhvK0rViFUoVdNTsgakPODQEZTj
BxvqvNKg0wcGxSjkpmhsiUc/vai7t00a6upg2fDc6rwIVFKS2LUNNu3EgsS4JHcnxf/8CGtpte9h
/x0aERj5FuydPA70f+D6HRODJm56+rNLsOWoQnb9fUYHs2Cb9QO9zzvjMaxzOiUIB6iX3KQCnFvF
tH9FeIR9jVyg2xBqaJCFSj7VwF3bT0jSdtlsEKwU58suDlmSY6VelXv+t5JJGZAdEBBhjoFxY/S3
CPrLfiqzT1aAQ78q90lGT4QFvGOycpB0E/yP5h0g4sTTqK3KMGHJUX9+TF67kAdcft+JHlo3hYNL
P8H3vk6mbehu/iCFElE5uFX20zA2nOTruYSQlUI7sj5QOIWSJwis9yFw1RGKBBVVQ8y+TYCgzDYA
ZYgW16oOPYh7PVsaPne/vovCNoHfdruH5Voc3drAQQjBZB/0KN2Qv3djkb+u5mZ9W6/H87txocUG
3Im8qPWB7llzWwoLnzqUi8PCcNjLpW+SPLPdZ2dwMXNqLRXaBmaE1/2CHhy8jK8S8GWwJVwmlNFW
UAyIW3wJr6Matm/dLb1HnTl+cKp+I45zh2rj0WRZQd5f0mNA04nytqjW23fbCVz00+jwWXiHdmFf
WiAEC4ZBTeTX8S4WJbpLS/d6/3Ofbo5uCf8E3DrcOrNW5uTEt3JNM4brhSxYe2FGr25KSRoWOBHE
rcshPnu9sCc7m+riy5zVLa3bsbfUxLElRTFjOlH6POISjuPxp6O69IUfrQP6NA996kaL/mWd87BO
h+VuH4wAzY00B8kpq9dOTIaCfZiyR8fKoOtuZpCHw9cSReoeis31cBHSdhTnPrUC64njx1Hmgp/f
Xlfu7ewaIlhTU9XaRUtuFjLpsr2vKb3Ck3fdlN0vBxz45XO+CqApBuT6jlcubQDRcB6PzeIpwGgd
LPWnG3cQbCF5YDQVeFB/u0UFyC092HkUsuAAPmuVgsXPLmivKrPtY8h25X5ljQZ4JnYZ8qdARgie
qsIt0bCNY0MXUwXvUJMqhyf269JTARW5v0QM9g1BMontVUUoN9gQWdUzizkU1RvL0WjbDE4PgHp9
qnLsjW4xCrdJ54Qo5kGqBzhfz+7WSSxIQqe+uly4dBD2sjgcN40lUDABENK1s8DTOoZ6WOReT3VB
A4N5L+RTW8MRj2s0/cuHBqkYy8Nqabe4mNadjYGGaiu1afyA2HLxhA4CIdkhyiQ6Jw3oq6+Od4RT
ehUwteA9FOlf1xJm5pxHmil79MnZdJtCPokPNzFMiIuL6AjsYCcTFQpPore35Q2KLC3AiiY29KTF
FnA+agsqp1BeWH+fm810ReeLSRda6En3JlWu5asw1lM9/7J0gW/En1QhrLt9KH807/tAZ7ZNkhem
rWOL2b5ZbHw8sKWx47WA/5RbDvADthVMqeRSfEpalYLPC/bWYlyhV1VDXNmdocse5OxYjJBnap1z
87OfowaYIQPfbixvFjdiGZm1LPCrNl3746ZED0pzFocJj0mH7lC+7dAzatgchxbbWM2GFiANgy5p
Dhdyjznnsw4+FB0WHYNihwAPHlsFRYe/6UR/ji9alFR6b7/Uv7eXQ3crE8+W/8pxTSFCG4W4s4tf
ARyLjgWzKJGqgV4u8496Pu1rv++lF04tGnWliWi+rHr0EEsmMww2+25nabDqtBbJp/AHZrZ4z3yq
Cw/LEnFRGHtEgxDAeWeVupMbNluG5q3/92wN+Td+NGS/A6aZrNYZI10TnbVjPDxG3qsTYgJ4BfCA
4i+FWHieL3mFWMCXDOYbyzfrfnPLa1xZ0vH+N5T6/2h7Za2xTlcJYFLz87G9etcZcjGYaVAaEw1r
zKltW8RzKio/v6IGdZYeCErylXQfBSvr9pxUl766999Q1zDt+5/Ci8fs4bJPVBhj4frdOTSf+e/p
pRJINaE8zkn9PfPCVJJtzNBeAWe0tOxEnEyqkEiQr4cTkkDPLj8EZcPadX2aOzvibJMJ4TiHfFCf
ikSYlqTYyXWw1gXcPaHkmH6r+00r3nbV6S90CvOGBOBfHdHkp4/nuR+CpR3TYna2ZVfLxzgHI/Rm
rBY8/+RMLUpv9pL57LQfrvyOu8odedtIP/MzEmJKMnvOzUv4cttUyNykBglR3JPErshm1El7wUUE
7BaZDUkjEvdXRy3Yz1eONiBf6a0F07HM3dyMkbEfFTwBHNDYevvGs6ptnQexaux2hMuO8G8KiSFF
65NtEYyXQ2gIbqAuDzH8dacvudtfFwU6Q5pf3wMY54B2uM2y4Nx36GW1RTq2mBIk9JNAL3DWjB6x
a/IASiUCCFOs5Mih+od18pFojIlaa2VzF1Nb448CNWy/nmM8KYlz1Xh0zMh0sUud26S7hVdugXhC
NdveOqY4BeDBndExi8QJoM9AnZKJS2opweo7g0QT4AQL3umoOlRP9mOlsIw1500MZkEyPSyecMe6
GCq4DM2fuwBff31z8KyAkypNo0GVnnsw8cQQVWOtDueB4uGUMYCwwwAIAFfRTFl/IG819R9fF4hy
sYb3s3i05iNetGb+moiPPtR7CNb+0bZsKGKoreKbkjjjoxV3Y9bB3PQ0ZE+Y8HxfEuogcK1iYLav
vQLXkX5fkqz4X0cJXM7eY6cMDV4rlJaT85lyjJfjxCqBFHGumkjJzizvX+8ht50nx5wePODzcUyX
MQWs/hj4a+nwl7GO5jYvnujNmaecN/oyt+vFj8od03AH3KpNQtMmTlybwD3viSfgsu5SmudBujjN
NOU+Ixi8wHcemtsEUEmzZGc4j/3M/8ebeKgodVEglUEJch1MAcfwxMU6WhuBj/FTODMPc77/zkKB
i9HDi945qP1pc3MiC8nRvPG4kCke//QeEP9XK5itSvAZl8nTQDGcnql98AoWSSlb4NY8qH1G3b4O
rhWiWEXnPWwUS1MAHlK5iNEtN100WdkZnyq0CqN5tATlVEQYP044PQQwhhB/qZkne+kXzP0vnbTb
tgx84g67DrofHaHjX71MGdhASgeq6+iSHYJnslSxFCWDM36ohtPoAxvfEnXWh9IV06mOaJM5nC2I
lcYnSWX8s8cSFwafpevO4qlu9dnoSYTih5gbPc1/kmGCM0uEuznTBLoJObuRmo/V6M10rh+dcQMl
5kgslgGv6bYcsDKdvgqT9BJ+6F3rQjrZpQh4aES81eaGcbQ1RWgJbgDQmeqYKUx5/MM2HW+SEDva
qRTMln1PslsK8NED/2A6+8ABJUFFCbKZzuFHYq8XZP2jtAGJ0auNr3424LWHGAT6AkALSV7UqOTu
lITy/D7XTBRW0bnZHkfTVHchkvjvxVHQESdP/Ca/LA5WwaSoaEXIi7LMnI9ZnfMVJ9UKE20CL6Mj
Q+W7Ov9SZlEDz50F54iNbq9qZAhFtQAojMv/bVc/t+etxBryRpxUPX+7vE9lYu6OKqxnVzT+wJ5/
059s3GG5xHAr4vzktzgjTvXLhSdcGLTBXW4qYogbW6UqaZJ/pHWV5MwEi2vyC1XS2HSKUscbSwRa
lgZYwsK7uXok9w9UkYEy3yA6KSfMtY+tgLJKf0YwZkcXKbkj+Hzs+uoIRzBxzgtc9m/Lb5hKvfsY
Z3k8Jji5pD9ORTczQZZXYKMp9idGkd0OkjLmJx3hIsRQnQH0T2zWI+MAKeNRg2XYI8l2AclMwncY
J9zd/m+2V/CTABeW2EobKClydOmbsAZXZnin48ywMKa1K33fZzzgzoY/3CwNEC4R0m8RllyMLPtf
2uHM/QRZN9Zy0cQnrCUHJJ9SooqRYADZSJhRB+FSPrmtAd4w3hKcTIWysT/GV8gXZkCUSV01oWiI
1Z1kJdgSC/seJBp9WgLPTdGP+E46rNZrMvc/dVMzymBroNu/xaC3jQ0vuwAtXxFFHMNYGct1/D6u
ZygY17CToRsxfucR979LJ9NifM7USVKTj1dLSnGcxuXc/kMMpmCMpj5zH2rytVzD4pJbOJePxYZ+
KnIwAk08o3w/w6VNfcDPJoJTvSLe01LAw1fqHivGY73fBpPE2drxsRRXdOZvcZGoriux5P1jhYvg
Ba/8gaFGKWVGQYeFlWJzog0ShNlDtS2yIbYqub+vkRp2irvo3r1yv6RNMoiCEWB+LOe8JAaEYUVH
qFsxqzPv6xm6V+ejCS507HKvktTmvt8Kh2DR0l6eQerZHb5Vhr8aJ0+GrJldyD6CuOIgxL6i7apP
VxVczYvHcW/4Kp2HgXMf/qdVQZglssAN8wHkna6FLaKNUTK7icYrdV9kYY1m72FFJVVSMtcRdTbQ
9uucjq6pef7VehfoembUHAO6WdW+LPegEqJ+7dHxxTppg0C0mhWrGwaoAW2LrqjlH2b1Eq70S64K
maPudBVoqlAA9qcYKXFNTe/x+tzfHbzgY4Tiy+GdqQQYDGWnwvJWo0AtcnCSaZrX6t15Xv8mGoIQ
rufNcL3CkWp/2nWC9L3TV50yYc4knQ8dcWtDOQwc+/jJtlwsfaZLVk7RvUI6q+yolWMYwnRXvDiO
mpiaBZDl90RFtlMOpPYc1+DRAQxshvGaLrYl/9TNTZuxPB6ZDxYAKbqSsxUuDsLbOjrw24515nm0
WU2SV09Qv3nwONyeQ8pSfsBAFhXXxhKCPsNkz/2SdAq/Ep2w7HQuCOl6xZFl+7zbXB8TjUcj++LA
KfpTKW6yCUXXT2xHn0udtZUygFage6Y0+0DTHfiAp7QVj/bcEJ2pqVRxJT6N45TpoRpgByPhLPa+
ZAcSvZLy7VvrsViE6XRM9GseM5OiXkHIDfwROKMV7R06OWbqBkzwEA22NKZh6XUY0IvO5U7oGTOJ
z9L8CQWGHpGP6drA2aqhn94KkJEsujdcssCcDH1+R4Jn/D4fO4Po4s4KzSR/oHck2qu05V2JpqJk
Ib85Ql5U6jdcx5Yqy2PZl04CgHl/oCxzwvCnHrhOHv7ykwJor0YMpedoSmbt1mUWy2ZNNRGKq0fx
SqiUT02jsC9iTdoNKtf/2Pviz3ZFBH5B1/kRyJnfrVTbD0a74E6dWmJ/R1bHYMtt3dUzWGIPuCWH
OCZ2YNfII0zjVi++NvDMuvcJcE9FLC0a87E1wFNryMYymtH94+sOqTvpiLwfe2n2cUEkykFKxU8o
X2zcSJ1x/me1nMfQV4qq/ra4zejc1jl0kJyNXVDhAigg+R88f5O2ExTfDPCbNxuzANFQBvnG9iFr
UMnnKfGlX7ccKY0FVj8y83nCi0ug1Ne2W6kfPTkVBlfObx9vbPqs1lYmgyqxkPlug6umz562hub6
vSkKg6C+EJ53+gJMeukRQxAgKqI9mkb/E1yc4R7/030iKn9xsW+I6h28i3lOszdcgdVYnsMhDvxn
0A75NyiXYb7z/2bWT6SjIaYwXEzQIlRr3jy+O01ZCBeLkFDXPNRH3YIRhcTzNYv84JzitgdGY8OO
rGkcVYVtn5yMM2IYv3QG0rZMQdCorg+41JjA0nDvdhbb70oHVJUvpltHxvW0jdlK7NHDvIm++/pR
0TPRC+ElFUZZPk09wizWK7CH5yDDrnzM0zcJMvzu7fQ6IZELuH1rabzJiigMzxRvvxyHs7UR74lY
BGqTySa7MXdEz7hZpbFyOhm6hViuBI6cryz1qU90vsQrVrLR4lof74z/9Reic7XckOr4PxMDbUli
WR6PZuCwLk4jEAynuZ/BjEcSv54niV6pfNnoYFvMMWKTIn8LsFQjj88giO4xX8tlIQIr5pVVkzPy
26mXpb8me1Swu0RYdWvzg9c6fPPohX3QihkGhXavi0reMgYrvvRKTPGj75Itm501j1W+yaZjCeaf
MtBKjeBCr4wRwXh8bzryjTqadvqcrSTbhGz0IqxVddT0igFjZCRpfz+OW4Bue0BN7x2iUXIvYpef
GlP0Oral4C3JfIcvBw/A37k2RO7+C7TWWCSFJ1grvlxvtP6hYz/xi7ZPHsUKaJQo2kCNxc0MWa8w
OFfNCf+afGDXDpt7gEHuAE4E2rvlYhfEafsDMFu3xA9L2uxWbzesSid9pLtbTVFcPqbLeboVDvik
K25/kKdb36MRvXtMGCiXlmuh/xFofPPDYeHc+cpMlQ7crZraeIjBl0jGthUZNfKI3OZ5UhRzannR
bNLgxC2qGhINlOLVM+M3rWa/7+I0Nwc2iE9cJAmD3MohnWdCkBug8oCGMsZNbW/5be7bQ3STgNWC
WMrRLZrZruMfJOUBxJQ8VGhJiGbNFnIoOJ4TFi1BDLmbLUr22/iSyP/R5dIvcaCiU7w7OKGDclrr
rLdbc4yft1G5clnEWaugqxfdDdFrf7J8VxAsQMSC0+9n90yoQuBIcxqA5BSVogKqTRVqs4I9FPna
e6cHFrcoNIs48seZ5zUD40xPl/uj+tYZ0Aib/dpt5wFmbu+MmrjqtLi3H8Mt7vUTeoFMxDWr+swS
UPS8fZyAbCcHxiYsV0pgtDw2B7H+KkHURYMMeEJ3+4PxMOc40HMZme8Q143I+pVNDZQbSIqbA6tf
8TAwe5g8S8/BQoAtrLQD995lM888wVIcIhSXJaHH+A4wIwSbwGWod4lfMJSdfhM5V+ti6Bu/pqII
JZVQ2W6iUDXi7RjVrsDe/rguztOQcn3tztv2uMegoI8vXJDiWLlUSjFA4JEczBpOJbGXHbWlNpN2
Tordjmb8zQ+cSyM9cUkiejjcON4mIpP4PA9haBXHGhMku0MA9xePljUq4t6m44uZVBwAKNXYv7Ps
8RbVwgRLIXtui1agjY2GxZ7PRGNiOH4zCF+n/Cyt5GMUw+HExhLmmHZv47MhHJSEm/ZARjCESE8g
U9+Yjo2IcfgnUI0udz6SqxOhRTIH0tmXZ9n576yPGRR713LlJzj7bMR8U2U2cOCuotb4aCj7gD02
c2AyOJvIpKFEPeEfYSCiTIeKP+2MBiGeQ1EsLNAvSClO8SnGlet/5qIX8XfgAhAV88bZyhLEtAg4
KcCBoBIIN5TDty4KLTs/lfcF71hGZ+CAcSSMVoX9LiKPkAbAolmSU8sCwKP/W6lY2eWFJyiGzYKi
pHw4BLxOP4xMlFLQiJZuHUUwjuyQ4uJbd1kiLC9Vz3Cv0MASh63sQbaOEmXRMLz5Ly1IVo2jbVzE
lCj8V0c/0RA52XMWatpxhas7AYLn9eX6MgWr78lFH1M9lr9n3aTEr36OPlR8+qAIcUs9Baa5Tkzr
0ro4KfjXJogO7IMm6H9WT7fbhVL2nuvffLSZlB5NUrAZOUXpX2k/EHlo1lwb/1odBoLc8lquMCTR
87zAM8nLLBNs6JNsuiaprwQ71+brNZJIxluiWzKfodc4cOw/vKVh7RHr/3Ttu98rSo5chIWpmdkP
YEuNCA3f2Nnnfx1SB1Zeo+9CcI+8ezIw2RxWdUr9khWKbzj4kz522TfIGuvLNIZG7EMoJBVT1ORf
VNnXP65zF2HyGZGCRS7XfwHk4llircyiXFQHh1wUGTYT1N44bG8vzlEk/MdAABcdADMofk2o+61L
AgpjpEWYURd/2U/26xqeX/JnHWyR3fNdi97itWcpFK6M4BZH9oHTYr9zPABmMGMUz2Sya0Km050H
4swZdbAJibcMMUwI9RshqqM65wAhKXJ/tQxtWmTYoz6I59ykQDFjJDcapnAJZhgYQzK29BVjjwjt
42qINkAF6nYMRv74d/XDd8CXZdTn6iXqco4DW6/nsK6KtwNf+m3PNclSSYKcABccFziVs8HCQHmn
HWn8W22jjY0twNAAr+E9GfqRNA1D2xWSZ/n9Mf6gUOaoegmG/55wEBC+AAAmyaPqQH8UgaNipORn
PdAy8mj+cmXJp/QvBkp1I+VxJJ0yb1S4/naO77ErRc8hky++YZVvxgf5LqAMvAk8ygYW5bZn/gno
G02zLyF7X8BMQnYPQzlrhOIfisvgyMg6OM0DMWArAaokOytjgp7GU4jFxQKggSpde9lPLSVHUA4g
QXXJR64AvcmXT959Os1Op0hOE08mPHy8j7LDnIqoNfPN+6t05FqQLw2uklK2SIPqekPu6nGyPTz9
C10mK6TY6XWvFdNx4qigdEImjcHbsZyr6HZeU1LA2yKKTTHLDe/FA4/iV7PiTW3degXPVpaaBsSm
vJlRR2WAUijs9F/86PlanUm7+R9c9V66+cphdEqc3v6rlVMeTCcG7Ho1LnC+1xy02ML5tS6cqH1K
FpI9WJAOc3MMyzP+j5BsoLV9HARV61OXL4MLSHTneNXhWkdGGCbfnNFyZSFH5k2wGRxDpC99m0pH
O8IvXGSQqbq0CGaRPvsa7LEBEc5330UtjasdQgWPTNukHUt85t+0oiLZnRMeVVMkz4Rj2e/1V9f4
X7wQxTpgaoywBBg4xtWZIR0ZGcz1UN5KiqXkmybTYbRlz0h/nk7odAL5otZip2sYnO6RJie1i5SA
ikhJBPWggJ4KBO4CaANKCwKFs0/Jor2WVZoEntQ7S0RL92IdWZFhFff+bibTd0h64G0FbYz6Bssu
p6mAYkdApo2PUkty0b4dfBKqrrFtSOMC+hhTIo7Xy+3Lfum4tYNvXzLyM9xyvFGUyZPeVgrJNIVg
WXqgw8Ob7NgkVXlsrBLFJNIVZhOeXf1IEO1Yl1FNZ/uovwCKxgGxRl2K3Z7eKx+7f1X4jG3KJkqd
31SpbAIBoHrIzMzMvyvF1p9e5ShvlIeG7jQ+TLtm8nYRbJvGAf5NAlrcoYQDZwyw2IeChK41Vj0K
kU4YdsS06JrtJzvyjrm5L1PbWLNiE30Ur6G10cFgjVahxSpm37FeZ9cQnTilIIGNZxJtnZFUOB8m
30JQpPrn9o4+LOZOcwyrhIzCih2PmGR6WuFe1U+JyeAvI2vA+NHV/m2x5/7H3k1pNgB3Lf9dUQ3w
qrzQIIp9i28SG14tzABMVf4nY9nUDJPrGh1eVyU5/D/3bhoYVKN3Wl7f1IBXWCL0YwIKMlj1sVwJ
6Ufy9QHy5pl8butsdtQU5Pu9lXy6P8Zxd8CD3M1I9oubzWjmhzDdOV21OzhY5wJ+EhySBAxJw/Ta
2A6CtVCFugy6HuEObt/g2EfzX23fFi90gx7tOfRrBa6T9DvvRmt9YAi0JzeE1WgYPMsQmsOq0y8T
AEfdiTuJlO+Tc10V38uHsWgx4DNKw6PkvHwxvJH3g065VFyPkHi8g7lcMXUUy84+ucL8QjlrQd87
vDdITroGNxz0xcBANBdXIFiYCFW+m1+MCXeWudlh/Rwfa/5TOAWSpFBd1oKbzN5l1VcOFpppKOlj
mEVyGFxp6H0u27oqQGMcwWUtX2qqCfMHsaIJzwlMzQXAF+qcIc0e2EUxWEOSSSF1zyvBCYQ0fKwS
am/APZRPAvkWfEqkf5JEixHi8jbO3eTA6FSeCqWXaK7rcVl7POO45UwdDjKM4C6Z+I/U3I9JxYVw
3mKghODyA+qUg5ix9VcrtYgMGXPbgWi7SnJTmOPc6bPBejuynDl5NoeKjCPz/q8UicAz+TbgN1kQ
IkFVp3SQRCUSoE/lfErUq7sHyLGwwajq3nHUdJ5HzRSiSYcJHu7s1xeJ0zTEs8UdhaKHLIMI5CUy
LuvMxhaw7HxA3I6jlA0veq9WEQHdGKys5Hr2gnIogvFs2AaBJrlJg+jOnQ/6rt7CHxLW4AhseCzD
84cmn48jD4hgPn39g1TUuyEgi+ppL+RiUiiSh47EzdWfeYVow1D5HSVKQZhl3yi+TJ2bXtwcCVkW
87nMCbs7s+dX0loRZBBc68w+ppS1Q385sCRy2uxXm1Sgc6NHkzHRd4PyMtUW4d2XeVHesFfy65xM
De1j8Ek814xJyGiGr7PSHx6riDAzIufExjvyHxcKf+bnhlsjCu7IP4NS0zOegQwibLHTHz7dOysf
F5bN03yvlV2msB/pQ/OnHOBriXCOddZYEdqCjYs9krTQE4Xp39SApXnyaR2DuvxC8HllUzWA3FOn
3cnZJ1MmaQgA9dNmw5Ns1I6gabtCVKVdwVg+t8RY4k8JB6cwMUwEPcBxoj5kQJlJ3DPITSN+6VSC
+1Ac+Rl8KXPHMPUjh5f0OnUZTyfgRDNEA+VtNG4AFbmlzbXam2VA0Au0EvAXWfNA8dD80LKhUkY+
R4M6B9YXjK8D4KMwgCQ6yFmuOQcoO9w0OZE5iCkTuVI1wOKufBJ8zks0UqyuTTO8f+2Y6F3oSDAo
K7DUHE14SDRNVcuI0MVjPXB+spUw243bmFwKKdTc79y3uJpoOKqIy0wVXPi3ltTPFhe7sdzD0lnI
MmNVROOrsGpmP+C7AfIyPLZ5ROv43Bru08kQk90tY+4MYyV9eSGwUPTSzK7uWuo9Iae2ulINTdoA
sNI0JMscZgADIzZRCi+S+hSiL69t4DeCe5Ql/t1+jIAQYUGBAyhPU09GhPvgnNntyEw2B3VGbI/s
B4rNaepNoo9U3SAQPUO/kd2rcrONXSPkscFkeYwZP8bVAexuovRuwMpnMNzGtYZQKrV2+K3Gdus8
wpPX5LiNTUK3zU+nmTJaD34XzC4GiB7U5vTX57B9mrgoMLs0QtZOClx0tf75vMj27xqG+ohhQjCb
NERqyGWH9x7D814blufUpHrsARAGqg5WTfpZAap5L47jbFHqN63IILEhGogfZKrJbHJfU2QXhhQX
OpUW4Xj0aZSQdXTBRSAqjjENK1f50WOX6Gb8k/5zsa4LN8KofMFJUeJbDLHE9kDKiYSJQrjm1I7S
9QR7ZCqK7lT7bAGG61ZQxsr26qNiuqykFGiqxOEpAIpOdFYL9YJMA2akw0CtViaMzqfndTkX7OQO
EV0Hxai6uXREEGXEnp6y0Bj4snDVVjAx5zI0ta0iwXTZaezBSrUBpWbMR9dSmDRXpEFpANndUEtj
QpRKGU9B7BbEoDYAlze7RupQoLv2wXPvuJl4Rw3pwgnFUepAj3pWWoyoFRMd3YSYJtteXo01aoYI
BmenSU1F3iJ9PmWcJ2fVSvYUyACOoph2j3xzHVanl9im9bTQeVIz9s+cnNxoJ+HctimawEwh7HDS
wiDhqKkxHsocGS3qr3OGRSXgDMk6VWKtkgWA3cIgJ1CuQyWAWEbQ1DfDvKKPENbJMuShWwuWJaEt
rKmLwak6HfijX76e4BgJjy5akK+CLsbpABwRfT9bnxrpuMmBVck0E/FmZ8mvHtUEAafthW8svwDG
dfVMD+TZAKQ7+/0LUD0wePlhuvtoii4eVPjtXPpXHWvVlLvAPTOVWkpdQ5mlMRljTmHjdz3D+WLh
LS+g2E9XMc/7wPPyXMaC+fI1UUSoA9TnLlC3Ltg/FwV+8TKtdi1jgUrNuSsULn5YXF58HDMYUhzW
FyNfnn49UTMXCPkIS7KNg6hGSgIPJ0eLmZeNSQKyfbIuApCIALmiz7wrHoPudkiSy8XQxjNlEi5d
qIb/IWahcj7SCJik9L5zJthyfwS74wj3DH3kam75ej+xBbXODTZ+QYXxGRBM7AWUojwAT+25O4XQ
hyMbEl8+DM/Emuga3JIog3DLcKf0MiBhwoXaPQuZPHeOQTVUqQ6Yb+k2F4KFCZTNl4CdxVX/s/lQ
txuBWeZ5Z8enanIJRCersTSEMqCm4t/f/g7GugiIeMOKq9fcYQzhZqG5dnWr6KWbWvtA7oen/RT+
c/D/jDyuhiwUzOdXduMsPXHXS1GBq6E4RNSw/rZ/uilgNgW7RqGntPFl2YRV05tiCBcN6Y0uh0pj
4ZUR7x+c4eFrmJ/VFRyYSDbx0Q/ag5m1Wy1FGs3nZn2a7RhSBKWooGO1bLV7HkhK8FkD6m6ZQ+hP
zTjPrHqI+AD+E5YKORovMUaZ6P1uUHalOw/+R2LCrYmvWVothpxlNA4c3H5uU98TlFudk+las5hC
0leO6GeIBhum3vmjgZlqlJmOJIAxvOSVaA7i+lucoQo8nRaAONbuitvy8OOwSPrUIUk87I0+VNKY
8EhtO3WWxdlwP4G1bhEsR4a7E2LFSMbyLroyyuwWPb9uz74n68vzelBEt0w1kUATKk0NCdYbdyTe
r8mH8a1QGE3uiahLCpGgbSHyuwDH6cYDbhMKlcHllQNflKqSCmGSqQv6DO0yZbZ+VxBjWFRl0ajp
H4qThUl6STGbP4trXtcXXIIU2VOeX+jH7zdu5e5N2Lp1kBw3DTKGwZJWvnlgmbTUkJeOg6MRud47
QBbhCX1PuHiWwTrDPkVlE0yYcfhRJ58GchD+TUHm/fn5n7hprGYaaFH4aU5J2r5rNQWVcjnjSscV
vNwWI9MJmOYQq1SBMNtcIZm0rdVTZk3xbBqwHiOi7TOTw2vKc6FmWxixPmdnup+GhG/xKWV/p+8g
1VsEktmzZiKXRbruXWR1U3jy/ceNnqVW02XuWIWddh9VRi/cDE8Zq2HrFFKYqotTomdFnHX8KfeF
L4qjvoMuxT7q4odBmFgSdCGkGZBicTCILeGzAMOSHz3Q6sBHTOjby/0ZCLqaIrCsf8XOUGdcvXJh
45NZPdfsEx+3eOPudMMY2Dp0DcVVcOkCL7r5CUoHMkEwYArei2O6buVQ4txLN4D+CsMIF/kMGIMg
c3BccrjX36d/zwcDIWCcBPRcMsvcDxnL4cJ/GCnL72DgEF2O7scwqNtwJPPAVlhst1iyOSObixz0
6Or5B23fXs0keeO9UZk4wRwtLpW3cvRIh1mfnP5nMdNFVpESfjKzjPKh+9USLACCT4mLJviUmMdw
JGpEVj5ETM49X8nRLHaKsmR+H5ZpyxpbetPvBkhDeoLcgGo9n8UzPffkuXf5T/rWMwEJZeXTtrXI
aKVwtPdsaK2d1LphFNgY+x8GNoP69pGrJohNy1nBdVEAuuQk5k03+czr1OHOHqh96dqv7gHONqnc
qM7XL4Wp8+Kzxk+QkVX1K3Xrhcn+0hZEf7Zo4g6IO1/IrFyXoPxDGizjcB14ZDNWLp14OgilxDD7
GlVXN532udPOKaiQo031qVzpX3OuJN+mDgpliMVO8GoXHgtamRlQTdlPpg+ZSqjYeL77RhiKEGXz
wsRAnflTbsGF970yvwHivQE1D0ZBj4n1c1uxmE+msVumNgmc8yhbOZVixWF4jpGck5vbU2nUJA5y
P4WH+nCEwHyEjI+S4hOGElj9f9g3XSEvq4hydJGGQ/p78OX8p0e1OpQn5R5MLiJk6yxlPVcILzMj
FEWgg8No9A+TLABFiDonbbDU/jOJk4fjslgl3+i4SgC8EMF/0DN4OYK1weBPpa7jUFpk7ChZbRHF
vuLtVE0j4S4ym+6YxegyIhUCGolhwe2OmfUmgqX1ZlX7dEXzWLpvRXN+SAE8Z9nv2pWPtBy1fkJy
DnhicAc6NTLi6IA3ga3pD5CoMsAbxtpeFgu3mehfGERBRqhOjB12cuxFTtnnUQSpIOEK1JHXGL8s
zB1OZUJ0k3qy2Lyrxnkau5kC4ZhyhjiUbkwg3FxEv1g//BpLHkW8pzZKZ6VSthUdLMU89UF7rZe0
IUaSyqLbui9oawGyArH9RlOrBsOcoBaMxh2fd2s7/LtMwjDyoxaP3OlmzIhxLgGXPPj9EQi74jYf
mYJIXOXi1rlVadGZK5FBgtGpAEL9OT60ihE+XQJtLYF3vXzGXa6+5H4+ZC/Q4QuIL7dKk7h3I70S
cLW44ilK4UIl+/JZBYtI5PaWnODCs7n0XLOj/9t65QrPMlbt4QfwlqeI/AqYicLHAQE68FV+L3/+
Osq3Spewj8xhnm0n1+6CAzwpiI0oUiRXrzLhLDiTWSv9jeYo/Dq6CkuxeDV5mGR91nitPxAyjIdM
k/TtDjLv8l7g0Chw7ZqnmHXitIivrdILyFqkodMZE3WXqMxUVr4eLz1Mu4Dw0Mevz/YhTqITcfen
z4FpyKFg/aT5+m9/20evbXia8ZDCZPr864o8vzRITgmnekZylS1YNWg15A00rszfGgqmIRA9JLRM
/ka6zNKdVRlTcXUG3k+iwclrI7rQGYlKCoC8sagyLOe8n1A+gmBkExSUPBf3QMZ/Ff4Qz+NvKfSU
OZcf3cvrgux3RH8K6MfYm27U1q56fmUXs4JPmzhq8gES20/2QWqNP/zwjilS74jNnJsvELdqn9Fh
NaNI25bnjP/UP+V47/suMf5UBB+p6/b6GuRBwZnSFvTVmbcs7tzoIo/HHDw7aQwaoEZeJQI3bkLO
ZPtovJqJ/z30paBiUET1vgcxEX542YJnbgksEHqjNKhTavdkEalNwW80sIMnoNjN6Xish/BrKbKJ
kXG++CTKN+8XliOVu3pQUnG9rBOSioN3NFr3xIihOmaxP5bkLhlnw+OcntcBollkNIR6sOhrfCFZ
C2BUXK5kfDz7qUZUdO/FL5ELvBsY3CEsJCqOLY38Cnjuo9JjiFJ1/ZSbLR3f9BCnWw0rZKlu/rJQ
sgpJyyreBC6Ybo97bKFr7LPmJ78CZ3BN8ZBb0EUiDNRVykEMwrpP5cfFx9yosV+CEpIDho9Z03SE
2DEX1zSN25MyaLCeVabrHyt4y/aeLDGqqHt6yYYCbpAPAyz76SlDO3f3IRVDLUaeO92Q8koYA5hX
GpmQB5d+oWsq6+kD5z8vO4xNk2uhDJs/4Iyw8m/qcRkfUGY0GT4MoKbyvB1DWX85Xp3ZXmlwWNxT
1fZqOkInw1lG2tomR2PtKsNbBLTcNn3mGFesvr6xym3SIrrX+346DXo5yPk153UKvgO3c2U5kGFz
iDksE85BiT8heXx61Ms6+8ny3BwhfkLISufkH6gTaY04/ZKlVCEzkW3pw7nvZwvLQtQqZStM3b9E
H3Q3G7PNFZ3V8kpy/v6Svq5gJnVq05wETN0i5mANiF8V2uz8zBco+/mn2HgpFM8Z7kYhNErQ2BKY
3ltgxr7/S9GkJcnvy1R58ffGUJYe/6oA0BiPi70OJXJDUA3etp2me5tdcqdYSVK28o++ugUDiCCS
hkaLZIgsKtBMrIxODhe9BxynHx/mkTak80om4LbdW/h0CbCbDF3MW4fBNbqMONajEv5Gl06UOTk7
wYabI9gAilA+6Eokq/tDRTYTisPFxbd7vd4JXQny+XEh4mft8GJ+IZb7XeHWFcmkoPkuMUtnLWrY
bnHyfMOUxfsBSfBdbk1o67lYvswpBpFAj599AAerZI0yCqpHcNLTGFGkxrxCojtJuGcnCca6h2mQ
FcaF4FMxiMxp+3AxncdqY0rzyQALSKM1t3+n2gJsezC9dUur3m1gSZiAS9zoCuAHWLcEJtvqA9Bn
1c8njgs6PeKd0DB73shJsdlw0htOdAp6g32Yu2yLnl+VkWFsF6b+RbxE/Vde/u/ZLpqvlD090euv
84P61uYUynBMBs4jj4IFEcYkS1RgdlTOSDZkPyPlpT3ktOtW0Px6ycVNY6HcebI7bGXFkXY9jWVb
Nry0cf2NP3ll3EZWMYt5UOblSLHzWZzcNkijMCJRMgpEMZ1J5YIzm0hCkkN3OPEnUlwWwA1+gxDO
KIlepjO8jbnIBaEhj97VrnmLAdG2gsxPSd1nyBOscRCpMhSKXiKJH9x+mMTDzgeffwDzJjg6lifj
b4K6ai8MU7dEKDqTRmSz+uMciKqk3z7FlQbGixvROZnw2pBNCCLnjDVSioHMMWT5BNvlPbqDXHRm
vpbd+uni91/sPDGXUQeXe6MwMPMpkgNmLzRIDcHS03fTw9evUrl7gcLlCEXZUnJWhVBWrC4gemjK
lp5eA8pUsvZ4aaXPSRfo2O2FhMUB0K/fNRfo0KtxRH0GvAOOQmI+g8CT23xHLQ4z8hGxFqBAvkHP
esILhW5VVSxE/JiLrcT4vXjcE1gSG0G61Mgbc6Ajhr872kqpOwL/T4vzQbecmJhc69HtSiDuux1+
JDKtsNNFQAZ11tOH09ADfcV4UEilSD2lYFaabxubVgioXKhKPhUmvt7JLtUlrgQW4OkK2EK/E7hm
AeUa6rJFnW6uZr1hvpR6U/r6UwwyF/B+KQrRlAgeW94WhRsLJrMOxTyZFvW0Z1N1jwl2ndcD0pWK
c/D2dwQfr3SRdC9ll34yJf1t1QlxIC6xu+ZZi9DTqdqMp6dls0COYTbj4MQGcxXvvpxs6xOQOWTT
ZxHZl0AS1I9FW2yvNaENm9mR/7MfUVH882aY/qeIy10aZ9zm47uXDin/JKBlT6Z1Y0UvWkocMmkw
LZDQaG6IA8rhh8saHDRvNib93xk624TK/zsPLuG1lihOgTir1AwzXoso8Jnpw35Ame3xWRSUSJz7
H4OoAjVrZzAtwM9gpjrxcFef0tD99IcIypTBdehqH9J2nXnwu6Koz+Jr/VNqHiizMs5zvNV++Nyi
z2e8hkjUChK7XAypSdUhayJMRGhskmnLvA+FbaC3dXA9o3NJ9Y3DEFMPkXS7dyoT2sXny0T0E+yQ
gPd91y/Of9LPiRx0xEaYayeCLra1asLFTjbJnqG9KXu4YE0l1h4eznnlWcnHmssrX+NSmAnMml6P
6bkbK74x2wsT8oxBPmffpg06/XoHYyv/Ft5lmMNUrXQHQd2bAfsG88PXjp7z7dgWQrzHC/N1xymO
IgThAmCFwVckjQsYQuBL93am2FvjXA3OpK/oOSFM9S3IVyx+ZtKl3PBm71DCRZO11hXyTG94mFWT
UKdGrXzUnzLK74/xErfYS54EkHz/8AFVlhqxnCYC082TKWUfeFg6jilbr4zu8O1FJRh02kjYMQkc
2mpWYd/rRqOz3NM5eP1/ODQGZ7qu/xHLqaYJv9+1aoJ6jAD0CwsC2/Iw66uCyxjNtqdbvgRpC3tT
5m57oAWtOuGAPoAG77LGhqEgZh4V4GIbVe07f9DJ076DsNvmCdAvqaMazxC1Ff+wQpBGrfb7X+UN
u0pkVqK4pYXoA28G8EDYbKxzmi/8fSqWLL8mcj4pPOfacaFWrPeCsSjHgInlB9T2JyWyq353qb+R
asfhjnbJmaGAa2wfvE7WDzA5Z98epZ8yyE04GWlI5n6gOOjlCQp1Cv3LxI/3gw/JQmU1vKfdxbnj
8otFH6H+kx2/UB1FtK3qewMRajXlwMNfwjVfqQ3Gef3reXE5aYzLzZP6nMOrsFGc3joyWcRF3ngM
qd3whuTIDjE4XW8ZQoDthtKHdMTeB8JOCry87FBq4L0zpxcwzSIAPeJQCApEHpjLVxB6jNhMJT0Y
dQQ3dw//xGCddbP/uY/0qs8vY8r61GnTPoMcpg2P0VJjRRKhvMIhGYYc1Bo6LCd6KLYkrOMBK3Ex
q0vz2BYO7wlDULnwYFL+qGmOsZIImURkqi7AiqPxKW4PJ/9tLCSgCqNC2rsxWVUBVEAfm/PdQP8q
GAaN9OrZ86nl8Cbkh8RtlHU0CmNQ1mzHodsKlywzrIpLHqooUebs5K5WwOoueC2geXlSUOF/Z/U9
kiCzQOIausND2pKCPlBPbYymPFyy1ak7tYUaIbVQTrIsKyEK+IqWXlqz6pJ5DvuyYoLT27a7imrV
yGbLJmRp5ys4fk5OJe00SRKPSl5DQ0qoMCO8v3LjVneU6fez7Me/m9eU8Lb92nPSIYe8Spk/zRF7
FwVXkbKMqb3YaSDE3+bilvpgKlhdsSIkze7yf9X/liNIyuM8M/vcTpHSH9AQGwqiNo8Q85WLZ7A6
rnaPqoTmCS4K8sgTrPdQ3sfepbqIRdzz3JDJn7I0ZcGYVF5bjaFebHzspZtsjja7ES4kpOc7n8zf
BtRQf8wTmTWaFSbAvSFcBeUINYxWeptYnLihEE6JL23cTR5Yg1sBbP8LOe/aKTeAqQ4bBDkk7uSF
EHJTgRy3Uk78PlWt+KSDFWxAmjap87kqwl7zX9opUVy7zoKj0E27MzBVvWsQQREhQQw49dNLXIHC
uyiwc252i1l61o8U6VXaSP2YolRbm5nURziDfM9XAmWVk4SlvZ9HbkzkJSe58U2Zt3DRLGeeUUV8
/nO/INKRrbzWO/QOAxc814D3h8u/Bu45zeLO/6S2nd78CUtCYP3agtrdYCsKv7ha4i6dlVKWPNs8
fatU7e6t5W5K2rId1P3ZxnE38p96aTHF6A3Nt5AwYtq5gjo4WWJiLXC1TVVAJr1/IK4h7NNc1CD/
ED82O6ddL8tCgmOXPRIrrCDS90hvT6ziM4EtTCDnHvCvOE7XDxJEVORZUflLMSThhOiGQzF+y8ny
y9YJdKKtCL0fKFMsohCIu89k5lJLzMNdIJp6P35TPby59vH48Gdf3pn/69VQ3ye6bTx7tM6y24j6
7+zI71+VtzJgmAtQ8K8n2noPYLbzywbWBxk5YIosvt6j2x915/eDVT94DA+u6MgazHWY7z00r7+W
pI57CJwQtFCdZrD44Dpd47+tyV/bOzBw1/AkgvG/4UaR0ynDMyj6XMVnbxXjlxV7OdAxhUzUjtii
2R+bEjLe/SZVqilBw4/n5G44aMvBf5luyVtgDQKDE8ncL1xRZUnQDh9vZen/0fNvk3z8PA7/mx02
hz4LCBmLUOhOJHRxhdFiuEtPqkuiZhx8Zgu3+TCxl6hOH2lVAji8dFi2HXG/9vuGHXQsi3mRNy0a
27OQpuJ1FlUdUQ6Gg+UQJ9b+0UP+iwhu2WlYOfXSPnUA5sDeChL0raVBQbuUoqOatHmlYhA2B5N9
jGIBXLhPH6FLGpKWeVaUnZkYOBLrmjTWgVn9VqL2i2cRI5DRhumryBmCrd1oj0gVwNFIh7FO41ay
MKF8Q4tSoA2VenGjQRAswxT+OrswTR4NcmOEp9apjdTPIzYgSVj9yujsZZcs8gQ3OiQOFPPfZXlI
v2Ccq2tLYaQY2jLUxmA2Qr6A8f59ZziXBDX5fFwPvWWFy82IrOEpwRhv+nT/mcTGvhRKTT9eL60S
qI1WQc36i3uOzu2icUb9x4tjGMHgUl6xx/5tvfmjwLIfEVW+C10hn1HN+H6JW+gDssCOn7IdKtuL
Tnif59e1rF5xsoBem1L5TnnSrItQ6+SFYad5aAIA38Amm+JdLwmUpNi5jPnNX3rzDvvQoWzcFeH1
HICfjDuPOqPNhbtqREFOm/N5UO60qehFmZAxp4aw333M2iftGUo/OLAqGRqu9tiIyWlsuQJ9BvzL
a5cy54ZGwSC1VT1fowi1GWIPwZSxkWK+WB6SE7Rt4inexc70b3Ir0qWn3qcPBpkJ1KpinZsniIDJ
Fpjj0g/xfk+aoLvKvMqefY2kPARJAdUILLIVztDAs7WtWV9MLgZ9ztgaB5G5DagPbgkk5k9m30MM
Z4A5+wOi/PHh21BIWRl2VMCWLjzifoHaVMT3jSf4mK5I1l2FuOUYNgsHAbq/1XwWaz/yS+KBcqx5
uGWTrQzKHg1oQWyhyG0Th8jNXlqYqy/jY7gAQKV+UbPKcPSwtYoWcXSbUoElA6MF+wOpUPfHRTgL
eXV0cyTntLZ9UVqlkWPi9Xcz8YXSs9KHchKs3ipRkLbyBMteFX83Rd+rrC1kOzsbLEYvAOqIYLqU
BYaIQnTLF12DX+kdqvjp7nnjLtb5iJWWF68yflIx5jEHFYzU37Ud+O+CahEsANp6hhdzMn0LOgAx
OrylNKBoHduXbPKGcxGfqLciurVTmlG/ietYmHi6rH7y8MFYeL4SUtBI9bnLM1u4vJ1l8ZPsQq5m
SEABEAzR/GGY4KsI4y4eok7JhZgo/xaGV2u5ofQx4JzhVEDwWt9ji3vUnDGf0vIZQI2BIM0yUYL7
pqpe7Gm48kpNuM9ayehKFOuEtx9IHDkFol2U3d0OzVBovJDZVO032ysmcNiqIw2zFF1bu0IqrFUt
fzbTFHFwqfCHvi4MJPR+/WKAQvzYU5uHr4/9E8YVGTKOTmuPvtnPmRuOkNsPHUGa/FvCGqb7pnF1
2WXC8a2QHqfwGL85akw1rq1NbAXc64ME1QvaIvsrcjiSdq1fUxGaaBHcYBWUggonu/IQSouBHPiA
CkIePNFUZ98hCDMvelYgCnF5HNH5Soer8PSVJ5ZGb5V9Ozu0zgai50XwW+JFYCQ3xu6xB/sm8MZr
A6bx8RL2LFJrVofleJR4egWXwmqPjTSdYWNlQ/R6eUA/S2mNUaRBumXIgwXhcSAhINXRo5f7HAl9
oyscNaJ56rtR+OrSrMPoTrZMtxbsVH3RWc8cjvaxHlK5DgVZbowPXs8aXOxQP0qO0lX/79J9fiCV
/5Lz50VYO+HGPcDDbytbppWpuPgXvg+clBRKIDyYbBC9pcvtvoqxDwGvsfDJWT2ZZe3Pe/UsGBgV
uawXJ2aShJfNvIh6/sYzR4KJmGK3kwvNhvSMJvstqYZOjwewRLuKnywl0nRqfAN+FTZhBnYocuiO
+8o0NqWc3yLIG3bEIcagZe4llkX/0qZ7VtXdyI6gWBsoo6ehhanoU1za7bYEHoFXFvmYqLMnYVQX
DId6z0fCWVKUud0+Cl4f6EFM38pMNOojYwWqax2SdySVgr20wrZ6X75q4gGHV+MuQnxIHKDQjcKO
V9gBxAMi4hLIXUxZcjJjb2StW2h2/NvWGV2cptKDpFgxUzkTio7vl3P3tAiYxtu0AoFXkHEX0iRA
Ca0dNV3WwW8suxuX5u0v73poKtxt3zxRJ1oEXOMg1jVsy4rblmnI1ps8J7AUQ9YGs5bSg4sbQTgg
JdPL+84Nr1orb3niwQjT/lCpSK29gMhTHT1+PFYC+nnjbzH8j9KUiJQBhMEbZNQ6rToh6+ovnWFK
ja3BBUogp+G3zljjzUQLYjt50+OBfxvFQzSTtRHlcBDF1b98ZtQh1lX/SHQ3VvSLEF22hPKCl04d
2XkB6YfqFQF8ZwabMdEQfRrk4mzjR0/eIERES+jFPbAG5ZaXPLzmfsn1B0cvP0E3JqsT99g8FRb2
FBz1/jDL5vrakZTKEKqNFltO18X3cGZaEhCuVA5DwaUEsrjp7Y9HfDt3uitu4EM4efu8+irQbsj2
cxdIU51xnbD7qxNJKkc5ruROixd+erol9ydeCS+mQoYsrJX0l0ygQ9Em6rGOz6FcoNlbCAIJ6ilw
jRIQZ7wUnimDH1w944k0Uninc6Zq0S9+K+yLAq9AtTYAOVFl2TA8YJEX8hrbquQEPZz4ssX1na6j
BJRrJcJbpe3C69ky5xLgtSh5ZFMM8EHYZM8h9sjaIejjU9Ui3IS7AUegoPMXa5h+Z2hb+Rshqvmd
6whwTQdAR1ZfkKLusE7A+WJp4vVicE3ctzLp+LXgNo+nPU1JCcvex9WBbk+qZkAWxhHcOJcH6sgP
c5WiyBjFTqB5EUqk6orFWhWoe3hTIoEr5g27llXBL6GrYA/VVE6A3/YLuA/Kfx0h4Yxt4e5X+xDq
thp3K5wbLwJVStnnxtfMz3bKmC93Pg2p8yxM75vgIxlhJA7CxugMctQeWfy6FWkG/CPH6u4xMgjX
mMaLmR2SmyRQPLjBZxADflJVG/PeGJgkTnjpXMhd6oQX/VvqKcqYMKhsnBj3c0WlvciPXiy8plJ9
zu1h6/713VNI93jX8BDvArbxgRhN9iPk/CwgxSrU6DxbkuAHPkoYR4GkSVLQOLb384R1K6Bp8fst
vHcMT65XUZuuV1QlX3Y2D38YTG8g56aC1lQgVoqbwoUOszq1NkEJ26K0xFiuRL+GIi8bmv5OEwEI
vtu//niamlyeBF/irNLMRo8yPvALyvAbm6QyNup65ntDnsApQCHQUAxZI1GbZe3YhGS+nBJliZHC
nwsia+kHOgLmiJABuTVR9o687s+u4vRASO+GtQMljF05jLwdjr+jF/AGZr3+pR8EIxbtzEFjz4LE
/0lAaxhgcppBd7SbfJ6sdaiZ/OSiZ43sBBmxIvE4todEgUedXoDGGus8qrif6KTSZeGRRuyEbamg
5Rzxf4C6IZ/OaVJry/R+kLG6ODEyHyigo296riC4Y2lZbiucdb6adq3f/JFmk/HQN0ZuxZDFvV+q
oru2QeK/1VdwDWYlo/ut6Q88ce21LUZgkjtlQ+Hf/4DCinkFQdxvMs9EvLYQtRIczJ/S9fLn8rZD
0wL+APji5MzEUS/eOMeSbb0bjWvVzbndf6R3bQJwRm8TTGz0Iieyo5HwOJ4jd1oqVuhvpQCXfo47
fnKl9s+vx+p00m2SGlvp5qtxvb8LJ20ZtrH9eBx8AyEDWRyASbgl4IT174ffqoAqenejL027HL4M
us3PXk/IbnB9RQCE5qzl6rwbzTu9b08XWsSol2b34Dy8Hwl16VuPo9aA6uDxeF31AgKO00bxyTm0
zatVFNO5ejdgiyMgm48gkOy+T4mVnii9/Wthc41AsaCv0Qo1TBikY+Qg6SMCUVZX1gCUhrlY/gHa
++iK4/R/O5Xgt8P+GIFTf7vf7uATSZOlED4E22oTd6NpWs2yD71vYkhtBEx6TVl3WNAcG0qMrwVw
AXQgDHz6Sc5ZtrzTQnuatm89o4DTsykB3wscT7BgilYzhY38WR9NA5iHXIM9JjGpiHpq+7eqabsF
WStzG9ejFBuJCVZsjPt5vnx3b9EK8GA4+wBYX9GILjoskxFSvyWG04F039JduVHbyFLXqwQyCsGC
p9gdQzFqpPva6UXdjMfgC8YQ+9qDGWjSuYQJ/lVvKLSm+RwFCTz8P1fyETYmjy9Qsm6ydYDLtyGD
THV6C418JnekIAzAMgmDpJh3KHnBSD6qT77VPK8LSwsO18RcTAthH3CcaB9OI/iN77SUbpMUDI/S
k3MZNjE8MYINT3lK1GXm4fQNtfw5SEUloAxdrFEN8LNrp+CO15v2nEUPxbJJKMF68M6epOSE/nPr
qzm4Ry24MqJ1PiZVdPCfU2QC/AM0WoRzSrirIWSlA4x2QBfnbgWwVXB+YGzNY11kLIgw5mV6BV8Y
viGBtwk9RWQgbVCO/WTUuLljlwO0XMd0XiLuFlDoxsybAPUKdBGYTWNv5zwHk8dlU1UUmEdSRKyQ
NXhvfacSIIoPhq1q+V0tlazJQD3MQeT4s+mQEtpqPB9iios0jgxgydF44he0XEcnG2qSLxYcv/D9
+tMvBvGxx7aqGtaaNtziZKhnlNmK7wQNJFcjqSbEXOGM3BWCqYo4NS9lSVCy4MICKfebCgeMXDFi
0axEi+aTDYPiY7LJyDkFNEjRk0zf4ZYmCRhqKCrUiRc97TH09NkPcLyUPBZWk57XM2FKa87+/Ado
bC6levxIynIJscZUK+aqk2XE/DVXXFspk7v6vK5/Ii0B5QTk+4fgYUIzfrlnid62wGXr65seewYL
6DJD57P1zG9Hi9+RO/0STp4/IfZh+sw1fu1/2wcYL3ynjjH9s5oJ++irk+8XroU5I4gv+RTaC0m8
qyLx7Ho1Ha4ESZhILbsthxW3EM17fnVXmPmD+hqo+H8VDkASMJutLUU1EQZNc4EiAtyaQpn2n6Fg
IfbFCuRKIAUSB05EKDh/WkPWnr2YmzamdTPoYNJKfT+Y1+wRQxuBdtDuMMMO4iy6h71BhZRyav08
93vgH9RNgq5Glhpbne0hlHzr/Yp1Cz5YJCrXAUHKUW4bGpFAxHrjr8jWtkxZGJDEP+BER1xuSQ7g
CUbouIO9YFXSg2OWB6vRxrd7R8Zh1LDhaPGtcI+2n5T70vnONK2JNp8Az070hIPhKe1DFbXGddIL
UsZB5VubivrgomVX1oZIGwsejxH+jYT/LueJy5s7Z0cDvenO6lCr0ZyJvCcfbEZYTmPdYFO/F6Hh
5zzexIogI56Xk8+rqUSGV0Vuw1GSllf0NQjXxCnN6Sq7HjEAaS+BI8hfIOInUG+Nq4ZmUkia8WFE
cTOHFC2NfosO2+vsdyxsmtTZSCMmZmeKUndC31c/ttbfVd00dEkyvTrv6ZH0buSKmiqiJIKLdm+d
jEUVdLm+ohO0RM9laogfbGzCvOHOBIxfJ1NYYj2uRGmL/FVEmJtWZVDQlT0nczibLJCEhIpD+umc
nNNzg9unOTh5r9GQM+MOKvYwr/RXZJ35ROdE9d/nsF21YJzrtDI7PCXzzRDCRjliZO4zFKEEIF6+
o0yCkcldjur/5q4zkgaN36Pxsbl3Z910rMs4crf2GBj6bSRjk8uYVV2SsH0G5FQ2zE+TkRPKIGuq
Q/nKry7QqgUPRCubydzMm3VE0G95bGtgBqxjViw4grx3wfXcZOsTCAG9dbcC8Q2QIu7ssXg6hTdH
XvVoo/pxANG0K6MMIDyQHwF2EjI3Aqg4ZAV+bOq1J3jdlg+ArO5UCB8RjKwcROI+bMm+7JPQA/J3
BMWBbpndGxBWj6xHJVDT4fPfJRmzjuDnOsTnGNzjt5jEvXIMcMZuvOmzJ9CwxqT0uKSapYKxPy6Z
fA6J6Ef+tDG0rx6w8/wpo9tzsrspaGfJ5SGmd+xr8SILyONb1lxtmTIyY37MTgDpjJA6ID2nx2Ic
0hx6HYbCZMA5e9X/soek60zg7SyMQETpf2osV42L+cH/oAVvFx8JfSE1QxrhXha8BhUGHOGu163Z
8fv1lcBw9WGJ12VN2a+DzjE1Mm6VboHV9EqHsA/7k9MR0U3+R/sXurgmEc/ymPh9NDnlNRWyDEZS
vD6/GJSeJr2F1H3p4II8Un0ajaUfaprrV3RLYO7l9GVtWM//1g5BuFg6xzCJGZo8vxh+QRaWTmx1
UYOlOP32gVxupuXEAh/rjkgQe5XBWXRtuhDvla8SWEC4PgNttJ+M7a10AlvCYJLQ0QDHYe1GXHFU
709Cc3kt6qbXrtz2hz1fp+wsMHo+0HUKOd2eBICCAvj8MD/jqHlq0fijNg2kOOduPb9FWOxEwi8b
kPoEWMLFsUAmF4Y7KyJQIMqM7BKzrjWtlKINiJzBOKcWMx6bU4MAr+4BiFg+RIeH9joOZU1PZaUu
4NF2vNLZj79o8gwSpkZHX830ab3pipgN85hsBLKDAsI9Tc1F75I9WLElELMRZ04GtXMrNVH64/Fa
VXP6z7cN3i1JMLAwsSH4GY/ca/WPO2XFnrPAx9Hf2eLsA6fDdYAYT+6xBJvZ0om4zZbnWzTFGsP4
Qhd0ToYsVCPxuhKI2l0NOwQyyG63mAEde1H550MwGH+ADQTyMLPHhhrPp8IFt2SLwmpzflVVVcOo
YAUGTfU7E62kf48HdiVSLUBjS/JgPUiU9bjd0PmLRYOkZJzAavX3Dw83nGHgMtQaA3k0AF+XC1BN
RSyzNi2LoPY2h/DVZ3k/3XgJXschVprx890QGC4BMxxUy6+czMCtTp8E9Lrf3E7vXffp4++5Dbxt
05tDKIUHrDoLfshY4wf9w821seKHrtceCzAJHtM40cp/xZW53V8u/zeACIwYAReYp7qDphWJweW7
yBYvpA4Bbu7AtyrfUCbG/AQ/e1yNZnDQHhaCIadrN3rZlirKGtooIjDCJ7VrFi/bedV36DXPDdQp
PuaMuMo0gDH1a5mc74+HZ5IJPhLgYvxsZQyPYUAdgmcmjD6UEllsezuTFuy9tSegumDF/nIAzvp8
B0lriStNgxZJNC7sY+ml6v2y+s7M1V0+8H710BRDzZhQl+LoJywO60LZjNEXRZF9kHXZknYgHe7m
8p3FxqbxpJplzUigRDiTWCZ4M1nYJve5psYNRdCaqop/ZIjPz6+sg4P1NVrkJ+XJpLz9ypaMZiE6
kmDV6W2el8VWvTqFKPdOZyndcdrDdOnfXtK0u7d+jbK+mDWmIJ+Uqj+LQ7JgxjSzbRGHiocESXT9
v9vSMDOO16/AN0T1hxjqdx5UWy9mBCJk7HVTXQoy9av4gGKiemVmTO0em66fFblKMRckW4QLAdc6
gaXGfpXGvwR6JN3sVB+KIdaiUh2jXAXT0pe6FGIYGsj5HbUU8Nv8ud2jDtgDdoHSeUdOT/0jwIHO
+1GuP45WG3/bjAugAY/K1LQcZelu8ilvZQUvhj+u9M//cNDoLSr7Xu7LxPphV8WNjojBuZSbd0ak
kiuGiaCEptP4riRF+elkzTsjY9oPgaS7drj+QxVOv9yXC8BpTi/lwwimBuIPMxgXSJ2NMRiqo61A
jRHkdsyjm4qgRCZcKHmzVkz/KlJtk0e9x1thxfRHQiwD5iIiEKMgs9OFCmKyoCwaZqUR8yEb8gcT
ZjRZj1wUDfaujpQ8SrRLXzUrp3polteI9f30dPdZtWbwxOzEvbmVnNKrGbjulu56xaNxup1tK/Hi
T3uTY24f0J9ozd7GiDnF6Ck5yFHkasxED464jgC/ONm6CApqxXxeoFUEmD3GBbex5k/Lks0wcTFd
bt0PBtNnZilRDPFJpsLvtfIinVW9bYuxNPViSBEpHG80KVKBoJa4DMHIQYYWdtQNpf/VI/Zamd0T
n3k/lOv+vmdOGiBwCVWwlga1vqjSr9+Grle6NqfKOhvqlDHlPvK3o0bw2tF0LLWE6YhCeU2pfAvs
RtEVmmxS15vO7sD6bzi8HNRFbORUx86KCB8hgj5pBp5iJGQCAo6ozMLmpJkNVL6iFYnvYBdJV1+/
MTANeQ8ihadpeLBBlwWvuqdkNCSQAZ1fHdX3tbDoqUMOOgsFp8stxp+ufLWAx6PKSK4NtzBKH5jm
D64aGXmWj7Da2pis7JpfFjpmfnkQaWjI2ykZSSM7jy/ycFDe4Ykjmp1gkNgoJSuv3jNUSm0TzKVR
DBkBMTb9uviz3Ier5ETg8WrOSGYLI2kcuPdPL8/7ui3s1iXGp1iMePjqxxpwmOA0SD0HoMuw10hH
y8atq+H9minkTaSky3H6k9XHUaCy7sld2LdyC5kjoAPGKbhqHMTNQbCv6wRTpvQoY18B68ncdleG
E7yxo06VjxySFtr152OlP2B0MDuQB8tijA/p3QR/c0UlMEvvnu69/aQrjjEHc0kTfSrsOkiTy9vO
0UHV7C1IsxyDzhZxvc95lRoUE68TArnG1pAMysOEbTA2w0SlULeNXRkAmzo5IShOn7rOKXqSbeTp
X0X5UT59yi5np3L7TT/8m6G+HL0ANKniTAIuO0RuGLzZRY4NCHfYSgfHccq8iAMrKIm+ZMdYAI5+
q75+5a28WsaaZaikdyNvBzLMI/IeUl/j3Kand2bojprA2I7f2YMmglxWqwH+Cw3YGxIz/QJwGmSP
8886nhhFDonVOTyqjX6ReG8zE8JP2OHj8E3BO5C4bzRm/yhrto5ot5e+YB/+iQEksqpfedM5ZZ+W
59WObe1qHDopaucqaAaRr23vPFO1x48FLs9ThgyiAigDcdjyzWJo2kDFzcmZ2H2ZUTFIwNkDcUdv
UIrIAWJ93A0piQ8fNy9IGFmnANxQMvJcoZ5N7ZPtOpAaoaQ2qBST0jHNvD2D+V5OVs+RaHFjlz7O
/dPepU8nCfBD1FpwtWIsRglJjj8pbAEcvD/jNwSTqCB3EoQhP+6XQo1llQKYBW+g4is8luj3SY9H
t0PNuZYR69XRq6qLoQSTfngw1uS25Qc4AVNfcKW2E4LV7bm7h9mX9I2Gbk2nLFNoL8QuK9CMfHjq
BxvHeOp4JY+CBVYBB7n+ZN+ievZfjvdRkhRdmkbHQXg2UmRtvxLuxIFt85Lwa1kLiBkvXt7dPWyR
J4DfUcf2zBaV/7s6YjtaztdQTkFwtK7rb+JQ6uPGFHjIAWXEOboKD5q59rLNzg2Sodtg8+lxl29G
KXyCVw+rS7kOaiSzqTO3lDtxecbrzum/gVTSVOslN6zAK+FVCTxuW1vUTgCkzcI15D/eoRL42jJv
o+5yNNWKTbvK0RXj1fAxGWV1AZCsePwA5g7/0Kta3ZFDwYABzYl517iH9PPS67EbhbOYbrNu7va+
QzukCIikX7jPXh1XBU7BobhKCypojZ3oHljqyXC3c3Ky7M70R4UFWuUnn04cGim+ZT48fJZHuTEo
R8zrLTUq8o+wYVsAgpSsZSte3S1pjg22oCx0cH9a27+n2qZ3xkRjXWngOIq+QzhLVbaRCR8rJtVK
VI5FU2KVR7bCrmDG0R9MPijOowUIwdd+KOGQIymA4EHK0AnIuWJ11SpOACWn1G0zPuVRTG/lVwN0
ZWqYIBn7tS3BaM12RtTaMaSfUjWxR+YH8xhm0P1PSpHUzs0IfHH+zQtQQD3l1QRnx7gzl289Wskq
vtqFT2GNKRjUvsXR0kSYX6vcLY+p2KEWZujdwbKlS/EOJWFSxRRva5V7PtJt45Qb69pdxIvbNZco
U/Fk+ft4SVR4lJR7d0txWhVQKkr/+sz4oi4lJZygmnSPSfA6Ju3dtSYF+cGg9nXABZ/XCiGs89kF
4mcJF7lKp906nqhJ4yps+TuuNgdM5D3rN089FfodeI4ccDA/05BF1lXWAnkUkjnHzUI6gZitY+b5
RCTvOGVFodNFlvKKVhPO+TWvK+j60FMQI0l+J62EQKjlxq79bwicAE2/cqrS6i14f3xXL5kp6STr
w3M6MwfLfyhiuInN/ac7i4Xj44AR4F7hnSTJ5i1veihqcGOF0gA0luKsjyyveYbwKc+jiMxwTGdl
y3+WVPQujOY7zmaCEMTYFouYBw6sntV/qbrCdny2Lg3RHDOBW9AB0vbLPhmCDMnC5Knun7mvN5nX
FNBRnwRQN+n68ljgGBmnajE8b0dDXnJcfJZQZ/TTYpMzvk+TVAjRPZsvLlNnxGcd3dZaObgltAnh
+h2Bqquik/kIGpSVKIj5a7FVy+gmPL9PS8KNW0VZNlpsYhy06J3xqPGkLpD4ndu5//O90JHH89Xl
2mSs9CRhR3h+LpIdukm2Rmks3UrtmNXHikIrAPp3XD1/QQ6SiO3MHKyrXHMPoFs0MpA1iLGoykf6
MrvFTOGuITyUtliCvm1qHcs/1um2+9DfroIxyrrP/b5DuKfrvnCwM0ZU3Tsmj7sccc8ybjwO3b30
BIN6b3n/NqNRN/+zgBOY71MQUtwS6hXyM9J4kaL4ELBdHdEiwnzrdcRQZP/vSj7VHHYOj86aeII2
LLLHWsRNfsxo81NNXkDj3Alg/kPBGtr7P2A0uTmPm47VwBqtSjnlvmteCLO1SmER1ai//9TsPUOw
Ob4lsoaEWOOIz+VDEF3u8WwANMwrgy1OP4B87kUaSq3Ie7h3MZs5187MLRv7N8KPYgCFdDis7LB0
LwlW35ea/Xz33aL/juRyZeI6sL0oNHMGkWV0FOckfwyL1dbk9CDqhC2H6DIZRav/bSWwX63fZ0Q/
ky6SwZYJiI5MRLfc/L9hRfGkCUpdYMTE47VQY6Iv3Ehv7rguEC8k6sFm14zhh32oOQR8ttTiyCA4
V9HsQgy0z78eox5kO/Hp8COBMRy2OWVvsgApyhyODCc9YGWEDsqlus2Yxf87aPppGh6ByF00AupJ
pSAM7Q6/ns0RjRAuGOxj1D+k73+jriVq0qQald7wiCI3xmEgqIvMLW/hwhjK6ge0HZBgan/ManIl
NC3kdSd12WV9oLzVR7Syy5pUH02Ms441vJ2fahUXWX3uhQwMor6SevCRYlwDIs7/6rmnFM+LtrsP
sy+wGiWkruGtKdMOU4DLte4woc6tqKABkFCo8rVDIw5AzwDwK/D7VKSumdm4RmCzVcqtHwYb8C9R
CjRmFBhCLTVwx+nWf/9qoxVPbUWd6iBfZ0pU8z/L8yn0TsWn/Tq39JLe5sEripy+QS9v3W4ZghgL
T2n1tUIeCX+0OD5EWnZydHjsZgtT1VYL5lmiyucxUiXliM1E/zZ8IX9aPAHEtZACigRZxI0LVGPG
MpxMpPg00MQ5bq8h0BZfCNrpWD3j9Lm79NgsrOq6ksoe67Z1MI6m9S46+R5Vj+mOXeQcn41Goget
d+usTRbjUj5bez/quwaHGWewD6uqdZQBpYV4M8UPEVpyv+yl5TCfI9PO9eyL8UH5FkSALj2cHKXq
PxT5DZofTCntYOBVwjhVgOcgArIWBla0lQMnovj+MnBDhzzTCcnz1shqzOfnPcWWmhhcsZIp+zE0
f7TBc8qI3EjunA0U0yT4vQjfFIP2UF3OG+lIcrsUDYwFVdDC6tO8WeJiYhyrA0VUkIBXT/kD+rYt
TNYSq2wHLMJkEZXpb0Nx3fmO3iLSWV2aEN59gqmb6NnpfCq/SATZ83ibLDVDQpRkTi8Ex9RR17Hj
oiSVtg8krD3Ac/sy5MhOkBci1O2PKrYn4ZUVNDeplPF0pPyWmRsMl7+L3+2dadrrHiLDLJs1utcL
M3bxHtTyDIHiULRkOkTHoatyYyjtjuT/z+Y38gQo6AT2yljwL3UMSOG1YtXdVj3z22RqyOW0idqs
dskZXHqJ6yjoT7RqTvZQInKzpxjk3VGB4F3O1nOfZ1/MKI7UkcPRdMbXIrERw2fxd+DdkyGXnhTr
9uYztL6JCRCkNOZprcjBpne8/HDBRsqFRq4oPsngbYzsJD6ByfrCs6oLYsFdKKsxkU/T89ZaQoa5
axGfXnN37JSYrQwPqDcdXbxuSjRWJW+lG2dafLr6jk2JzPT+6Qe1u9BY4i9Vd8TwuEwReXFsBrgG
caRsLNR8TbC1rAKAaUbaUiuNlCpejZCs/nK88fASoM3kDQ7y1lxMCHEeYzZVWVxGVo2jSIgH0xx+
wWmSE0SshkKLCQkcmMx7Smc2euFvrlvLtnCLkv3j7ZOQB8dPE2I+/qAcbBsq2yN/TLsV55Iq1mvn
UyOzJXeyOqj6UsLzKMJGZQXto/C/GMNFIxampbFh1nFNcxS1hriksdn1fSQ1NvdDgyaDjBmA7/48
MtgIrKl2/2aPywoyUdJnl9qgJU2guKTlRU2SMfTrc/P6MCPMp4PXrTvh0V5tSUAR3zwrNW/HF6NT
9+LwBBOYH5OKzqglylzIg0Q50Y8WfPM9GnCzviHX1fxdXpoOzHuAQcIiSV1BhUx0a2CfE1t7oe0O
JhOJqOU2Zsf68DFkrFOdn26Hu3IHzS66Z8SGg52Jhaa0yfQssHPgfa4U0XaB2TjM0VEHduhs2j9L
o8E+tkCBpYs2tjEMgx1MYBzAvt1cmn0StnvKTi4UxktH9CDWJp0MfHCdjTP5PU+6Ec6/xw98asOj
5iEAsHT/uDASSx9/zB8HjstFKnZDm/0XfRq0kGEfCk9/cRQ5SA24swrY92KRrGlhT0/MwRF8aYOW
7A92J3FLuUW0FR0JO0XEnt+8h9VXKUGMXHht0pZWlSZnX6gqfmE6MybYgmvEvX8CHm0xbJ2zxEqs
jz8HkSWW2gQmtQRiUjd/uj3Tklq3BH0jBV3A3Qz91cebqpMC6CDx7e3SiSJIRiBCTZ4cagv8SjyZ
ltVRABAGQiqy89KLj9koEp4Bzu6+fK+7FeNQnv+BLrCsd3hmN6iRJMnvnycCN/D3tcL/HuajTRTN
rH+ts7rweMMiKfLk5TDq8pZ0jBwy529Ssld0ZwNAHuMoCNiaZ/0V1GI0rIeczMYYeUj+xfapLZr9
YPwFSv58aXN/FrLsQ4SEG/UULx8dDVM0vGT+n6MQrm/qUxi0JRwdkibwD2Nc656bEkNbMiTMvC73
Fj+AVm/Cfz19twa6lUMkVA1X/rcWmX4enuyHmJoPc2aSMYg33438Bb4Xe7jfUcQ+W/8V6LcPJSRG
UpCsocM0Jc9JezNTsacwJ2W9WVIcS48oQxBlTVaJ8lhFCKgzZByJlS7U7bXRJOJfNCQ0ZxAkk51s
0ffLSOK85QJ30qFMmdlijYeC6gLzLGKDfxF9+t55wTh1C6ISApVgHDtdeFTyWZtRjIISe+hxg0N4
elp39TOrzm+gVDDQL6C6We7wrt54aC3nMfXRClM9MOkn9OeGaIRUg8VtI0K+gkTs2IoCzTjlh2ME
MotQJw7TCM4Ndt5eXuL4reAvfABT8pHRIWiMfUUwTUEFwxF6MpQmpgnUnSefO0A4qKCkRIgwIsO4
ZL/jzp3uXYMcX0Yhl8II6C+5itmN02THoU6YGUS0cgQ7cqrFu0SVrscwFV9s9A6OPNhrFB7S4oyJ
3Z0z/E0IQ9OJSuFJ6sqs105T+hfD0+ltrB9LSiXLtVgs93dvfbubHBm/2tdRRk+7W8nrdhUUoHRl
27eTSTRLbtIssqYzCxXEck8CzCI/vRDfhQ30kewTkBAWS4w5OBx0ggLLdx5CsZBAonpakX5y3i5O
3f98KF3s/PFBktAmmSCO161zYngGvUHJb42wtVktM73mnxwochfmeK5RP1KfxT7EbiclqMHqm8yx
firNd5/9Zte9sNx7qzyLsx1Ka2lHLZw4X+WbQeKGzcybVHYhdxigFg7YPwGPzFR5BBUTGsm4YlUn
tTfwZ400hRxbOtyWQOU7415jaqLXHSSpTfLnH9sGnWtD7IAxkfBEvSMy5sZhAMTsYUPe/xsyrReZ
t96RectdprCn6pAzA+DcT1dNS9fG9nztpcoZzeMTg2BnfW8y4tbwKae3FDfAESpUFBuO6T6JUXyz
izJ9slDSGX+lNEXpoTfVLZXOZYGFOZrLgsDWGiJ1l7hY50SuSSuXr64hTXQc6gOvhfGAg0Mw0Y9m
jw93x/L5RdzFeb7hCguB57BusOSmBAgevmv7iRvcyfB2QiqJ9JCqYjNAPMaE6c0+JLbCmqRwYRRr
u0fMwcElaGpP8CZ2okQFsBmFNpEe+G9ZDPi1t/eF7sb0UGaxxdFkc/DSrVjRQNmu4aPH5y7Nfcbd
ncfvYij2BSwWfL+ewvrH/nGo6tSxTMYl6iazfOiisLoQK3tRDkNJO7mAx9pEWUj0+9b1YA1oElPh
b2Ebfv4DyVZ5Wv5rSU+VUxqgfUS9/ATIT3eSYaMUi5Ej5zGNot9RdO6mVCVSweckmbRqBmg1PH4u
pktnDCrf2u70RVmfYqdNbE0+z6JVnvqB13LM5OIoNHqLVJU7nkjfLLIWSmz7rW/UHvhwA3RW7ify
8biIAcKr5u4s4lx9kQH9nj7UKZvTOIXr9dmpw4ydEvxVvvEEgqpp20Jw3E6QWj5miSDgVRM1Z29x
0EZ0dEWZ2jg545jYowMx5QH60jGo7L0G5S7Q4iPFnSp2KNoLiaI2HivZFLzhnJZ5tXXoUjMPWEpX
cJj6+hjMr9BwM6HwR2a66IenGwjHj7mQD6J7YDc1Eva1fpJbqLv12b8P7VfvtsfUBOUjec+FmZhK
quv+QPoafpKTodqhhAUZiGQPvBteyAaW73Speg3NYfqhRaMBT1L5VwjVDc2PzTfMdOtJl7P3CqlS
XOnPRGMz1DgMtDHS5GOQyQ1QBhl4ZLuN7DKwVv/BUM1RfHdeMx3D74FMuWffXhHYCfcvBrXIvVmF
IAOpidM1ze5cSRxfAvG/xwtwKzjwJcIiC+jjN2spbQUSOagZ2f5UamCoNs7G+DS1bhwAcHsLBJdN
d3lSqYR48DGqAow6f9yZn2UW+hOM35o8iyDthtQ56uVC9KiBBvGtdFsJBbmeZhHD4FFy/ak2EXzI
BSMhjjHCbm2cir/u7PENS5IFxvYJEcOhMzyPdOpU8fYetMUlQYf76M1RaPLdx+RsQJejO6ulYgcV
AoEnWEq0xZaZ+XJa8uGr+Zb7qyL/Nky7ToRei+qukqk60gijAKDtp0Wk+TN+cqJssSsQeMk+3+Tt
YDuO4fkz4W2881PCT25hJ9ibR5Z262W9NPsGIKCDGzVaNlRYtQLY4yu8HL+zx/IH8FRuu6L7AtbK
+yTE06RXl8DSJWLRRPN2nQFruY7m+73z7byx8mK9MnMvSwhHc2cCMg2Hfj87d3WKs+56gljp4kTw
zsifIY1WBGD60Zq3HMWyee1uCGfZTe9OyN6PblKuV9it01t3ikzkS03hkGaJCKylcP3haeq3/zwk
pTzxJtdUfyz9WsUwz6u8M+L9bBsvcT0Kc70QvU0YMmofhLQU1st+VxCVpiylrqSrJFCKHLLppc9D
oymjXLn8/aXbDTHP6tjFHIZ88vYp94kF/YrqzLwayNYbeQhaMst5Ckz4f9qgOHuvjV23oV0cJdtj
/5FkWQoU8baUQ5SUlS/0jF6LTxIB1sB2ush9ITVGsLqMZkeA89Tnq928FPjbfMSCBxdZF2fvzu3o
6eISqPNAo/fg8ysr1VZimUN6f+GKVHGBW5J6aoRSeQ2sop9gneiJt2nUrPSO8cP1ODt4qcDPxw/P
xDH9rO4maiBk5jIGwObMt5I40AqXBDJKquqGpoGlDSNfExksJcfIZ7wzJEXlTCwrFPNkfVKOO0Dj
Xe2Xl8PBqRPAFJmvuI5uoAOnwVgF5pH7G89gK3pKZFei30fXkIMKDtSsXFtNsNzzvpTrGUd/RNDq
qJ85lM+g8Xp42xZ4yQnlLqwzl86vRczn13m96Y9cSa/SNZ8TneBYpRlEjPu/GYA8Y8Kv9srvBPQe
6OCGDkWDq+uyaHlL6umpk1964ww2unVewNxCBforAifAfIJjSD8RyRvGqvSYXS3tCeXfKjVQw0ze
OtcYMzbGYnlHci0BRvTUc8STKIGPmoruxytimIP6ID+UBj7sU+Kx9HCJDITOyqV/0d/XCM1QW938
rUTCxY7HwjNX6RrxT/S4gsnpETl0oEzVfTaKDhCXIgm3ekDYzdYuJ/lyVPPvpkg+HocvgtqB8xFa
QCS/yLLbCVrYKd+8IdIBMCJ/EroYa2pGxy6kOSK8pSe+Crk3fxOylhFlNmdubugqCALGeWffZVPq
kKnlcjhZM/ErSW7kJSpRCDlHOJzkvg4n1UCH8PEkWVmW6Y2KxxaQLk9l7uBZTkcKv/B++up+oJIZ
63FxKEN8Cepm1ObNPyFzckWU+YgYf/tsdyoB+j5DtwHP/+nFhLBdtI/PVxiCcNuJOZgw3XXRZkci
Hzm2sZsXiipCN3L4jj1O6yU6ZN86Jho9N7xES92ZXQXQNl+GM9i6RDAdX4fP9SiHwKvU26tKDx2q
1F/JBxP4HbLdRqdW20dNZe+waXLsQofskEL8JZjpM30BHdK9YMU/Sdi9asJ4PJrSEwEq6cTAEUj4
UymnSFomSPm/0Je9rwZn7fpSk7oMWP9m8sLgh943m/pHHFXs3zzpbGvHd5IBafPXpKewvOdb2cy5
VzxYiMpcUbadaWHiBaYH6yvcQSOKWhZglsAUkiBnr7cMlBSixwoueAKJXrFXmZFZR7gdcJ38q1T0
BtU7o8Iz3TyZ12fCvKLxjc8DAt8LnsLQLsHnOUH3sZUlklFc188S8JWu3KHitUkUlB1E0gjEGZvT
z2maRhwWH47DgFZsKLY4ovUplWREp5wVm8O6ydgkwVMEIfPoz22EQwksQE8cqqrwTHz9Kx2oZmBj
oTaIpyqbi7GXLOz+EyFLV1SPLz9f1osA600CTUnFqL9JSs4ztK4NnGRxZWvUlLoB/JHlbcz3iH7E
G/+Tlz3yq5U/jpdJcuWey9D9PfQtgauoLwz3wR7L+fASV5QhPEDjzZJbGf4cGAh46z0Bzo2JfviA
FvgE/Nn8p7tCfLdzrDeg07SBTv+aaLeh3RMoYNVJ2W8Eub06FrQe7ijRIedD1JxF/9kP9JjQRG3w
F6IzMzBMg/Arq/9Abs2odiIwyS1NOpZB/maYsg9VwphUk4dgXWoO4EIDqDmiS8di00F9p9N8psIu
Py8+LNc0to/LplA+IxPqvu3pieWChr+K4/gvLmlBuxhvhuIkEsRw+vw+gm48DyI4MV42gRj+4yMQ
cQze6oBYfAWoUUoXgE1LrceKTgQzT2OFDe3XHqnrwce/2da8Thm09PPNhaq9iprEqQIylNMhxuK/
vR1tzDnAee0Ru9uPL0m5TJkHdVPmMoTrI8R4EVd/4ndEEzEZUXYeBfIGwfDIfQBWGvwPzrS+FjFU
LlTUytXULnX2hQf8+Si4Js22/gn5dniuKiqqjWVyl5jzKGzU8kgi/IB/3kJwLhrNHYZySLnGtFaP
rUveNMqLjcGTeSkOca3N+cerzir23D7VCJWqBe4S47xqr98GE/MOi9Qhf1SxhnEEVc2PuOMoYlHE
OTyiZxUhOBnWVOmJiHzz21qkUi5ou/oahlGLk/vNQU4zF1ImkNv2hL0LnV+rVdjk/nxSdnF3CQc9
gRnqMYrarNFaFU4dhc98hpVLSqLc+fSIoVYibWIZvNNhyGbFW2NYvG63tP+N7Zy03CVeZ11IZLgM
hI2V5by4sNtYGKO0bk3syB2noFxbbiN9E43Y+VAU4vKBoy6H4JtFPC/QtkJ/740DxsZq6fDurwxK
LY9G5CoaoDk6I8TJPxjz7bPmEXjSGiLCs4Etx4WuLaKFIc4Fsc+6uitsKA6Zoq3Oj5biTp96/Lyh
NbqEaPenJ8oXu3NLMQwfBfYN7AJzJmKLdqS+jpN6q+M2BM3ZGaK00IpwYHQuPohY9jGSBLuoJRcL
C8nmjyaq7XLNnS5o3XBO2temKMpbgPrXJoij/KH2KPbL0M36lCFD3qWLUikoU0bSPNwiEvxK2S8b
FbMqGUFV/rCEoXrRCSEbJdJIPlm+wiYREA09bwqr4b5uRLWenPuFPMdNF294sJtUHbXuFm4y4fbA
zYYWuNUYfF4GwNEWtzgqPeAJdWJM0Tkfaey5/8ShnEbBUBbzj5IX7VZKmtxxA+RkvPf90oAi99ah
h+WRx7fqllqFrB0entYFQxPkk4nz0i2uRt7EhyyVEuWtP4A9JJxIyeC3VlTW7OYrDqPqAi5VKfKV
kI3W2V6uxE5j7kxrNdu7ulrU2BpOTMy16DvBY7DuTJhjUz+55SSzzUgOh0LAgr26/nbQdP/Bhv10
B14LoCn0uUCyasA1xFpq682Tih02KX+CtjeYeSTnJi1p9YkZbNhwHWW51VnspW0xr/r/7cbpqF54
grQbF1mzKxKqF5oCluTjg8IgBpYtBajrv5rA7VwxB7J6YtfgV/1eZi2CjcTXZz7tItn3IK7motkI
mgDi547/Es9nsrXgCO7WF7/66CG2miM9LiPpMoXDLuahXBYwG3r2ObD+VHZJvezWgqFmwps/MNqm
ltslHKH+tWTU6VrfPjHVthuPt+G7p2WZqJMr5hMpMdYgGSQLF1N/maQXCJe6iWxDQUy/kwcC3R78
broVLr77yyxqmJ+r9nCdfCAeM6LdJR2QQRcm/+nyBa0Q9EgNKsplybi78Eti+j0ey57uYGOdMrar
nxyZ2YB6bxamn3tY0P5n7ZNpL8HgvhXzDHTso0km4PoBonVDcuIUrf1Kv2kH537lXksVowSGk0GW
ddeE6uV4p6vt7s0x9vOT7R7Su+lwZQjw3rfv501GK0ala5a9F2U+RAi58JwJrt9jtpkI0EubrReW
kgzwME8acCR7+ArHUOQBPdenfCjZ9s2s88SZiPOr5t9yNtnmMxfAykZpF5ctn4rkJI4iL2yAK74A
3hyLa2yn/u2DZx/wKMwhgS0IpeKhMDbW/0/qJSCKKu+IZTlnohZblu37QU3KIdHqgo4pM8kddIco
tK084ckJGFa5qG6vwEQnh5beRawGFkDfWC/V8qzlmgc96Oa3pWTB4j0F77QAEkVbAdR7q/WpBLRQ
mGqyfYK1PdpX+mlOC3nZIOyfbJwEqVjEbwMCA1RYqo/lSknOT/iTgIPj1GQ2bs/hP8OBZHnOv4c2
97hsvysV2Y2j1Na6Be2DtUPO9mC/CNtjYMPp7ueqkIP9lUN0dE52ooLovU+yLICsG/UzURQkPmKx
E3uvXyjUNxs6WtmrqhSKdYjP4ujcxd9lCn7Qal/asiL2mjGgu2Uil9C7T4mhC8dt6WDVSUcbAB+x
/znXoq8BdK/wvGiBCqB/vTTtLpJMdN7MwX/96evhkfoZ6z23l1iqdAIonTNp0rzm9hhJRFWE9PoU
9MxMemkWUOuzl4q3fOZnx1zSYQhlc7/zUutMPv71NOmyakJ07P58WIx8vHuAvGzsqZxd3B4AeJK4
lPqcpaZyxLwB/JRtm7bir9AkTRqVaBVW7114F2GkdCyz3VXyCN6CMus6slHKM7zcXHecjfHAH5Z+
kFPhB5760SD7oK62s9KsOiO80KBO9vfaHmKpmTQo0UXI4cl0doc2zn/LM/x+tVvDpZY0ulwumSWl
vb5BpCPnjzKrleQuvSkcVr6TaDJ1vfjcLMgW4hT3L5G9NTih/NEG59trDHDkhhWhMiy7Mxa/+knS
eTyopfELoNETiUyMdXemhr95288gypp2g1YDIjxwEEU95MdLrV3oVqK25wtpSZBxD8UUbQSGAVIZ
P+1r+avpfHDy7RIYVD0vy6MrwVRSz7/b1ZJQ2WGYUpuZQaYh8aB5Q+Khz59ttQhL85iKQgfx89LK
hjc5gtEzBzSyNPgfwTg5ysEJFhTc4+FzgdYOvs87eEsW50H85aMK4Z0M/CJ8C9vw1PdH0JN0s8Ns
Bpa4W7nHIMTSh4IwPQaxqwaInv8hahn/iV/fSvYcQl4/1DTR7WhQowTK6d+1n1c1vejad5x0OBAB
L59nBNVjE6V82tte3dRQwPWHGVVRZtS8YAjJBT+1apzfsSkgGdyWoIR2HQoZetm/waqpgWg0Vd4g
lWB9oiCvj2IYjmYOeioPppqcSzwxfip+clgQKxg2p5De03XFOiGHFa/5uQZaD1kbv/t+iv/PwL7a
InKPnEENTKNh0rQ7WFK3lcPb4tqAowt0R/08ZjaWFCXeSHS5Fe2b3/HraOZaRfnem4LCv0r2E5Pp
lSPoCarfyDDJWSk0NxXvyUpM7leb3rXr2BEbOi1Qp09UZf8D8lgysuj6qBlAZzd0LZfnTdIs8Q/f
gp3OUT5kQaPzHJmrNQgB9TCEdzru2nlWO9F4vqKQ7sdP8CFkUoP1XX5YBTwJVBsMaF9Z9tSU1u3Q
F1dqJk+I7O/vLUv62uLZeoF2h5yA4lQbwcfKNTqV1WhwHyXcpAOAB7vMzwaYuPtf6NBUWK1iKUQu
irCxwMTNPphHkhISejxj95YaS0GfWw/FRmwAVcGrDSEC+kZ0A5XHI4zoQcTp6899poqV3m1KeBFS
NVBqYoQeiONA5vsfhKxQsHmH6jsqeZgxNGKjsuXJEnj5bTHDiF2ME8oBMLlEYmYidgNc6Hk6p0aM
jUOXWhaK/E9iCeMRn6Cjpy715haDsS98MUT81GVw9UMIhQNtNspYnK4DJRq0uhwpj5SCUfx6lk0V
aUs+rOZkxO330DPpIne8LvatNySzaoOxRObZwXy/jQT45QZFj872f6RwUep4FwNcs4bGe/nkRr14
YRhfTWJ0vp/7TRkoarpYU5Ih9DzxGCibB9s/6SOBu6BRHBuZDYnMepMOLxJjyhiZCpTbGvHL41Be
ObYsKTZaKKZy34FCNaaUWne0+APK+b12L4U9ILFz0oRb9obuO9/eDIvJEHI6NBnH6bNvJMA42R+0
I4ECyz7xQqtXt6jLraAFR3oZ3AcJl2LlF99G89tWQtIebGbhNwzRlGfv7XJCkjdJEsHyu529346S
wg5exA5/dBfL2CnC3SkBPfaT4HU22QhyazKrPHOIB2bR+M/CgD3IPUSPfZhoCFPktPUOpI2Z/E+B
kLpQBr0AEFUsScNecNUGn4/RbsBzlwHvlY2T57e850uKL+M41yTB0Wu7Wcd+dDJYFA3KbJK9Bqr6
FTFsByDqeQbE/r+vQjKrYJdwk8/CNyIXKWXN9uxLIdHqQNiByr87Un2z6oeT7cJzOEwtHrQd8O04
Y0/XGc9eva+uWNL239sgFgr6q8ClWnSDY90zSlDVmjgmTI2CMARRovg0XVHa2LyygkbHaDjbAd+2
wcdgw5RnYoCFUsXYKCMSpSjmypSLRFoGTOcYeP2rktnbnp7e+o1YI/vDqehEBmE2aoOVWwGxDnvN
bOeehEgXPUJuhsyxfYV7qQ6krodJkPKMwRC+Lh+h+wZDQqglweMNU/bdqBOz1SUEI+wYL6N7G3AA
HjF3E6UjBdoXE6H8aFcVCUeDWRQRrGZ19EN+V+09MG2KqTxnqwjIAooFNEqo+4kvHxoHDjrljQTL
3xBkReiI1dLxmrSibodvqnMQtOKGLDz5Hwy5NTqhaeOJJgQtQgO7OjLC4LgS8pPcX/l4yNXo3elr
2xOkNyapmOnfzxaa7qrZyBgiQMOBPXA5lh/8kFgmuVme1hPTr3zIIVazfa8ADXG/N55YDsBtjAFe
WkuGJHnrWsqcTXdjKgFNrkd/lW2soyw43eZtYX3XpKJejKQCGTGCE8s02V3bHjQeXnBp1elC594P
QfqiEA7jzUozm+oMpA+kLStVVS1pETfKkXLu21Jq59w6X8/+1JVxu8cFni94ZfT1R5c09B6G6v9K
+wICXovOXAlXrLKnqx74X+oSuDYsWBB5YaM5pIeCQund+XoyXwxTiOhQuIHfTtYJJ5B0Y9wot0OZ
DeQtg+ubcw6EV9nSLfcr/yzG6iVzl97pdHyZwv/hJF3XA4SJFkvojlP5skOTJ2IPGsd5cRF4Lmx8
q3u5CkQQH/sVOXuBWTy+ODpNqciaYMl9kSKOX4SRuCWcXhPpK1BkDQNU7jB7udDVYARiEx9c97++
XBXs2mBKDOqyrsy4QddDnTw12EEeaPuKAam1GUrc0YMWVNILiPr/HxXvv1eCi5Ou60e8g4niq4ze
ekSJUIxXVMg7XN15JPS13yR7u0rtywoiRS3h0GBzv5qjHLqasB8ARQ7BpWDnbE3I3jEK7/iUBWxH
qdrjCkCgF3E7VyKSb5TBuA+monZ36aCEyxP5Z1uIWxNi0GxcBE08Ie7GQiR072XL/UNDvXH/0ZCj
NlEzbETXXLq/Shc9A3FiB1Z9V47Cw1DBnnN1vKaaG78MQEiLLklHtr5v/88b9IqRkxteCzzvdM2a
gTD0ddUv79p4x9K9a3kUBTTutXLUsK4UjGUadUBQo2/Kxe/yNYQCZHs9azr8TMhZanT9Q5Jg3UkM
CWtoqnTrvkS6+Ld6FskSytlp2m9ayAl34H6RPUWv2/8dDmVdB/dGY6+9gG4YabfvV/15uLCoeOGS
g984Dzb9G9688xWxQ6ekAwrCZ9NEM1tEpw3f6hMMGl6Kv0YXwcVEP9+ttaxsdTgSTqL5x2liZNSh
qYXw1bNxYlaTvXv1rc1lwJc3s+jHl/t/tp8qIPzkSojMkYWXZ/pDEHDIGu5l5n58GceJYtS6dK+P
Ns5QQYHvsroYhy0+cU4hStuDlhrFlFimM5s6n0vOVvCmteYlcENA98Em3F6yyR7zVEIIxZpxjJWW
AL+immkmOWGLJvGxZJjHxz+qoWSMdFzubSuoOF3qkQVvA88/f/xNnk4t45IGwXi+KKyDSmrxA+sA
XS4dxOmRIJdqopUej/U6nVlVzgnGBA0T8LM/7mRx4Jrzwq0Llb7xn7ePZ2xb2Fuh88YBBvAgiMm5
KXwgs7PNos4ukniFYHX1rQ0iP9O29+M2cr9+4H/1rsMir47dY9DTrID0CynmQqZkmKQhd8WhQuJ/
antwlWcdynkNcRk279ee8heEkRCtIxCN8BLt7wUBrm2I6lt8XSt8MyAVfR4i7r6XAYkmLZ+V4mZP
1hT/A/Y639mzVLOVfddS1A+rm4qEJ7zk2AFZSg9EMMDsEULUiCqFmKXWTTcmnK2/uCBTy9U6rCDa
C6KaRqsSaAw5m14NyuS29n1NZeTimZH9o9Cq4MNwM+b/fgQ2G6si2Es7DvjAiNiIILQmQwkCIv1h
+U3LDOCnBmHY/VSWKx55lcEFXidYIwS3kBFAYX2hbEUMuLKctxlIhQoFyfwFYiFrfPi/JqgFsu70
u21wc1uQjsA3NXP4042BoS7BcI3kfqFxXP5GoqjKZ+WjWOfj4nWG6niX/lmWCtoXzmD/IARJoZXQ
ZBNRebXQ10G1wSoZs5uxQLrMYO28QpMn8gEaM8uaZ82aCKb23bFwIK2eMrt1avbQj6hKGuM8ofPO
CHcp1cpFv+uZQERN4W7mj+ZrOVzrJA8R/AtUlzc7UsMVJeWWLCqKTXUPLV2uHp9F+e66yiODP8dl
BIn/RijzARVYsXtDwY58575soFoMgqh9rh8r3yt/KT8VAMUpP4JcQMgjxKXCTucD3VdZfkK8bKLW
rbvANEEsVVkuFwQIg3ujkczdfDt3/qQr0mxjYbtJFKVdXe0uHEnavnC8Gse5XzhA6OD8h7yPuLvf
jHVykHV+a04ZyDj30Tf//erP9J1aEKDnD8uR2ZgbpIPO0ZkRV17wWfj2qxp8Dg+izSp4GjHBVRXV
AJO+JXw+2zZQKajU9k2hChohgPuwsHVIxE1a3XDyUZhlMngh7cCuDB9EufLR0HPMxQrJ6dAVe7Pn
A2wivlEyRQy/ynP5H2EIWudJhuRMIPjF40jGvTHzUqAtBOYNHzKDMb47ePEv2tt741UTYzYMo6wM
IIrx+8s1nhm64BCZ29puIrG+rdwdSOUl+RKqybt37bL9pPXh0gJ2jQ8r7Plgl5pCh+G5tG7BwwiB
FBPSeJxAqq7kR6BhlVYdGAf8V+7iBR7khwWjJR6Bz47eceFuDoPwhlY6otRT1Bf/I2wjRmr1sQ2S
H4j7EKqjgBCBIPL+0OVD1vWjvPvn+LYX2Yu0BLmlhGE+tPBgrl29fErhb/jl5IpgmEXojR+7KOQJ
PLekNORjRYqJCBpDMEZPhr/bOURW2fT4647Y9fz7lLSBv41gEel4XEEBK7T35sTPn9uGsPT+nkCf
gUMJ6syEkDr2gmsYWTxvKsYm0IUZu/F5SlVBZxboQ95CiSXF39FUtyCfhJx6tMKBC8C92A3U+OTt
LzOiDzbaP/tyZRgmXVvifd06OQCvxUEwrbm2eFB9qYEQmCRqx7CsifI+yFU8/qqMQxrxgrcQP/nv
DVgCFvtWH8ECHCJ+PHprl5WacWf8rm5l/1M79eDB8SrkzyYPSOcOkQwSyl4ouC+M5xBwb/J82nIp
RjXIlVZuqkNrQ20KymiBdJ1O5pkT8NrMAlpQl+yhDFQ6hQVQicTGQqz6Al2+YRBqzbipMMw+R7u6
8t1TUYumRAzAdeccBvaKSA04Y03o7NRteE04iUqzP77Tqnynemt+EdnZiPTJnMbyjtb5lsee6nys
7E9e431BGVOIymtL2VHKKApjXUCTDcTRo1iGiB2osoCDIZN5g5026sKW2G3qhetlVzFHdRNA2EeY
J6mvcG94kprKuUCFe+8YyxR4XtBmu5F4nnlH3ot/UsCBiW9o30calD8ygYR5kZDLVTlE/vU5tWf/
B/78lG2jAVX/EmDlTytxixR5F2/i8mKIFVu8Qon6s7tVMk3S2QidCo4atpMRAgJYn4jQ8ueZGFVj
LBffCmbPHaYrJzUTiNhC+te33P4mLiiZiR2DXF0FzJ9dRk3+VpVnOHDhq5so7aYNFWUi4vwH7EOS
tje/5eHFi53xU6PYKdCysvTmkamF8OoTn73Mw5jXMaT6ikV79afZabwjT8I6oD4Sd7m1vlf/5u4w
9qXlWRi2nSviO1Q70eXqICtoUhg/UAeexzAWJrlz1G0LG+izax2VHnC8fm1WnbhNEXssRhJskm0H
NGVWN2/MRDxjom+6jJM75jMZoBojsvJdF/styru11qSsNxp5sE78SCfM4vJKU3FotHEgT/5khNVa
wk52QIdpBLgqaEBqLJhwbi4FmzJe7deJJtBaw+X0j7vQiYKMoEuiHCq7hMKsNmt7WrqVllSYEfF5
lQ7SXEZzzQ8t1S5VbNieDWhDEapI26FGSWkVKJjLv8om9BW+zPx8E4rMLpKwq6xxG7bd8aF3ENct
yySapTT6k1u4QguPavuEzCockVgJlAMxdR0R1c7hlaBmB+QFGv07XXAft5R6P1ULCArKYUfhxBdK
kKB78UZvCzZdQBiPvFa744Rz4FhsF+JuitEqQHhnLFZUJRMmB7MIbDPCpUYcgYalrR8Ms5HzYs53
C/HEKQm/pEv7gZWj2Og181yeHQi3QlY+PQT38yi+7Sn2wZ1fuR0QMAgdAMM8pKz2BZHcjQgqpf9M
bPkrQlHTS3pmbLqIUQeNjmWI25dcdWEtmbrmEvRaLSEx53/j8Sy0juG9dZEQYh8qwpEOGXQOaL3W
lpxKFWPMm9VHb2ZwLLHqhFUVYJpp28tCrkjbtjh5UrRwVrKOJMV5W5KSgBwpc9PjYfTH2occxXi4
px4ywbX6ktJi5EzVuLHXFwPwnNBeYTHMypHpOdStD3Xd0BzB0bQSRKryflJpExs9tDKnWSmUy7qD
yvlqkxeVL6WeG38kqYT/5ay7dSMTtdL89TvruWNdCMMkfzcuBgdaYINUPHWXwz3sIQMTNRs+XVng
bd8LIWiyjjEG3uqaBk+Fvg58FX5Irn+z0tASn1PieZwjil9uVVywDTl4CZugDrr8srmR88nZZ2/o
WJIXd49OuSc27EsbjIkjxMCM9wK+p1ntVLo1oYEV8qKOIgC/yiHi8AaqmbBMxEDoKi4xxUsN1ZWu
U3mqIu25x2SXvkKDevdYGXnPGR8A/pZ4y2cB9APFxo+e0tlAnYabw6L4T9ORkq6CkC4QHIIzfmhu
2bFUesywLCKeyOWAYYV+jkX+ioB/g057FUngKrJ2CvWO+VoqwtDfKLs4HQcwlAYqnXnhtL6JXhbe
0CB/sO7Fw7ymJ4u+8mScKvRjkPIn13bLwm2arPSXdaP/eVeXKa5+knXw7bALadMPGmMsMedC6IOv
Jb2v821bwyYkM6HXI64NZW+tZpBk6irOf7hKWQ0+iCC163w53Lj7JUSPaKUuQ3NraiZR32n+ZWG4
Ol4yICb7aUx+CfzaX2baXJOXZUHq5rdXgqHWaFPROSviy9IvuWGmLc+m7gl20RQZ45rWUJM/M0IX
b+5ezX6oX2kOLIOYcGBRZP49ejFuwMaABDfj9+NeKh/zktuACCV682h4t9PNMNl79hGMB5gcJ+2A
Gd6Y9wlB6/SsTlDW4vqpywnlq5upXNlHoFqX0PpuWQr0nycNY5K93xWMwLq/LaccQUdZHf5qcNhg
iMwklX/tnwAurT5vUJUQ8dadaC6pvO7+kiP3VlunQV9LLrIf7hDWHfQhrmeqiYVUF82c7ldgfOBl
ETDkvrBuUgBzEKbRBX/hknt7XlJXtmHs5HY8pKJzredLfSwdToffK/s9+CvLPodv/4VDKgwPKkQH
YClriqvVboPfyBVCpsK24yogw7CULtsT3HXVH/Ri5ZnYi65EQ/sEsCo6adkg6A3fE4qcF5SjARlD
h8rMyCrAdYbnfrELHC3RCMpWhSmHW+4+TZhid5CBm0OEltiVtOu5q/lojG5a6KW0p1XLtgxTypAZ
rBSH/7yfFmPVG+j8YfudsAPKKVH7XIUdyBdzmO3nmti18NbbJ9C7uOyPnJpl/DeZWsQ4grqRf6Em
GnzmwEPeYNN0HHMwCXHzkXoapxZRlBeI7UdcBnxe/XwA6pE/j4iAZ8nRKNdjv2guKugzQWY/m3HC
C0k2khgBQqWAyR7+8oA9YYQdfjHPk5+Lx5aXGI251lHJYKOiANZ26T+Y0JImqA1P8y+dqppA5AN3
0V5dkyqEggFtbpjjuvWonH6TJWsHXQveGPKiGq3VTHgv8yxDr6h92WMFWZFpWIqdPHzAYLFEYgu0
ctm7ROsEU6t/5w19QVmFjRh/ZYlW7HGPxbznM51+uQMn4oiXKHZ0ZCFs/sm3csfL6GiXWcd7HCyx
XO1Dt9TkRCPNBYGQUVWASNnuA6n66ICFx3Z98gPjVJgtJjYQIc5pyLuN2PaapwllVQLRf5+wCgPz
S7XeKi37uAHKQLOqlSVMN5rlphjXh3R9u9JYKvu6Oya/IbRBnPCtQ2rCWoPv/YMDkjtoXh2WcSdJ
paUKhOkvvbBZuAWPSdpXY41WAF01GRdrKt5maKag4Be6j9fJSuV4piCKUG95Q6OSF3XdKv3nL97x
WvauomUyD9hHnVFgn9PCZuBbp3wsR+OOMpR6SiaaCn7hTiHsohJjBLBYm2gxhMAusoE066jsRIyL
LYRL2b/Zi3KHlH3wdx4YV5PE9WtCtKlTmujun1M1ypeKXyC7uThEERYhtLeeiTTdxYgQqKGde4li
sdUYcjvyJ4Uv/ckvimRAna1OFUcHuM/c650VQuVdyBZiXvkZLZEfc6plPbKjzz3LlKjRTz3M7lhM
GW6CsoG8PKktN5lhGEMa3xRxTTrHGiU7EUlBWqd9+Q0gdv4jNJepcn6iPlXLhV4eEzXNdrMJUko6
IiUTBc6DwYLGgr8JThR5J2pyiLrvO8ZKCSf8AjWsaNWKGDc0L3/QghsBCL/UIdqSxr5uwXbUH/Oo
DW4rUYnGte3BUUXLdrKqiQfJEFT+hF1I8M9U6pVpZuZ9Ov25mE5QSfzRr6GrvYg01Y7cnuktnsaT
SPHcvbDvUT3UTQW8kWlqwdfxxVoJSzxfRjMesF4SjGxTV9MSiD6LUphNdQGuyKWatBnw2Iul4hup
7iiP6HuqrvXUQ4QTNsfPCtWBUrVUSFu6S59Ixa3J1tLbxKsuYPr0bVgPor/FI56r+jwOy0kfjIrP
A+0+oyEpIu1Pp8zDO87Cpt4ZX4DwDok8CtyqCNkJt6oJYb8zmGH23eRk42UOPD7Q5/jTuIS6LSO+
NqZ1RFQ5QdSymKAHxrQ6jOUX+Ax+H9FsEMvbi/+dH0BlLJKuWDXyV5zkYp0wvJLbIlVwI+L/0KBp
GyiXg9mI/9MGE20Q/Bx5CdRloxqJyh7z01AK/XSYnn4FyBQhAvG9OeHswBQllbuS+2+8EC6nnnIn
LyPZXl9yemSNTssUpaOg6OZJ/rfq2VouhDORa4hBJ1gPjmKQbQ+KdUTkUoOzMUXBa85oOD1uevn1
YXj6IfYyP0G79OAgs29rFjtSoemu8xBS6ye/U2s6GN60DJqkmfrX1jAyWK/DZA+ekCZOXwYhCrrA
Gm27kUtQXtFVIwwfK8K8DzkLerJ+bqqtfxjItjIKFN5HbMPCjb4d6YYtTkSCIguo1JKc5EtWVGhz
bwgCWVGBQouGQWNAl/+hzOdWsQBx2vLkcLHNDZsyZSVJ0FbN6ZlxWs0NbDu1+xiDjdw7LzuiovX5
xmOniASAeSYoBhaG0q9Ysq1Xcs/k37wYHy8sMJ61UduqIaNDURcf0DR+/9F1eYlg9b6VxxcgxqXr
ex8UXL/8YbWQATjw1HJ0/hc8xJH8gzu7iZjjMVPgp3Tgfa4n3aaxUz9mWbceUlYPeBojKz51QYOW
QLcQWhgfWaH/JxnSILLDKXYLekoGzgmJikmI/uWclFPjTc4ved4Gy8RCxagGHpu9C4HAuOhTkCY8
8VNljhQKfA6RDWtQkXPAX2Te+DikTEVTB62BrNwIzjNGlzesOArcQErcuFq7VM4ujEStiZSpawoG
E3sulLFUvBPlmRoNzvx/pLopcnbAJuvrKjpVt6PqJH+b9C0Ahhc19oUZ3P6j+8rbvLf6Ro0Dwabc
0xQcABcEn2FpeGz2QYd7Z8tugMp6npxIFTf/5d3uifhTDsHxqMywnR+18ufH/J5Z8ObLZIjQAaTw
Q5vh8QA21tM1MhzRKONgfVuEPWPnjHqnJjJRtUjHdFH2F8puC5vdl8ljO6WKv0fLoa+1holYk7Px
sr/LyNl4Q8qO8uUoh4RuCcy33N1nUdLRyPKXtczxDaOt2vfzh7oSI8p3j37T+08yMoCcI6Aqh0h6
GLgElJdWTRRFUZdbUZlHRYhPXxynMJxo+FKkFN94B17m5beotmbPnqxdN/3WqduWhFskaNDCQFWx
4F7qnKZZy/z59STyP7uxOv3U6q491UNrS7IdTUZB7FMbwD8cDxyR1jEK+o+wzEuZPZxais1US6RB
cIuP0QHgXvs2VHxv7uqtXb97SUiOQ4+7qpYIABeQ7JjIYUk2NmmeYB7rr2UjUfBzPciAtFLpKeoJ
RaVVXZdwrxuSbPo83yKraajkRh9iNbNp0ipJnihMD0hz0OROwSwc5wjVSGdirq0Hek7PHaQD2VkJ
QBUV56U6Zps+t0FLmrxm/veXSPBZLsAJowM88+JaBrrUuRmbaE023YJXVHoE/xW7ibtcG0aBPIw3
I3RyTqI+sAe5Briz9wYLQ41Xjte52BpKoF8hVvuqOp6naHRA27qWLiqUUkRPo+0PHwMJ0pc19FPs
Q10cA6FSVUmZaaiOSWCbJ0WgPn5BBPivQBNyTERXLvB8LNebSJZC6GeRkHK7YZoyD7oRbnOfomgh
jexm9n1uXehkcpqyrl61fmgCvKoXhwkN4lTM/+a57K+mftxaT5KyXAoTXQhhTiZ1QdY+FeBYIfzk
qgbZfB8GWakFMX628+WW0/r6ipJB+wPD1/yUyULzwk5sG3u6yMpm96reCWm4qhAiGJTFIsR9C3nf
BJmByD6YB9VXLGQSlhQugVGdJFWD/fzl3DPJyBHiDABAsd0HWqiYXKLJkY8sEXspsdEj/GbtNKpx
IV7zeTy+soeUNjxCL79gBmSZGNPFaTyp9lClq/WspHLlvPQ/I46VnmZHVFWKn+/l9T29cj5Zbz93
uJvOUxCM+laH7qNBLOTC0QWE3n5EGcwW2iy4ekG/hfVSIrAN468LrlLnzdmqCP9U46vXDvGPVJGU
U5sK2hqtEJE6HuWOeIKKYlIlfKS/Or2Ohq3vsKzfSYRpQ2Qs/J5vSWLu15MiSVHBmF3wR9k+APiA
Nvbfdoq/dFkYOSK4UbsjH0FNdQ+kjvOkeD2r7JFHwQTmQnE5vXVU7KgTZi63mPsWahewUZlmWKGh
REf5d0ZdQS14N5FMVHZvnX64cG2dh2tSnZCGliyN2NW5mj48Mo4iPv/TcU6tpWN+n657gh1BXozM
PruddP0/5ZZzduhZPxT0HRyPK4fPAV13lI3RKRUbNO7137hjFBMrFJj+i5qWiceG0n8fb2Re6IVa
2ldjOBBu6AmxxFwsvR76kDaJKnd9rXCa10MKkQ9w0pXzCE0ZM4Og9MfB1uj8Nyb1f4LaumZDETpR
gUtntFzGe4oVSzNjoIUfzwzqff6nZVhcM01dw+G0jSXlm5snnuiiWnhBOeRLxb9UQzEyebP2IZ7y
bwMZ9NIK41FY1Z+4XcDbWcHIV00YpUMtcYqA66xJPf/RpfWUpHsX5p6TupJVS/SWzpIJh3Dpbxse
Wqnikl/ObxOJfz5s6pvrwcANXp9e/EwPUErLvnOLo7x2wDyPULISER5NJZMwIdsdS+f8AhhwYXB9
w85Vgg8fuoODNlfzp5mR3KLt7XroAc2fISDIcjdDx2nNKh63r2JYfAKUf6tJwinGI4QMYB/ETmWb
0LJ4AOqdzayTEhEC/70eMezh9uz/THI9MfhnSd5TaNQeArQUHfIsP0TungJnzLodp0z7cH3AOjpq
RcFzAI2PQZeaZithOLjSmelHzfOA83Q1s+WZhnF9sBqhCmAKJYSgonDcPIMrB1Y8SyzQfnCMsCuR
cQ1A9AuIzhTOBptD+6Uqwd9RHQEUOCnI4L9IijRP4MVBwubJvldJ6SYTuLeX0D6Sb24FD7C2Pbt9
3Nup4aEKyj1FIPIU91C+27lQq9M8e1KDIFtE+jKGX42dOMc+S1shyL57u9gdI2GLwI60EDONPLbE
h08F/Q1Zi47XisEAyN+QaFIne8JKuTJwA3UHAiVKCS0qOs0QcQcuBBGwCMDrTItDy9NNV+5GVk3W
CLpy2KRe3/g2NwmjpDJYUbsuS7Fpe76rREoIxuAkTqSPtMXXHAMsfw9O6dVb03n3jB/VpSq7fs2P
6+38BC/2fGOf/lMhDqcDNICuekS8MzTdLw+SS+8Y9MGph9Bo1ORPlzJr1urnPWj3wn7Bz0Tx7k9m
tGehVYGFxX7X8Bw5fUn5iE5W/26qRyHvUKrDhCBTQHaQ/QJeowNa5w35xzim68O5U909y4ba+S6t
yoL4eVyS5JeQAALW/mEyE/YWTwRtYQnnvEfdlAxezUrl6ynXjUYabTjcDvhlGo+lKjkg/zcvD220
eNzc/IOcn7If0nQBa2z4VOjNtTy4a+Fysw29VD3Vt+pIMryXAE2Kloebi6YDxczA++xpTovy6qKN
DUF8DoRsewwdnsvMiOLAdY4WKAgJCtrsVt4poE0QcaDtv93aU1jWA5T0yHN+Oi+7g0/F7AC3PeMZ
xl0gM1HNx0IWg8smA3viTw098Cza2k0vUvFBvz5ade+Qng6jS1yTLsiCTp1XYmEVRwTNF0uDUaqI
ZMwqvnjnIRJOvwnirgeZ1Or2OfxoZUGToOeYJHp7J+oTHwLSQF+sWZUxgHmzVnBIUi98eVJ3GHOX
LIbMnnZE0qt2bBDYhTFOS/RyPX7G9O1A4LB33tnwC3fSyOnrWgPuQFtXmA/O01MjrNQEoDw1QddT
L0kk+YKryyVPplllbBh9qKMUKynh+iIx47+7b90pLv9UmkFcnRyHjPQJx/zaRNjDrHfQRb0UG/NK
V55KyWOvNGpKrwPpSVzXI10HOhFsnn720unxMX2X42Ba1/HLYTSkjLCL3eoHcBH9OUgYQHIT8j8v
9WszOlS5V2FQ7FuUnKTgKX8lzQpu/RsIBozmwEiMKrcRCL24Uyfu70XHIgC0itMqg62jvu8m54Du
YofeTya/wuWw3a59VXaFTQIRVBqwcIrhG7QCxe7YpiRVsI94WFhY+Gdtc3NIjeAVCgQOHyBLHupg
TPH2pyjib/AyqTWS0+vdpaKGq8Jf799PZ6n4dU7wu57ePx8WseQ1NvWwgVuW1uZi5oYkglWBa/e1
CMlwy9EIkMWG++VJSK4NevSJVx6d1+UPPkT7C4fT+UGuxDkaLsegn9UKOL8lb29yRB7eiV5hd/sK
CEqGzfObImkJnjAyetb7HlPvnEeTXBMOy5q3EgkXhSC+gMi22dxYSiOqJhU7bD33swO+P0EeUv8o
0AfzOT7tQawenWP8QKmW2dgi8FYE85I+IcDakyj9M2axkPQRxC8jGA++4wRYNNQ8abafhD70SvGX
yXTX5E3l5jh3ntRsdbWGqA9TC9JS9xJaablvJfRulgA/WPyi+LkaIJXSJ6phV0ibAK4NCED+Alqb
vBPghAQO36P8yx0TL02hqhUYAoWxbS/V6lCDoaKW747yDRFvHoAVJ3PYOSwByo9sygJzZGENHJuS
jLsYLlPrWSseSk1SUoPay1KUoOy/3WlteMA7yLb6Rhy9BUW0Zvu0SVfHSBajk/YMiyrldF/TXKU1
nqahqys9ZiqAJaML79qPWSBggAkqfnXke5xNlNskl6WtgX0SVxxPsNRdd0vMzTCZqZV3Q/5h6M5D
hA0GzZ7YnxsJMYAJaipkdmuRlyu4mUagebiCpTnKoe6/2Qnpcqf9mbaT+M0knIqHyLQwrRYSID5i
sW5ehoKTEppdjxFuXKZIAnYryoyhDoQ7CLob3avTRetwU41nYQUB+ZmaPy2qkLcZIGv1DthEB+kb
xNUApnz5XYl0iBYTkClphHVBXnYa1aQvfW1IvmZfMjB+iYtlMZ5JB5LN/LBM0mUBlHXhQngukyA8
YEn3Xrtk/F3N10omZWWEWgBfhAC+R0X98QispSXqVFyt78nuWuJhFTvciaT5tITBX9stdvgbaZ6d
yG+eLZmfOUkkB2RRE3WgDDE8B0qSZchzJTl+9ANmWH/gYeHPVihTAnP4XEJB8xnIyQ/IcfOjUTlF
on3Kc8lV5IlKi4YBn7ln4haQVID4ot9HF8YIirStf8QAmpQZ9Vvxv8de3vsjVSPnLS3R2Cwtzhnq
0ylwPljlZmQ2Gp2k1fKPTxfVYm6+XHRQoRi/EecEs/4rZhssmqXC3fGCzerJxxUapJxHwBLZN+Gf
NM9aLMZkqRd25TkrYrrwXSOrSQ0kbbAXlMfZjNb8ItDfqitiyWIgSNV4P8diiIGokdc5pOu0Imjc
QDbk31Vj6T/Ag3p8Yjd0eBTsSUg82KqnPzMe9Bnt2jdE4Aj/RaqC4LFXrWZmN6GqeIyFH0UpFAnt
YRhYUpYTijWcIEOhs6G6cztyDTw/OdcisZdsptoAUevQnWgdrjMWLdMPpOf4Qql5ixqOEcESx18z
SjtJ1VEVwrvY0KSRgU8X5yw2FEQ9bGSpIF/QNpkxIGx1xUdBlf0A24nDu0nSDBQ34nY7XNjZ1KFl
NoQ1qjaLizXaCKLsr7Q9mfUH/lSLSFWApZt4tpG9lr3TOtktKjRejlbnu2RdhyXz6FlNG4rB57bX
wB3AZWRajj34FOITeDNodAbSbjy5qn+438Py9v6d6EuutBaeZ6YeNF3xTN7OH2tWgdKFMdUUIvc8
ijR7ejWZPErbgFD6sjNdSzoYEUmS4rTtzaRfg+cpS15vUTkuoV/JQagq8IA6L+LnDrO9YWXiXmOb
sdVNydDl4txWJLvpZZQpG5Op4hQA1D8reksGmKHz32l7WygeynTjFxMV+onxks5wEDNoH7dikQv5
ryT43VNJCf/Jg9/xan5HQIpoZHdgiG70dKrqJu+42PLCuDY67eHtsbdtiTbOeasmbTaANKmO18ms
K69+5XhJoT+wfexnTdO8DnybMwX1tXHtUj5KaD5VSiKYJ/hnJEApaNYjruhhh0S0qSXCR16hQE/G
9Queh8cePZFW9qR0rOlfv7mIV9K8O5fJJtvy4X3rk3IelhMJSYD6mtilUC4jCxtOv/VLiD9xFy5C
0tOVHvQWRLpS+ffGl8jItRMnOTAxktlkJlaaldb1EjwElzq2C51ZZU6FngN4E5mZtPN/EO/X58Lj
fMC0k/YsONZaryHFuradeMjM0t+obnyMjl4yLxGy4+rTDZqPkgPIgOmLMZ30k64+rortNcx49PQm
Mg7okf8XGHBcejc7B641pjUll2eT75o41f4A52/h9dE8oUrYipiY6D3B+jNgeWjlhEvy58ttdGha
Fle+ZdOXt69Ik0xzg/q/NKOLXnZwFnstisYM8y4L//WP3i/EgfRYazPjHHgOCVgmjUUWVfwMXd64
i2do/QzGRfWVSSsO/Xkk6BYCdueDq5nNkwSeAk8ihejfy9kyE8vPuc7RW2P8G9lemald0DNaqViS
QMSVE2L/UFKFuLVqcNLrMO11pzF1akFv+3dXM9S4dGQpmKBn6JnJ0c5Dpdtrjk2jCxFidLgicWgf
Jb0W26dPuPXRhZQIBctRmYchMVc7KfvHPDdKjKEGbq/Ucci8dDpNlYxuoHcoTV8mLcKd43g+7Szl
Wqw5iiZmmF5uPtpwCXOaNyaPY7ZIyuHYP9EhihgLopeDOK/A2Rq/o3LZHHje9L2zlQP3y5PbRjsw
VIkSxpiGVYWRo3Refs1t+UW2sdVFTXxbITJRMnXY/cIaXbnuRZQfiSiurH2HXKZm7gOCVqRqP8PL
6r5/gVUMG8Fel0DRhKXFVUt4KepGRON3cabTo5RwiFJ1H/5NDL1xVloORFs3LFaxdT03qg8XOl4r
N8zpO83ELk08CnWjoloQjvqoPT3MF5ukV0SvzDwHyNuwze/RrkG4Pyd7XKVS6vpXFWORoBQeHa+t
tM/IMlkZWhn3YVUYE3o4D5EbwRhzrNCpQ6kPDnnQFHP5CVQPmRiVy5kbRUGZfjalzv1E6ODkHPk4
h6LH4DvQCqQ7TKHtQggHCeUgONBprfSsSQkaE4pWdyPo3MalcVgAvyNeeRt3Yiq2dFg4IBPreGWf
o75Y5RZjthmFf4R34JBrB6ET+sntr2jIpvSYfnyKitrqAjHnFkSqLcryoodsR+Xt71YdmOeqm+a1
rk2b36+Gn+Z+zWdDm14PsM1JzkzRgn7xF9C6D6ycdju+hK0LEvA4MkRsf5QWDtewQq6Y/+sp0Q3V
V1PFeJI4wuY/9PLQW4kTOOcVhpArRYNMz8nap0bUhwzQFJPggfkAlRws3e5L4IAzMz0FQhMyrbNL
h3rpNA/Vq5P0PKHhPQdEWJy79hipoFoMRSLaqugbVlG9azxl5yiDxyeI7IM4TYbeYGkEjQgmFfnT
xrNZfwZrFjAMYIXwfjnQdig5JO98TVvdLKvpfOiNnWJoiuJ7EmTFabs/GlJgA1z3u6cG7j3ZJPZu
HX/pQYgNuG6Hfy0EgLFPK+1/Yi+/Igcn5b+6Zg/S8wOGDTnTtDQ1pHrCwGdeUg3Z2aAG1P8STbLE
Co5clnZdSfRHRnWpA7LIFzW+DF2XrnK2MC9H5O4O8TzeP/toIhDiJJXjtyNLqZPSAGICA/feyF3K
X45gQ68mka5EQFGSdwhi5qlVdVJ4cG2dZxg6/exjSSTA4Fmi00bkAP2BbKRMbvKzLi9Nk1KZitRO
y/SRtEXBZiaMAlxIB5nnz6iscra1X2ggiAFJPG8e81tgK7B331yvBEZ+ZE0D+o51vpG8jOCT4teL
3hAuGnvJXFeouAPsEN31aTW5mXNyHn+F2TCzl1+IR3b16voY6GPOgyiJSGQO9d4SxSENrTHFFLJi
vh3I547MkDNkmNqTv0bffJtwSGjNEf8NMCxjNjBQB4b8Jx96NzEgQzv45qvZlPjNe10Y1gGVhhZh
Hh1BxOTTEFCkwwmJxtnJHo8U9scluLouJzz5jzjvhX9PucCrqEeqOORWPI8Mv89zfpUgLCwYunMn
1us7UFXMRiYXNTgxy5a9ZMGEnqoKoWj6WRun8zv45BdB9ShIG0Dyhc+NCxJkr23jqI03SqzM16wD
z+5H43yhvOA+PbQXiw8lGr017bl14mhE0xHDc6Lbx6YdkSRSArd6ywe/EV3nwVFMzVCEO4YYlPIe
F55/lKm/gOJD2QK3s/N5mAVUz0U8ExegXBwA/mMA+cZgIrdolHwjLIIwiA2zK6R18HBxH/2iZ4DK
ETLp8nlGCuB5Jc4F1i9JA0gCFFN4MR7SMpiqgrLTQ91f5/IyJVQETLiMOahGyKlK/Crsrp9NbJH5
dzgvC+h31ZD8VzdQ9+gI02oWQwAhIoAWwfvy8bLtl1wqdsz8wtIT04VHnBUDErLmfJhQUAUpc1Rt
YNgX1XsGhngFQtGjobTTndL1XM7q/Wr1yeN7M3Rvu3wfKYbUmmyBJ24W0ZVqYt4YXq40rgKDmeu3
eUpKc60Z9mdUKKZQtJ48Qd+jp9LQSdjmxCQKF1POqJG/ZM3wzOA8HWbvA79UgysxUeQoH3v/09Ta
Qbwr72ICzUl6eG3YTzOktqMzSXL3y08BpzOjuI2W7Do8bdGG+wf1ZpvcItAMqTxv75n36qpM0HRo
Xt1YUnc0cRBd/FYPnbmSxVihInDvyUIlXuqFcyRov2QvTElSyk7jgWvt33ZP/jQBrJ2X3364ELuM
kQyVPXniyez5v15BY+FMks+/ZJtPpv7upmDuQh1DBI1W3y//jBLYxDEE6XjMbxj/02V4p+RSoCoQ
U1dIpXksNSUD63OelA9kZ88sWQGtoJHMFA55W5BfxfOLk3aqTRDmsxch1HjF/3oFdw5i04nvA/np
5HxUdT8ztYKRu1Tjkaqa0+Tw3UpwyYV/0kRo83854LdivqQz+Ic3deFZIDXDzmD2tHpdANE+N/eI
MKFiQ6Rrv6WNwouGm9Tu7jfgMFSju7WwEaBCsOSBaQNzSRfnAvYX5xpsOZ1wFRy6J/rib/YFHBl2
wxwxUzviJ8bvSEXwKI1ykDEfbyrWvTO7+RaV3++ARefrrGOCykgxax5P7YnRZO15Tq+lUWeWUqY7
wPn1WsGxPZSW1146PQzM1XJkqt/aAf8Gc0z6WfL7v0RQzehKaATfJMFkNNFbE2EafgZhPAg3yaH3
futtaLF91P6Ep3pj0IMCkNJd1jTeElLQSfagg2hDJynarKnJVIX8idkqEDzbKRncwldEMoQmsvB9
miDJQ6CtdizcyL9CekDgikeBV1hLeoj1JYgeJq09P8fI6ObeJRubaYS2ynRBJXmiaDTv44aEtlhE
FiTw6/aX59J7yA48mcO95rC8Dlkie83KaxuxqzOtLDXT/MbcSK9GDgOEURhuze/Piz8i6QGJsYSv
Xxwimtbpf+mYnu19X1bYIB3fIZFH1raTWjAGSmXtomFs0ov9erGKt1k6JRI9c52nYkHxUCv7xtlw
O3tiy1HTIYko6yCw3XF0bCqxMlBvblIETb3srePmIt74wtny1Xyc7KsZAzZSvan0GR7rZr/kmE0A
X4K72WNmWkiheKgcNfBetpwg9ogXe1Kdt5ehIH+Q2Xf5LBQNgFbmxXGOKiOFV2oV+dhwH+jP++yJ
hUPyzYQIfiFFa50eIDX8NzEl988IzMvkr2J6aRiMKM3iaOAEAAGqxQQh8FBf7g/NGBSuo1OL9sai
Gpl8wC0HJa1EvpskUoKe59X4I8L2tuCpMh2Qu1sB5rJP+WfIx+Ju4CLgB1luqVjFmCUtr6yqV/ao
9sUpA9NfpsA0eROqG/PyW5nFG4PHkmdHPbGJkFc2QIEG+BU8WgK/RLgNNV0wqPMlRbekurG3aNlr
1HKa+Qp1SraVV5PZB8UCfonL+/42pr4b5xoR81CdSmaeaUmIIPLBxaUk0Ljh6p0g4kYRqP92AUnY
khHp1yWlKUQxWeRzdgFD6pdl5ENcveW1Lmd3sd5fJH8ES2Wy4lf7/nSoyqRyAj4VMbwX7GGUBJIP
9NDKRFvOkhIYSNZaMTUMQfpbLR1F4MMbfpTlzXBVylO6QEnW3HVJqN7Doh9+9HVbWEY1BEIQdx1Q
6/eyDKrfYAe5BmcwUPuDUAonI5noyLk/vW+vYClFRaY+l2pci7aKSsLUguncBAPp3LRji9tu9EHC
sBF3mYykHxnotG+MeSRXejPWKNAYkB1cC2ZSpnieY8q6/NmY6ZExitrpbDarvZdasQbHxu7egeJF
BK7uOvXD4tHzjAnG2XDJdoXn4+SaHEEpOTAIgMdSN4HGb2lc2H5scJ4h1V9xGnJH/bFAiK3TnvBy
LH6/WcF/kDxrUGXbGS60dIF4EvqToPZM+ZuMZLoZX0YSwemNfM507glAhLxKpa0sRitP9IJPjBl+
tSj4194mQr9f8CSQzzeBCeN6K136/qhT1DN/oUT7wcqI9ynR/03uSn4W0L6fpLZkmly1RxJmlWu+
EtTYPmMvSlcXyMy/WJrDOlEPDAJ49qL6p9ZFYeoTXugko6Saz+fkl1REoPC5II1TP/q5Q6cDEDpk
DG/JDLQW6dZ/hYvQE2Nu2ijE7q0yOWC3V6RKuIkSQ08r7fDKOM2U3BbcAM/Wio/yLlr8eaTt88oC
e8hmDyJHUXabT/8eC9NyboXI5wjNps6M3CNcsrQf+fEBTSRhssEfnWJq6A8/u82i21K83rc0vxnc
/mvFrwXTJgsymjku7TpHeDhXEzm79wog+OPZzpbGNK1zcwXdaa66om0lmIGa03CbOLXYpT5NQ23z
8qqmmIc7Z0FiNcoiO31xEsU5x6fwhKyZIc+OeUUoClUsQKkH1nLTh7Ij3TqF17V9+Zx+67LMvodO
FP4Qr/50HMWc0wV/xQ0lBnSn9/XsoCib9k+O7F1NWP9piFyg/a5rPst0nkICD3PRGMfrMIC6mHx5
4Fk0pMBF47DHOlRNDcBtD4vqnnHs8ZGr13jJiyuW/BWM3cl2KQ1XIY1wES1dh2U3KhiEqaI3ubWb
D0Q352KPLzf1djuYZrkiD92zXdqz3cshklZP/7w1cRIR65VHLL3gFxJSomJCi1B3xs1JbrmrCdA2
dYL59BNXrU/iJePO+Pa7n7Kr1G35wRD+Al/QII1y8SISD3lz4yd5AfDebVOXqI9JwxefGEMB+moL
+YjiFXudzG858LashWjpeD+89ZfaH44HasKiuEe5OwiHl8ZfHHfpZ5uiba2WDj+DVQ79b82Xo7Wr
+3+PfZ6QrYpBNKWe/Khra79mwBprZnvcsu8QttNzHAE1C11s2kNSAn2vgQZcZnontK+QzHHA/fBs
fMau7yYRKd25o5RNvEakreLE8WSoCKrsixzL9H1Gmyw6qn6FRNRC1sJLrqz7kgH+KIydar5oCCHd
rMJ0AgqAro8+wGKz1okawO/VSwuOOlrTP1sz6ZQYn/O32+nKBXUwkAlS5Xx8LuNWd3cT1XH84esq
7tzU8Imt7n+r/zWHIY3HhD/muAVe6a+0OiuM3emsigjCubib2fhbJmHfgjZJVySDrm4GLiNEBT8h
IZBTb0d8nCezfja7VI5fKRDPFxL1uBVfYBiaXegnOwcg9wy2kQM5D6MkC+9kVNT11bwHUwco2aNv
LT8yzNN7pMkYjhbfFCAxQ8yqFB7RjyUURjl4cDJsvPA9MXshGp2UROEjsZ1zVGG1rNXqYD63toPX
UUotKfriyuByaWvdIM4nHliHvRT2q+4cJ1bfqNja2xoqooLnCw0d7ry0aq4i446Gdbv2LJzRmaUm
OwwkSahA7YXosSOIerI0NKgzYCyyptRGt8ZFXDmfBAEvUksWIX+bUZeU3m36fyFcCvBHgkM+LXVA
92ieun0Wb4Q3ySpJQsNP1xY5i0OhzkZQnWwF92c8JQqHcbS/3uHDFUBThJvaWeF+TgSvKGw4vBAp
xh+qiIDA7AzqwszdykKRI+oasOLt5C/PYRZ6hd5iNL+g2ohoOxdqU1tFe0xqS9z6d3c+RY8FlWy9
xqD87txmkOn+IDzXO8V4kTWkXy1U9efquZ0tW+pFzF4BpTOFfl0gVWax5PwEDH8WlHw+lM98PKJR
YMD/6jMPHvBhFsdO9XtJnyKBClrmD7GRpOvfXuU2rzftNdNB+KhDqrWbuvgFRwgGTrqRXtfWiPZ9
pLvZ5GaqtKGio3E/aL4Zyo5naMWlvDAsBmM/Azlm/jlyL9Z6RVqOgjDOCE0eVjg22SqnyqxlnQkn
XFnqdSxigcTrNZlGPOQ9m3YKazC/bWEcgQdL1duYkxqbV4WbcqQmsKvoPFLa5Qd1uO2pHI6vi1WM
VNh6n5t6/ONRrqtTREsqOyy2Yiajlc45IjL6GCjTCbgNo224HhIzZUsCpseIOWAuCh9RiMknebft
lZChaGEAo+WCFpcGEoGlG6YQf9ulB1ST3qb96nCMus2HyeX+U40vPkCe7Pu7zIQrHS+0OxiENhtX
rPsCxexiX/q+xYtBRE6sVyQTBBynYQLmZsh2MZnGA3Uhs0f5BYTQ+bZ2qsQIk5RdQlyFt9UfbG9T
nWG2qhzSfdp1lWUBN2OU3uSCFN/xSBfpsDR2dUHwxHbGFINYTyhG3LXBaaE7dKbIjvwJAU0OCfOR
jtbmtdZupIgTpxsFX6YE2DkGHDFtif6UgZZGIXe5kKadrSU05Vx3zYeNvIvqQ8QYrkGA4GR999A6
DCJfUydulkPl9b4Ls6UbUH/Yqm2NfGiKaXGNhDF+zurJ2tNEb8sPIHrSBWVijH95RoHj+9rVCK1i
Kuq1SUZN5VzBA8mVoDE+RR0rIZr9LbUhT5j6gSDiW04mQl05GxaX1xjf9s/zPQQVbMzh5uSwDn3P
AfQFADJj78QaznY5I9mCL2B6aE+8IkV86eGn17vaw6Jx+TW9KMGMBQ7tH/RrsCGJP/NIDm06qX2x
RtjpJtCioEtVlfK1xvvEXwEr11jdSnT1UVx3zS42+QBHh6oH9BmfCfeKOZS1Z2IedQ/gc3y4wSd2
+k+x1NtvEUsPY1+3ag8UJP1B9WSKHekfakEM8PV0aCCrP9yRKuCT1/ZFDtSC7R1269qw8qtXnXS3
zUQRzfXSm7jPgvVI/hKAPWzWJ2glnF0eXzqLgZD59Uz6kYeiGfD3Lwu6CBLdVVZdhDOyABn1ZQuQ
w7inDaoc1kVaymEF7/rcePIa4pR7o4RoXxwEe1LGlCtsnoP3ss857idqK8VYLvzT/WMXyXzgc81E
purqO2WqDSn4wd9p8LYGDvHDa1WW7I6sQh+WrAFjIDDA98zDsHwj8lg9ocmbXebkdaTV0z9koEmr
hdOMG8IsYYLlq3ajDZAck7Q4787VLc3vwhf/l7QOFZwQPA7kUoMKuHT4YZz00ngYY8gk3leHQgH4
9ajnQ63nXT7XY9WxdPVN2CRnZ0C9vChfZpnOro6wTLPNU2oijEWbd/oSzjFLn8xGUKlmvjMtv35U
tEfFvM7FxGGr8xbjrKsIRiulphQtgZyT9N74HpRlx7bINHPB9/AByq8bh+ZumNoGuJLa3nrjpFAf
UbJPXFbL3shprjF6BS4AMLJN3fjI5Lc9jijSUnNJk69VgN9s4ZYHkRa3aLXvv/qauTn+46buf2vT
59vGz+cUvyKdHQrMJMuooDTxRGHJDFIRMTKA5ggEgQcBq+9D8ioLNL7f8+7z6eB9VpmFGYYhMgMI
HEdZvWnLnQuW4oqrn76AoEnsh4c0KDwMDzBBFcyQ96/qnDduiWZ06RcovZOz7fFajW6VbUDLmWPb
IjQlcvZzRrZ31nvXpQsgtN+6w5SF4s6Snts+RZnycAcU+UfiXpEaYrYtMs5txfAqHRaJiwAaDlaA
8EuV+h/lp4THyrqkFYZ566ciE4EdiFY2aMfENA7jnzn7PH++i6gzi/m1MeD0MXKMViEhxeC+ZDYz
yvnPraVKEl4CXZijefvoOlo7z59IU1i9TG5llbzFegTPpInHC+g2RZpv4eVJGC+WtAK+dDPLO7JN
B+Ht0P8JU/K7BIviBEA6Eh1VsrJ8Oaovz6Yh3skrKiHyBRo0sWlpBD5znHlHUJ1HGUT1NtBObF4I
/M4dHs6Sni7pRoKIKHW19zMuWQblnOyNic5d1InqBeVPFzg3E2bM3H6Rqg1kHlKNATVh9tD+QYZ/
ysSkydGGS5e3zU3XSeOSUvrO76xAf6dEChzWurSh4wgeDmwv9yzCoppYBTjzQLBVJp3lAzsvilfH
miMHMUyyGDmOFJFktetVUkFRmCITqFHAu/zoFqZIlsqJbFqsHlb8GuOes+dFSZW6eY6/qtGR3e15
YTQqjxkh55Jmtqarl/UdjlvWwRQ00IUrtygJwzxfe+13DBBJK6PbKDM2BJWEUABV/WA6adwsvQnN
HG1PjcQMCokpMiWpXcS4ud8UvWP4b+18eV7dp7qJ+/qaDqr9dR1LWwCX6J1qaraVTo/GkBiAMtKk
KHwHcOlzAvtNgKb0GOuVUT3mMkZU+A67AKj4/2IQmoU/xsaoqvUGTWkCkiD9wkL4ozGUAQCu/GCh
9rbcko81s+6Xt14BeRM0w+JQdxwy/vZzbtS2VbZwxQOCa5BKdxigI6wcAd9UX1FynUR3a91GJFnv
7CayUrz9TRquIRGQit3av3bxACDO2L7uPeUGpCyzI3iR5l/MZHj5reeIWWb12C/fnbW7wF66tPzB
UffZWYwI+BRWO84zZgQT2TVb4SxIz9Lb86seumkXRP964LCGHD4e6ShuX571Fttb3/sQhoBPj2Gp
2rJv26Kap3DgaVYnz7HjTRso6GT8NZINQDuGNHziqaAppNYdgWohSAra5I9xQ9+pEiy7xmBoSozi
nTiAH8hP4FQprxTqnMMy1BsN0+sy4DNJNECRPJOe2QlrU/7I2hRr5M0xMh6qbfvrIFPYH8LepRH7
CJ0Nq0i+YhXv8Ef2jQpWUzk87Tz2DG7Ai1R+8dcRvcaadKS0EaC3Dq71zlFRZyw5YL99GlpsH0dn
NShGRu+6ja/GWsQLsF1PUIKJHzyGOBr58RYScM9Clsb1/PG3eemqp7rBPi/F0o57EblyocHtQ3jK
/AbSEal++Lt8oGEfVuebnC79s77x5I69YIR3T+qNpX48+yZXb/ZtBTOANNpLcQuuq1mpFP7C4Xyx
rawvcJbMPSVnheUcb/3EL0IrxdoCk9MhUjmTC++3JSMQpNSTVUuYRMTEGNoJrNY7XKkEDgrbKMdg
y0aDNSk8POsbSMFTS0wgjPD5qOb3eKoaIlsLzXfG2++3ECxom5XfOUOzk0AsU6TiG82goVAw5GvE
+kDFVehu8zwVVBIfVAHbo5ApAAMEEE7ZcFV043AYboH7TMI7YjTox5P0zQbR1pfOZtv+BzOq/Edm
w0YEyf9QvIHUsjKwxL1d6gclhoj5qeCYc2gpMyNDZeaN2lWCBqu4OS7tKBMSVE3e3hyjIQ9PIvxm
bUo6JvtPxM8Cyx3eCqxnsxImRLp1bm0YBrroCki5iuotjqqv1pHCIUIYINqYmqq2YJ+7MKO8/7yY
Ri2UfOE68VCa0mIQDXOMK2WxQ/v+CzRMm/na+kYABKOIqskh+7t1Piz4CYCTe0t/8k1zl/+uaYoS
sRDVeQ0r9XTgomvIBuryuaIJuqEZNdnpaaBZrI98JI8w8SNegZ3Ou+yWOrrIGY4EZVtrbFnZdzEC
HGD0EE2HuhhIjw2O4o1ArqDbO4OswjOkFRDRQ383NWND4P/acJlKD+j3Wj5zW6gLFQwQAv4F4ENk
mKcRAX8LT8bih1e8kQuROECJjXjiM0C66rd/u5RxhwtLOq/gNCzcLWKItVYbX85mrt7JLVPPrzDl
oKPEctXawLQYnvJn3W7koPvHF4+Gif/GgtIPPgeSwNne174C+iPyVGVJslCYWfuYKaUmQGZl402L
5V1UT4ZLYipsEyD+0V2lHdHVVMjorOSWCofACT6MKoAUoruliCNOvnAwQt82SUK7IAIay6OQtDzh
EsKY15u02rtjms+Sn+MvAF7kKTM3PR8M2WnWrzpkiw8hRgKZqbBCWZ1WD2mhE5OOoHjD0lSWnrTb
CYztDqIuck+X+TWTGRqT3HTDtp1bixzxqdNuwOwnkDfy9p3Ucpq4MJ3T6jPxN/kuXfITgWThelvI
jR5Gi4kzlTTf8xsuwGSUvcOc96w1kb3VWUmBSYe3YLIRwzKKoZbDuTtDaK1UQs3vkV//oPgR3UCa
QzBV+SCvBty2hcSNy/xt4B6qmD48uQoyBotYIsSppsJLgMM6/bkS5BCYLun7rYDh/MbQanCyHT1r
4t7a7rcW/iZlmRuA1k6KvjSL0SNMvEZjAqz57sZhxWgNJAo2iDYb/qaRdmP6ofD3H10/jzMzHcQM
B0qLfCh6Qj1Wr1aOJUvfuMN5d64TwTvdvolnMmu/f/dQTfnIPC2tN30sn/HLPdGhggZVOJ2l5lfA
5/zXCPN/7esOfLsuQjpm9jHr/U45GOiHfP9B7Kq8KRy5ZGaaJF/XX8YWAUUS1z7dR0pqjCNY2vgo
1i2Jwi0Dj2Xqq7Vq/N3LS2/5owxuBvVvKs+nJQ+4/0n9nX9NKJ0fpPkeB62aV6MjLBcWDCpRWX9w
1U15/UKCmq8JR7wCTY5S0johw2Ura/Poor1+WRN8nX8U5e+9wH0QjGGZrSIgsEETVcCCUfSfPyHG
UWEFexG6FltVYyQ1EKCc/stFd5oQXy9astZ0yPDRt+Sp8L/NzPA7ys6zljLUKRqp5p/0c6IBax4N
pSjWqqSxbIHAQfBu0LJWZg7EfVdSlv9vhMy4z49UF33Qe9iv1Ad99nz3QNq9KxcGVfD9HN8/FzMs
UTcyZqEZYKchi8EhaZ1aLUZ2xruuwGcUrYSqJelvWDBhcvON8HS7g/HbVJJSsl3IP3VPu5OG/IuV
jzehElabYhP/LkUGw8THr3TxewWDSBoeqyy/8t0XIV7TlBNCVP40GVm7eQ4W7IkToclgDdD0kRvI
Y1kzXbBFK1tts1pEpZvJ5vXvGjbdRz5GV80HpzagaTrIzdDkp6Puaky3xr0d0k2iMRjMMWBxjH+I
wqTId1tWgbkwTkiJeD4xdcLWxbRZPQGktYYaOAjSB1OVUa1soCSCzWRwEKFHHmE6rvqaVLYl6kCt
TLGPiELaak6WvBHhywChwKEGtT1I9mXHEW/PUxwcs855qvw9xtIhVEN2XrgtMTY6l1SDR4hnyid8
mLxzhjr68E/NHJToQRJPKMNOvNIB1vmKz6Af0DRV1aI8ZCu+ysaEzNJfl3E8ZsoTpB97dis4Qqe/
szuyMgpRmSu5BSYBEpr9oTtlyvG7svDOL69HCLqbYke/Qiw7azqq6mY+78sGF6vcOIN9oRrTsT9N
1y/pKJQkB1OMk9woWkzIRPxuIKFOkK5CqaTIjgrhacH1wwzHN/GJ9RIBBij4nc8Oim1WkQ/pOnXB
0MzsvUl8ziQH0md+dr9JlmUWuTdnpMIy9neR6l9A/2uls+qaiSzwJh/DU8LUn/l8xp6qBh1RbSpt
AMu/GOYH3DrMUrMfL9sVeeBtp6AAKKV22d5Grue4bkcmQL6JOCXazEoeBH2s1OzLQVvu5DFcLpBd
6OlCcf1G4/3mvXwroESjE2RiXWL+ERPCQiPFRi3erAL4ypVagksG7Hmo+0DHNvLPJEPoZ9/kiMMP
qoPaPqlQatllyAFCDvTXC98CJHYT2J2CdYWE0gIrQFJUTnB9BsITxiwtiW+/lveRdUjddjY3Aisj
3iRXfHtsmLACkq/TSjg3UtRRCe9viVoAMLVdnm9cWshxoyYnCSB9XGIdj7fvSZMpYY+9479Vnrfv
iQ4rGn2//S6gx17vXz7ygjzzeedchocuAvgn8coJQY4dwH6bAIZgTX8A7b3t3YMPSxyA9sUTnc+W
Gn9MqX+/RUkTy3esT6Sd4oqkAKhlI0miZUvsOLiImhS+IfaMYesW2H2COn9H53j833uHGhr/8LH2
99tiaX1XVObIs5jZXR46u6qao/dFdD5QW1k/NEW1hYHi3NU1owv6/MVmzkFH798/+VGVQPhdcLv2
YFTbp1sVS/Ye17FSx4SjEOe5CSOSh/LT/WiIo/5aJzSMs4Hy5yS1XqSZc2ZEJHnTEr9fC0viNd8K
g7qscXodr47K5E50crKn3PTnmoPpSDR6nEjJuty6Kl5hj8RAGsG864jPDBu0AVqbWoPjmMSBKeyR
21vQC21Mx/FD8dvFQH483jlK9CyRfjYgV9g6c/ETFezDJ2vwHccnCclwO/LukRTpIZkNPjiwY/SJ
YrkTVltBXTnqoXwPyLI3/aliL2IiSFUjWKun6dM3kmcEVEt4ubI07d2yejWHNExE2kDCH+QGdvWA
phx8m2a0tqC4WOMsepXplkpZXVTo8OHwc4Jb66MZh5r2TM02AV9EZXn86Tv4PdXndEYCUsriVCFc
lPcJ29/A56s0tXtgjMnq54tvTwh6dTt2yK1HM4DIMwBCVa/i1jo1Mx/KhxZtduAaLOySvLq2WZO8
dXK7LfBipKnHeAWQjzjjCyoR2lrY3nspHR6kiSM1i47QOC/VdMoOLe93v4SoFDPXX+CQL6cCyih6
+kc+1E1MRBhXZKUP6tiyh8XE09BHpZVef1FJhMw1xchnxVfZKNCQmqvq7SHWlOTAeIMhSz9rYiuK
+aONg4x0t1dUsUWkZLbJZmgV+1wdGiphpB8wutLTK53J+4850T/EqH53qu5smL1rsIJkaTss/p2p
lJFNhkVQfqXrZ09bJ4+hGOobOpmP25Sv9Dj5xP8yLrg6qqZdrcHTe8NHWvlfoBZpznblORIGyGeA
RtwsItm0F7HqgF5hQRNSwmoRZ6vnymHL9Z2tSomNRHaqkX7BJKYrYtb5K99aXnvaYASXljNtfsfl
Tpk/bY+mjgksKYQsNZxTaKwNfyL2p9zT1m9hxNYlzNip5Pz71qMsV9uZzm98/jEzPwMcSdtzlJ+t
PAAUpG232c/X4kMddF38jvSQDVbFYq77roGTFcJ0QtsVVbAkZHKQhvS9t954ZlXA9l01KQVAcLcX
scGorWm7C/Ne3Hifia26mbHd3HYDgKCGoLT09vstf2Jdbss0I+d48mzW9w/m5xjQ4miSA2MPeT8C
8c6eUcp5XH94HKxdY59s21nBQlx27wbNLbGHEOJOgRIZ61IKYB6X0ePlZQnE2gH4GDUmza9y7bKE
OBhNvPc2iwRUuPPgQyzBK9EbXp057IUPNmKazFnemOgDsbDbLRjELt/fjB7IUYQ5MlfteFUp0l1N
8/4jtHzZAYhG52ro9Ox4K87ulGQJcO4Com7aJvRELH6l2Wm2dpVAF77oHDugN38j9uXd0ibEmxIV
+Y9KkQ3TNVR+8yyQl+1R1hTtaRVsiPCmxqCvIVrT7YgByzrqEkE9Kxp5Dg6vpKFd3Kj/7eTPnmes
KimiYjqrIFJ5rLupW0OOTz1JTIo2AeBtCTyzs+kbs0zm3nZ/f7PfzK6muKoBd6RQX93Xfe8TixlO
C/h7REwUendUx5ooMGaYOTebdnzlctCcTaaiLTB6X8Oz8Bz7UmAYrYQUu2arxtH/uViZ4bNYPciI
lSil7Zmsa7FGVlKFE+Rkpc0nEbuSQLfWMngz8HlP4N1XuVHk4oikMxZWcZst/sEQJdnd6wGvIXJF
73tr16H1geBAEW476xBZv8oWt2dSnhJDoBHyg39NVspgi7osegkQ2O/jjkYK6DcYjm0YJAtG3a2Q
YXenWOHc48V03pmkBUUi0UsAdfRILd+usNFtTWKOA+KGOeVwAQCU0bDPCJ1tzNEjPRj8bIZAkgSE
HZ4Olba+n49aewd/Wt18TY/Pg9n+w0CxKUdOEfGJZp9q18ui88dhPefG3nce4sQ3SWXSsNpTMEeW
3HCyTt2/pJlbLhSq7CCDqxNjbNgZuWfXmoBamBHesVLuY32vxMaLjOjtZZcTn2vqrpq6AGMGUiu9
Oag5evKc3aCbOOQyAVKqaBEIxepELPIx3oUNGHCzGm4bsZs/1lCOEA1Lv533vP+HCZBGcNdzrPA6
zEP4MOuX023hzKHNH2QG0EKaUNBqL1M1C8DPKX7Ta/kG+/WL90yrtlkkzMo7pWeqHXjTTq/g764W
KxdA/qC849AXiutmmLVBUuqgC8pbGBJeOZ4JlTTdxZ3Rn01VEK7HdgBuh6MLZOtHtjd9qlXR8fVm
MrLhfoj6V/9hjfkGxPPp1hZVjbpO4aCc5XAQPPSAQwJrSz7qc4SI++tAX6buQtlRS8enrG1CmwWe
BpurjgweA121UPG55aKr9ly+J4Ad6pJPFsJIr4ON7DuQXu+LniJ4OcztemnCKyDM5neH0Bp8RjkQ
bdO7raOCTuBzpfobQ2QtTZmsYuSHjKpxR52ClWmAC9Ay/+bmao0b/N+h6adeKK2BzhTLfys0ss52
GzQKli9wGIbbAusuwJf5Bp4jH3RbWDJWD+KhLUVzu9yOvJyPv1dj3Acmzp4DpYUnOjVfQxAz9Muy
0aDvkyAZBWwYL2O4yo9+Yfty8aubc+5trWKiGk4t03ihhjk0tqL3OeOuhhrxKTJhV7v8EDZgtGbB
B7ZYw8Xp8seRlS0p9I2sd6YssTyUg3b5+fl8Y6xQEhvOpSOPSQdwgAEndwrEPID1GHS7CNn0RSOF
f/qoriiEk99wISw4EnSTNl8CshR6MhbGCmY4Cn3i2cyoCPgQPrs1Zc4NwV8oVO7jshx0i5IxqOeX
7GDGYFr2HNg2dilo6bkP6jMLetel1fhIjI7NvhF91J6nlJZIy+P9VZgMWGfyuYetgYOGeJWzTfsx
DqRHJACXgAfFlLi3gW2hszymUsC/cMeqeg07SHIHqcAxAFvX7DjJZcW60JJfYZwiNpohTqZqw0dF
XLODtlk6/6EXl6KIHnfPmpExxk+QY8RsWejQrkrDKnwBzhuWHkyJ7SgvLjM7uGhDK8T5S5NyD1zg
m5hmcGGwCYm/NV6GvjL37pi5vP3OiyoRy0CKECeB3pS0jEfwxtnlQwvRa6AMVrJ6KJVibOllm605
9TzSU08TxuvhTQDQaPUZnC1BiYY2KKAjTJsyBHLOmEl5sjoDMC4ypD23MtfKZ1cG6AYp1Vac42b5
CXG9+IagMMdjQ+y0mC+Hbi5rYLIk0o7Nr+o6Q+zL6xDfPdvMGF3NTM9488Zdz4qF+jtvdQERhlD+
v8/+qK+Jajw/tgmfEiElHEQitsSL43h+jgABcbLX3b7gaQTm+hULSkVGRRfH8FC0JVRNvpYuTsNr
YEE/ULHD+opqcxoyxBGBJcZdIYMMlTGhLwSWHQsSiRIyMYKVm8tCKxiOJ2fCOu0IWjy9yiIVfUfq
pLM0QtYbue+0OQW5ZIWon2phNG6NhwbGZG0aDVweAG1drt18vl8tI6ItZmEHVConYRmCO4RCUii+
EOTNaMifsJVvaC/B7ANbolRvJL23xsjyIiRCDoxn3u29d8ewHhB50AB/bvaWFVBB6tHT2k0f8Wqp
RzmAj8wdFZ/xJ4RKZ93Px1w1J8FIfzM+rk/NkQ0bH0vxFZfdDH5AFWtIZHlEVMmawqJ4D9gzGa77
dMLVLjpIgAjPFeRGV8uQHQ/iAIVEfgnDwAnaVUn7ewDwVMCUIR/V3YQCu39c+35oaRTZ8lTcslD2
PMU+P0OPvz/D37i6fNSi4Ee6+idaF4cXVAqTJDgHIQBXLx+dDX8dUOzx0Bla5TYrKxGIctns4FXZ
0wBInBBVM1LGPkZd9hJEVXYfjc3Lvcv5bzJY7n81g1PVja+/2VdzB3i39b0N1ZNATpgs7lVcs0xz
QveB9BB6OpFoCsOUOGDxx6HFtw4wibtZFtsHHp537QWsnSgJRVhLsv8YoNjEwOmm5/MVAqWWwVBU
i9R24wtzc7sCyhrD7Bu6lvaOrJiIMRfLh9NSJc4HV8DIICPtGkAf8TTPRqevUGKYkEJnex+gDl8w
TzFphVcXaEB16y9R6LzQZmnhd4usI0HDFe7Gi/jKmn2n37LhfyFWz9E/qVAtaDAeRAIAKC5D4J4a
tDi/qfgu8LXYWvQgxuI1gfg/dicckETFWe2rytTf9lUD2XzoZ0vEy7cqLqMKeZjlr0rwopUsC0F9
GYNoKmTF/3A1JV6a2wb9nOjoRYCG8tewSO/v9unzE5cvt+EIBC39fPt8TL31kemwOnjHBPC6B6Zl
6GqO88Onv10gLzTsi5CgAt8Lfef38vMVlld9yv6WN00SgGoDFh1tV/5gwq+IiUem/8N+e1JabIQ/
zoUvN5L+ZdiGEHru7tTnHNY+VKkOLgEeXmNjcDhsrKDqc0b5G+FWpAeoLet5kM8kIWolb9mqk/+4
gW+1FcFxxmSoMVTzFC7QPmf3/FrZ4vin2j4EFb2u1EV8BZ9D6vFBmAFx6ayxFcebqgzAOJl2GS4q
fhZkO4qYCIeU//QxyyjnOTKF3X/RMX5Nsz6MoRXW7hnhb7sKKXSxBEfdcqapixHQ7opLZl9nXGHy
U1MPuX2k2YBKXOkTRbgLH7h1pEfOUzYlR9m7U+m6fN43QTYyIHgJmqulSrToKro3RZIdAGI+kOgK
UUWMr2XEpZuLN7APYt9DVhf/MNBEk9OPf6X9Fgst6+SmcS1WNKSCRx6h04Atoo50XKAb9khEkDCx
sM2L/apIxEy0nxi/RDOnkmi7859z/o3KbpIZrk3dH/fDzD/kgnuOkYb3ULBqWVXBfbQB3TRIBeIe
8nTMgFGfCb2tPWZhKjY7/9wWTh/BCMVzgT+CAu2G4SW01jbkZ5RhDkzXUZJ0LFBfHWH5qoZrGOr5
sTcLsifHCmqlA/iUFw03/+XVdTUNevdxAaVWKg1SXFOm6Jj92KoSALGUQNb1AY2yv3tt+yiAk8Ey
Yu9clrP7WCJZrLByHahniK/JY6hHNUeaC0Cdxr1VeWJfUjAeROrtmumf3MnuMP/xWMAqZF4UlrA9
NFW0WFaIFuFQBzimhLc3xF4m70PfO0PZfjVwduGnN1KGBs+bsticG1P7lWmtabZSc4wlb69DCWy0
H/Q2mu7VFeEGlWUgFxGcKUu7jFbTvTXuFVPBern7dUWCqIm9J6WZkmBdNZNlb7JsrlrJRdEUUukY
xXHHJ7JZX6NIA8EL3ZKLdyp2RUblHGFC91TgXQw2gsCYxkhQH99VO4UaPCqsR6NPDjQbMiJnSabZ
XCL7FD/tjhS6UMGMo/vAlElbMNLnftRLYTh9z+KHM8EJcMVIqNVZXEo5LEegzhEriQsNruUPZu5Y
7h340mNkPbm4tyA0J7jz+dzv3tPbvmAdE2trAQjcnFeC7aZWP7TunPy/vsOR+dP0rXjB1urRjKxf
vGDhMB3Fn5ZxDAQDT+gYO8P0GO8SgR+h62Xl2OTot1KGy/tYWnjQI9hTyGhBvMtuBCkBa6jvTOkx
3046gF8anrSdrs9lQZ+uLKYXnpOzEuAbXxvK1LPucAxpI7pzkwGbH05DpZ7bqqOhLQLP/63NkuHc
/sbgcft7trpzuhOl6RLpdxBLjThMgu3xvXfIxJBrGuSt4M3AdNad42uqQgOZ5NPcKXrUvQsFp+Co
DQ8ojt4h2qKF010vu+IQq5BoGDyW+EJuTq1pzIzSEa6ohieW0n/9lkVcK9RQ52B53dWsdVutEIzp
Nk7H3HUzzs7h3lvHb2VvRKtS3veOPeOIJfVMolJYbUyD/2Szxtj0BBMRYds9T2B18DPkyasbsWQm
HHyiCLrrNWUJ57NXNNACo18LhEONlcg0eIhF1xZS15JZiqAh1bE7tuzAhJjHcGyiK/LHnFxaxRBF
pOdmkf1VJUDDTV0S1iWkoeW785ak412lojVm/V3qHUHgu79dyZk4KeE8oO5LVeI8+jcnhHsrChkg
FMYCcslL2rogGBDlQMw3zlDq7Dr9BDXWKrh8/E2D6zmhs91HK6YJUmg+yiLfBX/YtalhplFL0PBb
hDxMw77L9llchoaYx7PbvVxIMxMx/7rx2+IqJ+GD90ZjJh2dkVR5P7XplqtA5hk1Mhkli5Hf2vmV
yJHNP2vmzIN8f/PSg0fQMSSNb0y+tDGyddofPv2+6pljStyCnKF3QmJGsC3DWaDejKoK+ZO3z1DO
lemJiec2JTEb430AI+k0Ajyy83TglQI351eDBUIDTITZ/6+Qhbq9q+mEMsly48CDxOAkplk5T+ok
G7nUCA+/3QMI8G4T7K9f0TswGVdSeIoHNv5fLCkTNYWtQ6ergq8D9p8mf/OWWg2hTpEmORXSpo62
cfOTU8OiieVi9fDUCE3mxm9VTtSNYFXT4BQFaSxA7gFp76DDpTeUpImmd1dp1i/wDw+N+CVtF9yA
QrjZDZPWb+btmp6XuaDnDtiUHcm1CFDIosXpjgdV5Meh6kdI44ghA9CkyIZQS1yQgneOGMGIlOFn
FVUPwIQiWLMZBEMEM3533oTuHVh7d5FAPGd3APjxI5xiKd24sbWDXabY1dqDsF9fddWpF/yNG7ny
N7iMV8yqlycgiDg5P7gZsrj+4q0nTm9tvX9QejrCf4MZs330SLM0dPuVnKmEksBJ0e38+w9DKctf
fzXdupbC76mdxP11F0gNUvObuw1c/m4MiSBEC1vVwJ2647Sw4gvPS9UTgKEn/oEStHkJvvptiSB7
3qly83i4nKMpisAs8K4lFByz6SVU6y3BFcv1BSxoT/o2Xc5kvmh5tFFooUSo4aotVi+tpmON2d71
zeHVLMhkxJ5y13sK097/fVgQbhbCewO5f5alvKAFAK7RgKhiErqCU3TyvAl4v266Nf5Y77FM/3Ow
M5+L8z90W6HASscfYJOe5LBBP+4qMhmnJ6NrVzfT0wjUkw53QS8swJo5iOztOsfs5htZcugCDmrO
ku+VxfT8oJaE4iFzOUb0X5UtJVoUWoPPMIXOTkefK8Kr/dwaducwSIvLrK8WcUJku+CPQPQCyonq
rRHVnwBBDXnJ3DUjEG5UrHUG7qpK4GiFquvnTv8sI6BBttMORXif8oOOqdEA6htaAuflFYe0etMf
WBtDeBF+vBoSbHcHGODia33mA3Ape/sdQ4M4Bl10XBBMylel/BKNN2VPseLVMRqiZCMkit/IGwik
3eWlO+9Jj2uVwAGjZEbHA4aC5Lhizc8PImPGwFVnkZ3ED2bDzhROK9P5xp9PWtRD/z0y7FwfBBCo
JzLc6DZVL0rEk8n3CssP7cEhacTt33JZ8mHErQB6L1DckNCAP6ZLPFSCZyIc3TWx218Ljk4uN9y6
DwB8NtHeinurwcCK+eKeu+FzYp6dhamFBlDuuBoLhxVGqJAjZuIB2gmqnHT+KijYEJPsgl1cmdx8
q6NGmt1lAHhlchNurZVWnrjaWE31OARkG7Ohvo08n2eajd9lV20vLS9aVHLRdmgOKZz4bAhJgZR2
eGRcjQg7BwKiHKfatvjfJ7oYLYupGAvZkgoapSLZ37Lm+rei8/JAsbbyl8BERRPtB5qrODlFU8pF
z9qN83rLZ2VL0ShoksanrL16mIRtKVTq16S+0ziJhMcFbeuC4NWXY4sdyZaCVKhzI6SENXRu0LYi
A5Rq1PO3vGkiqPKuAyW5ZMOBfQyIQoMaiAApUm4icbhSmA6HSx2PclR3mB2NOVxk+cOphzjdy/Zr
K1o1sewzPDgwzvK75V7v0LVXwSUE3M/O5HpquJof+rI3YqIrpFTkr9pTjOar/tjyZS6vgT7BAkhG
g62iUW5JYIjGcd/j7nUn8kgu458fV01U3BPZqXfLyZ2ZRjMkW11XLEyG2kPUk7Xx3m6JDH/c+yg5
AKjvF8Opbw57ru5Zfo7GTq12CM7cD85+8Av/TKF4ByoN8L4S95nPlsS7oaMeSFK/JWec5dJOEA5t
ky8AOoPMFd1NTDfgLQeWFEafaudGyCz5PPUgBugSFpbhyEt5AiwEkD78uSnXlYDUFvSxymd4haOB
OHymYCWx56eDQ/YI/Xz3SBNVBuNZQZDsa1siPRZjrIEz9Fd/CdIw23ZmfFFJdhfMQA/pUNxSHlQ0
hTvuouSVIeQZVsiSzK3M+evqJJp9nhvzbgcsUa3iwBdC1mfSG+nXUF2iw1ydC7TN9E+8olhhv/L0
uzQPU8+fkJs9XVdah7or6A1HQpg1u2tYHqZKfq69tFtn/xZEskENsAEf2pbqwP2nVujv1Qd+b6hY
F63Aqv/VMgcCxGCNfQC0I57oXUl0UlXjIPq5AgNVteWlX7UkGX01GY8XbVHzeCjie0a9tWmcpT8y
VUKfxlMCULXBzVUvuviLN6QjDxMiLl5zHXUV1jh75n96Czmq5jAPmq81THGG+906p5oDwse9wuL4
pkznXKouzM+iQWHUqX1b+WAKzy31z1p2F6b0/8PqDT8uhbNwn8ANgnyjLgG+9PoYBkkZHI0TlSaF
QiaxytJ+awYUxgVaD8yd1cOSOm2qPwIdPX5TavI9zQaN2Di5gAJoqEJx7z2m+ao76eu9PgbtPR/Y
h9tmcVl5ZqAqoJHC/efvx7o/CtCUd4uGj+OoeR6F1vtIDTwOmMsvyHPt2PF6cZy5B/mTg5Ii7JyI
VqXobglugqZDEz1FVGdOeoOIQAjGlWatbKuk/Hr0qXEFbgaVW+ND2CB4jAQKkwI/IjaUkv0rM72j
WoEDqAYhr/8euNRZsSDEx4LNfON4OL8XQfq8IYYIHhnjNBG2YqSmxk4CZmh1cy2K5DuyjJqNaaa1
DTdaFRpeKJfLcziiyU8RJyL304EriEl8Xq+4pJpRupVGihm/tBMKhvBjCD+xXOL9o872lUyppBHe
XCRJJMKZnNQW8+jkp2tdnvB8uZF2Q/YkD1A5GXRqHWaV85pJALTEK9rwjkyMT979GK2Qk5sJc96i
RjgxsTzxgtcjIELvP+dSTAHzNtk0OcuW0X78r5diu2xe9y1azOTdXMiTuDBF+T+wkwfwBAwhpTgs
p02INOfzMfu20R3BkmHI9X26PeykgY1of3g0yLPtGw8dHu0ZrgcA9NSNSwoGDq7gesNX03XBmMvB
7K0TERoj4rpSFHCGbV9KIFhSLbccPY9EQ931cDIZeH7A1KNvk9BNWb60xwQNiPBXraYen7m3eLNU
P9M6AVAoCbDmO7LsqqYA+sU1tuPIKGnfvSmOgLyBjRPRyIVPKz7xqa7ZQDHaUhanuhMYFAs4klr0
jhf//mdHDIN1LUWyEguop6UMoNuq9JEs8KmmdvHWxoRMvJN3jPZDJ2ZPdzKtrxwYkp4eqC5kTqKn
UxVJTSa/KxAUkcFQE27O2XpmMGJXSAE4eGSWup9+1B3JYBdqzwYqIT0rx3EMxtvNw4nM5UJE/u3b
EXDnsU+/pnditwP/981+oggiFeiEDTv9ehJc3DG8F1rTf2qJ3kr7FW3zf42iClogJ24zcXExI9mI
8X5G7KagNq2I/JtM5+UsfZrjHy/Piy+VCmYRhzm8ylkht434E5ax0nWHKjTi6aeKAe5k4zr8gi1h
UoS0+kHccfi+0sp/SLibQItW2KyBwzVq2+0IESV4KYDcCgPdK5EGW86eos/fIdVh7Yn9JX/MOZ+n
lgs7+qa74mI56XEdRh2rZ/UOq7xi9FYZmrym5ktRi5Ftxa9F9VnRR3JH+YhwX9uw2+i+k3xFOZFj
u0aKijg3NjcHXE3l4Ffhbnen5kUua93BnFNxbjHtqNp5z5LPTyTUeSVY4DbdoYcE3Jwk1/Iy4O6c
90I1Bl3wWuQqI8pDGee3oED9Lz7e1O2GXPalJKoXno6T6VtXYJ+WPdUTGEdoV1rx9gyhCQWWW3vi
1RwsgmE2k2O6+7T+iAZrKpeMv0qVKYilaIZlMIjjCgbJuXEx1oHHaoHvpShzCS32c6vbgRHjWdzl
khP2ZPJFfWf+pz8scq1IzOp/kko+ihgr1WK9Yr9HxP1OtRdLx9A7eB5JcBhNz1TmsC7PXmLVIxjJ
PpDw7zdMMirTHK28j66cQJne8MXFOMR7Pre2HvdTWsBMM4weSmM5WHxos5AO/ABREbyOIzk7GEly
B/jGfqpSw/i6ekV/F7A26DQ5lWhLRbXvUjGMONIZkRClTpdK38YE9XfYLaIPbxZAs59sd8cdIogk
Zt6Npl1jgituI8dUnSboQzGbsimV8ElLTiWAzp33Tm3sn0uIaqRQTCfOIeYzdhn+tMYfNfsS3+T/
hbiSwU3lIUQ1cX33GNPH//kisgoPzPkNWitM2mawH8FuX7XNpfE7iWSsZuT1M0eIIOQCXXC/X0gL
mfgy8uVmjteUupBlrHxO/uGFRMbH+1Ppcl1vG+jqLQZvo/JS6UTHYzLU49a9Np3kNFV1Ii6KIwBN
UCGIMx+xU53adJBcdVYSKW2JG/jNaKr5rrtmdfSTVJmdpcTSS6xVJqSNx6KnhXQoJmI9Abn+dPmP
8C3uAHcs+nHZmQJeINjDaYkF80WtrGSO5fUnhyGjeFFWQyYi7FC7IuHF8VorkHD2qBRLg9UpzKeL
wN8r4t2cDzYIyoCLrPi2mwMXHebCM+mkH61ksDgvT3APFF/ECmR+F4KgG6dq5t7WbLs1IwH653I0
e1WyaTx4SQx84AQwwz4pTTICH6B4KD8rhcMrEgSEfq1tYyLsS6KikgDLOUSElzZq6vjCasfKP5qs
TKGkeXT2fxNr6gd/BNtbs0JFyVRzuz3hNUhCH81lRhnDs17v30ebQSNcx0Gnoe9+mlow6TOD9Vyu
cviN3cqZCU8H32U//MYXxTHA0OOAJSIiNCoabZiUP8123TFafG1Oj8YONZkjEMyWtKtagTppmoHb
FzY4mCRE56Rvzr/ZfToZrdNdbxXAt7gqiK7uzJe6/l/hoJHYqA57hp5koJ/HC+FCuBxXhHCvrhMu
EgvRuqm9xG7okIUN0Zh/J61TCd3bmvipB8Mce63kcGEgYDacn6EDpRmI66ruGKxTOTGYxGLKaHOP
4KzGGDY2vYyxSeF4AFNwS1eaB2IT0UoHuq9U6iFJDOqUzz0YShgcN5eR75Zz1x2TQS9J7Vfv/0CI
fx7Q1WjqPvvj9mn9JVXUd4li5JTtrcpUK5P75yoZCvi2gNSAt9Xukg/qLc5dZSj3IXCcA12vSfOx
JvIQ7ZIx2sL9u4VdkBOj8LLftXaz3viYFAmMcf2PZgiQbJVxJss7XcRfQpxAfVUYrUTm/Ps36ish
lz3FbcNk7qWGhJhXK34Tfj3e0SByn6hOZdYcq2CpcW2HNumwcKkK5UxfoyZ6FQz8hmfEbBWxDqg7
d3F6bLFEHGTOiZ+tkT2/Al2F/R+K6h4iZxSC8wc4i9NLH2ycFEkQKD7fCsZ/aVwKFwCGq7tS3GQ5
/hvXcfhP9GIHaTXNzMn10Zo0JGU2rOHgiinP7lhJjW/oZECf5ecpf2F6/d2DtbmJHoO23sbpDxHI
YCqshK0jxWgwEIi7phyIWq/wx3E0GJ4agRqJ3sdLBm6XNxryX3PEjfJ1kw7rLVH77th88++Wizoo
Lqu8n9L3vCrTPm5gqZWSDDgS55pd0gK+LqeZmahY4RaclQNzs1DZjcSCAvfdrX2pHxEhJnIjdg3j
s4gycps/un6gI075U7NQmVVb0kU47iAGuMQ2w2GbWrT+E3kx0A6vaSUcRChU+LbiUfLDLzzqedMt
Heu9IaxqE8T1+IlUchad+zdA5jQQ1quHDqOKC46g1qGUcMc94b4rpbmJ86X8/fOlwktOu1OLkXVY
1Kf916Ky/BlAvmCznLmP9DAAtevG7Pazj2vHFOUHMt1g8FNqbZWRNf2ioYZwOGXQSiCy/5bhL390
1RrS4VLwl5tDwkM0Iwd/CH0EUqfcHoR+aUvRmJQuCWhwx9PFnptMXZySypwAO1TTbvdctrHj74Sl
1ATgR1jX1zBOdx6ESk5/7n3/7E5aIetdz118BhtZF+wlDIu1y0wF9VRRjU//KgdaJLWl0vRZVyVE
+0LYUpy3Hqkh4RnEQLdt2Aa0xG3RBOv/lMMcb6MQZZEvHGcOzuZueAA1SXqZb+cxSG3b44XTQv5Z
yi9a8CaH8Wqp9/6/n2K2PeZM8T6QpDxFxtv8rpU+wtxpqOYdMY0t+lYkRv3+jnRDiN/nZuBu0ZiB
XBEfMBUwGmKKL5qmMnP/fuWLDGL4ks6QRZebLjQZe//0qyuAA1HvFEPRMvCzInIduAOeP97XjsAU
TYg7c0Up5ADC+AYRRcu40om1KQwR/FRlsgpHv/MebuTB5BXbIh5twE8Ju0t4Yf5smYbug5hIv9/u
LTKiKLlIyunVgy147MFdj0mlE8M6i9FNySIX9/aAwpmbQbLvkZlJu3+gV20SiNrfoIM3D8Vl8T6d
ej8lbx8Su29wrooIZEWufjdsAnPrEUmZl9s58G/nIzW4DOnVQnKctIAH/+zEKZTK41+65YT6c+bi
obO1YdwM9Jfnvi2q1MiB/pTMP4wgf6uOTyDVA3+N9yqjYagDywrVB2rF1kz+IxM7D7EagCqR/29L
6UL2WevxwY80ztBOZr9hBVHc5vwmtc8hE2o+xVNVequ6IVBXHWdVGAgBNhu5f/KCFbkqMOkLo/4P
uBsELVXLY3J5v+477zgKabLK7abCVIc/yOi8Ap4qfoNxqzSJcrhHh2KUOAlSxP5wiqWZ16OJVvk5
2UAUbHYo++OYDQkMdkDHFulr+AWhzxBQVUFIQ1MWAtOAuCr3StmF6nMophMUAZBzDAUNaHuIaOpL
ZbDvLHotehFC1r+OG3s7Hu0NhF+0AsSaPeRWtO06S8Ikvney2oCBwnwGpazb94fbu3s7J+PtZNNg
5KdvGSTqkHUXymx+mqwMQBrsaSoEIgPoXgfCPdNHkYp0l5RCZphDWEVf6tRF/TJEYEL4y2dndHBW
oiQIhmoJ7vumkXl0ocyJu+VcfiAZdCXvpOFm8WOzHKUc/HbQsJkCnvpo8FrP30LlRyXvU2QwQG4b
bS89nYRI7I8nsuLMgO/HGKHzNFO8NauE+R2EAJQ0ctmdnlgzxXZ+98gl+1LD+W2Wexsjs/Prva0j
Y9ALBiqyVGGGi7tZ7ntC6yZr4IRR9Gg1+rAF3m1WRTxb5wPNt7NBBXJ1/HPdOmZobaf+wWVA6pXm
f0NJKAseiNp/fLfBNxNZj1FSj88onOIoZDL1QZ59OK/GLJDxIzOqOoo+nrShHSUWTQBwSivjrzYd
alpZagyzc+zu+PsAuMBv/IbSRHaPW+pE1sPT2jGVIycATV4r5C0pq+DJzlx76owgzT2Y92CP1hzo
r39MrhIllwCRbSAVJsdp6QCFJoYbQRvVFOBWu5MfZz/DcPaQE9lp6qdWe3mr1JLQnpDunNrtZ0yN
CbK0vBZq8LZWwRmqzoSx2iHXEp/ovVD1mzgjByF4yzOkCYdH3/BztWq14zf1YWHr25+vAIjcYe/+
D/mKBgLO1icJzgXQNnyprcKzgpm8h9+QdcPa/QNKrZwl00RoAH/uTvRvZBtmR2aqWj0w9nRs19lk
+/ODbPK/gBZjLPvQ7ZfLpml1qM+ee5JPnTYGgbnFcTQ+KS/GPJZkeBXXQ8Foo1JJoHJxfeBRInkJ
gy48stgtDgKbfFoiQXjyzkSGz4+FWEOuF4O+bXeQ5ANPgZrZT39I40IB1rxEOkuJU9Zcm0vh8cbd
BktO/f3JxDjipvXbIzrTJvMsO4wGKMk3grFJCj7dJfYcIeM+ggovVV6+ebupcQugmc1S417r+eap
ZuKJOGIvvHBf+fAUupk7FVgQmkKkk8oJirfcckNIVPDl4lK3gvcR1kWRiogn9zZ4laW0MmOCivGd
3VXGEicFx6b4xwtTORue6gfdfVig9EKnY+zw7RORu64nXU7Lct+iYsk9I+N/TkQvvLCxpf6HlKdb
/r38B4b7WFN2BfBot9s5smziO010xL2V0B4ymH7eqIiFGO6hG2f5K2i2cW+NVeLRXeIx6wda7QU+
pMOYtA0VXLhS5bJkNP0aOX5uSipE8JVoxsaYdCk057sFBE0TmnXEb24C6cdd7njt08ucmw/+AQGm
MPnRUdZKW/aZkUO5YdgdsgiceMzI1huNn0aNMfqPutS+e0+K0sXZNSAiT0rslkc7rztSnnPoC1pq
DjijFUbcCILBnm9WYFxBSjlaQwajTjmCkF642RCXEP3ZEUUFjvHAGM/VzsOZ2MXdf/AY5q3i0xJl
QgTyAEVfZSTPF9EFC6Uwm83qCF0Ygag0PtuwEobWgds+RsheXt08FLj1IWmVYRuIinx6k8JCZk/P
sUzIwvAd61qeh7mWcDLePIITq8xNMp8p/XVIEQG24wZFcsU8SfDATu8qjYff49K26/aRiSfcd8eY
wmeUJ+v9FPVVivvx7liJK2Zlqnrqgyeu9MpWfVGxagWYawTDpdnpTvQKuOlYLczZ8hZ2EAm2bmaz
El0e8xTw8Fhyexenwwas40jm07hFesX4wBNOatslmGZgp/lpTDK/+3JoJzqtVIXfmPZkm47CfnMa
3PEtK3m9BULo0XqYCLd/iPceBbAdlnIfhZLfdrz9AAvipaysPQbZmxuhs1R2YgWlFA4csptPSe8w
y/M5/fkwtUwXf+onGX8xo9nbGfs9FZYND9JTRZ+5WsuSkCSlccxanwpTbOW8PaKf6zIxKmfHfRlC
FV63hdwCoPkR3nm6ule37+S63uC7ymWuxJF/+RITkq8IDURT33igrCZRYSjKcVow0faOgxstCyGa
CFTpoueZYZSAFVxSDBAIkbPhM7QQxKX5qPo3b2Nr1jFagmBK6U36BvYyd/ML3JcbhL+4UE96VsBl
6FfdQQPnryJx2xrF5RlTMttPx2dISK1iNsIJNo7MiBWZo0SPuQfxsi037AvfuLVRZGC99ykWf3vF
lKfVzCJ0Czy1f98oa1vPr5joOZLh4eyAEK9iDW/5APwmqAmFqJ/FcIQlIVjdXq1KIHDw9bOgcLXC
kw1yXJdaI1UwPJaLrQnKRA82Jva1e5u+uXgfbq/22vVX/yOtMYTjUkR92DQNhcc57Lbn8e4CPN7S
d+rBMH6PJA9uz3k2hPgmDLUeNa88vLYqdfxWn0xdIODB9rx/yvoqet4lgAIcrVpxY31ccRuJUoHy
dCrDZIaDBimoRyIPCEp+yQTHkpkHGViSbdrrmo7SQpiL9dFm1qzzvWwJRZCoxBjthbGVZcn/badO
dsO7ksxbwEq7FSu/PjM0y0HbkSnykd7QTEvbhsG/RpUbqnSycOA6tXJz/+Xn9sHTL7NzSkm7QDT+
C3ISDfq1VRqdrwkd9P1A3LPfmzj2X0Awj7jKrTpzZfFMAIltb18KvJFo9a++ciVdIGGVfvYEyrMw
RYp867U2oUo5G6x1X02SezcUzZzo6NkAZrnJs30LS4X+bwPTeuCJUCr64ymjSKDzBmCF39bZsOWh
R9nWARgYcnImJGfB/puO7toC++1/RBtkqU6P56ewTOjFjLUf9VbY8l2UH0pav9u28+PyFTaKw0XV
4EEiA5e1l4dM3PWwg2Qdy0BCTYobWF7qhTNAxMnPAx/oBMIQdgqaRMfMdpiBsTr4e4oDtjWxugd6
wbKM9JzvPuzryq5/yNC+qopHTgoPTQc1niHwdakqZ2OmPFKXNjHuavVfhJZ9yWXQ3/JVd8K8G+mD
er/e0Sh7gi2ozlVwvsk2DMHUZSQNBZIks/fAW1dKxAjiOjo/jJK/qwZolG6PwZUMl6+4SB6cvSxi
Z5zGSVunQ8znheuBSQGgFrGbIeaghube3pYm55McbBHk5OS9BJKwvxeVx0vWYvZkwAJnKNPhucMK
0o/+RRPcsboS9vCBvDydrYci7uwjyWcqgk9oD+mbeWYixgA+Z2sThox9yw3kOSWlEKJ7t4VfHQSM
gEVaVowwqC7iuDS4c6kCLI3a9QnOxDUB/tVcd5xzj7bVuCPisUIz7N/fePTrmNEn1IqUcpqdVB3d
3Mxwck6FVraDWv98wVwmp+io1R9ZPDMhJTC9x1TRYumoPKcW0EFUiidEL2JhVt4pQGU347ubawKE
YRyUQeVVuhkHsQBzHWtir9jxmD2PhqkCjMUjOYX5LHOFyy+w+EC/plMPZ/Grm/mSG0+vR4DoxW2o
ikTozRN/CC71eZxaG2brJBpXglXTvLyRETfn/R8UHCnHIIv4vpQqByQNL8nm/aG4gVHygRV7JWh7
9YqGK3FsEnAxrBSkLIvVIZFHuq+mDmYM1Jqo2WpEQzn247Msci3rK9Fn24V6evP2FBLd7ptal/+Y
dE7fS+e/fqMv2kIVyGuFsqiNIIAir3teB6TXIqNeYEkDLZVpvR0X90PaB8p3I9LNssFKVzbefAyO
vNC/DkJPgHJcXWWdi+B/qGbXVDnxeqVVa5gZngZeqZ/rswPD9JekGnAbS/fFVhaANeDAO3uqvfEM
+jh10rL//y185w6BmaAZWaV5Ho/oSgC3FtORz8yJ4iouIyvn5ByOuiEenDvTIoNKIJudg1cZEriH
C9Zi5eqgfuPt0bWX4nMSodv6A8XUwxQJ1/RillGxVvdF/F6jXoh7T2ZPsCXk91PBcoALqw4ROtBo
pcvQers3gxVwc+JzujI4JlpepmoIdxqN1e+ZRtrxUhYYhMhloN+F/KV+LTXpKw86xWwaJIfQE5lp
hgfetFxBS4YpkvZurvFz0nkR8k2j3Qxx34Sei7INhplp+gVb99Pk0HTl7rlFNXtmsjJMf3LLCN7S
18keJmIhVhpCXsB2SutoVA1dtMAKtAFB2K90sY6GR2P4lHnlwBrqygEfyx/WGDUrSJ7t3Hc3cMAt
h7Rv3obPU9odkNx1FWIHowxCT6Zov8bCdBbZskKbmgNY2fOq5Yg1emEI3VJVRRavXaY716sMRyf+
aPU/pzDKHW62bWUMowSAXJkungTHG2K17nqFyzr01d71Fo/0Nb03MCf1n/WsERvyvxp4anLCpXrA
OJDW6ZrvA+kwoHgjkQWGaEbqFyyfubQETSzztd9qPgK++SxA1mnGLDUT56V70iPLNGFheUQFb2ua
cG1wmTi9eWKhlc46RydQqKsTFuBuYjKdjWTIdoij+Q/kgcI5UMR3i1iXzN5gRkQ4sSbXrjf7PZk8
Az/hsvOWWup/U+v6uSXkbb2+oFwAVufqqUA3cKBNy4eqq+jHnJWt0q2qCnvvMO263b1gaLWexj8I
StURrizjnPGNdeAI2N3sbPp8BXYekTjPj3S3Gzo19gglwHBdYqf32ygHYRA5SBmX/2qTuYI3e9iW
4Yv4Ir89/xEdvGOzLFLg5evHyOhpCv0uUOYdl5j2i2tnEzQeKfoNTc/NOvaYEjcMD7Aq58Y/qOZe
Nc9pitUyKU0M7GccTGarnWR3Yu6VmM1JvavY7xfVfrpftc5RQ9FuRSdD2BBsGprKeANERnhFL5Pl
54fAVbe0f7zOyc+EmvadpPyhy9RBCsqOgZKPihxDJesGHFxbOV4gOUIbbaWBqsgNV/zshCx7P1wq
LSjVtMaOmolJxmyWew85g8yPRqdrv3ZFykumH1MljwWp3z4h6mXAMaYPtmDCcAI6i3sgju/EDAsc
R045bmKWyWa4Zd7rCCpYftcbiv3t/KnuWWa5tIVIVs+9wexDiZLBArl3mPQj+b3slHb+RixPgKWw
Ih0V7RiVLaNPbEHGnFBPAuh5EDPmQ3YQqqt0zX9UU12dZPHEyd7z0DBZBcwe5x6LL2lTdZ4MWaPC
FPvBxCssnNruHrbt8OtdZvauVAf+Genvo9tW5B94+KvHLR2uBFWR19YwtXYODuvPuIypy8OXg8C0
h2roC5w77WqoMd+p5fa176Kattb5eaC/sWIXyXJVRM+uCtGxMwcmTg5dlWh+pHm3qbBL/9WNwAty
CjdfR/iV3NONiQVforQav2NYSqjPCGo+Ct1yrDOJ2GwNBYScdPWLyIDCWY8Et2Plm9RqBObsk026
6arqTZdie+F0YhsYsPUpkEH/jWXfhBvUYOl7iPOIM/5QfwhwMeQbxGz8zMpGbNCdTJKqFfZh5EPR
uRANb1E1qAwytjrEgTJRG7x6tX3yL//6uhGd3KXBmV3bXj9RQjJOQ81EUKAzfTPQRXLqlWVzG6LO
vbeZaU23tWaZ5WHN0SQnyQVSh183fJ2PuOkQ6RA9zJTcD4d+JKVRNgcw6t0HvB407mSArpjoeXkK
t/om5wq3+jxCffAZP94OE1GCOfK9plgGEKtYProS1OdplU5czi2nYleDJ59654fhuEz2dxrCIPPF
/I8+FGNx+0EayiYvSnqN7v9dJ+RwfbQVX40d3DVPeduWw85ADuBqxP/4hWkxpi7nxH6haFr37j8k
eNdlpq13y21j46YAeTDzwnM+knlI0OigZbJcnn+sqE15HyLpA/yYA/razt2pnKo0b9QQfDNtaHnm
0HENIM3QGZclnmqiqzMnQOcSywEWvFCgZeA1oHp2hfPWLFL9dwwJHaxpfmIrfljLZi4YylmXV8nK
kbYr28BoD+Ohjw4vBfMtPCQs2A7Qj+tVw7L8H8y5PqTnmoopK0fMLrBG23izDbJaqKTDpnx0yKCB
z+96e7FvzQoybo0biYIPfcf2SoufuD1tYyAljk0T0FCxAZDAUKcdKhxrD5XCwPJi4z7OrtZSBfg+
3dge6sDJ5wEWiDAQHgRV0WFS/0meAGoxrtqG46G8qXZwiYn+/ze9Q1IOX4kq6/VLtQGFdSjn2NrX
pQdnY62Ux/cbhgPZGko9t8+XL2ulNy0hC3d5PRqaM+YWxSkx5UkhaAEhNUt/PkiwcUbUN4hIYFP2
BFgsz3a6GYW+4VEixq7aRm1MSHdobGt9kX/5qCL3UKJvBnmYUQCwUPI7mdpfI3zG6E9K0TZTcSwP
BLjKVM6C9mh2ILwKyOeYXloU+ZNc5RIxXhojgGTbhzCBHsS/r+QifQiLriSoFfEnJUK5kmi7RBdK
2UtZPP215BPTQMjmNDV0gbx7HbNkVmGRYEUa/ofVNOVF+HfdNQYNPSciemDNNlxAV6YgS9TE/Pqo
vmWbIBdRZ7SV3BPT/OjZYJdYS9ymic9b6lmj+XfAgpDsoimIk0jM752Icph0qQ6Si3W0JAR7yLT+
W17elhAKfSZpYYJZ8V09Dj/ZgVxrj3ELlOyhCXAZSG+4OCRCrak0sTeInNSTSOSClSru4Pw5dLcD
RCz4ak+k9xnt3XYKQY3Nlq4U14Hd8gnQTWZcWL4l8MpDP0Tz39UqQJhFoLNxYD4hDnroQCvTj6Di
JlhweSh0WBL6b8Pu31EzblLVZmTxDBkC1NFT3wZCG1KE1Qt68BFD6W5ZFkBfv/sHdJSXmPKzy/7e
LEBSIZqJCgN6vxmRQ2K61SPuS+khRNB5wIFVKJpQV/RhyyAz/1E0R03dEXjsFEZlq2p1tBgn1uP9
12OmjyBQtoojm+TJPmtetBuT7vUXQxQiZdG88RyFP7ojw9tWWy2/Iv4RQ83oMhkK0Xq7yqTZiwSG
sKmokq209sEgqo9btHHJ7gvDtPFnY/R6DC9vec03el7VanJS90Q988Symdps/rHgrE6baM7R96AN
vbi6Nm1PsrJxHraiN6spPxFtTiGP8mlzgRt2Ei3VEu+cA+X05+EqtDhsaEkKrSceYlvVnfTBurH9
kYD0y3lLER4IQXT65Yu7bQC0svFJR5XUkzx2idd7OELufOqp6Hx+lDumdIGiJzRTOBx76thhE25M
72IdeBt9keX94MIcjeVDxAStGlMsg9TcL3vLIaBB8+J0/eVtSsJUFehb1r4gOFPS/1sVO6KypSvI
HWUkkFtGLRxG+KMRslQpcYsB9FjyKLZenBZR35RY5jC+gee+p+Htidyj6TfYaebeOrNEU+wbOlPe
2i4x6Javj98lTNtKyA8ygAR1Ls1IEL5Aadr2EF9Nmv/qg2nO625zG1cvvCra8x2y0OfJeWaW0VHS
L0F4EEsvop9IlCEvezvPzQTrGi+NQaOaXYpP+FLnyKANp+Y9hYEDqdAd0sI+5qoMAPzSSiTjjFie
FG16NsFGv26aACrQRRFfT7nXYPRG/bP8RIVjjG73ZbbZM4whPc469iNilhr/hQ3/63xrX+b1Q0Dh
V7tt7g4NYf9tNY7VT3VKdLHoS2AnQka4SzJuYiMSyf751+OZxm7pP6aTY8TF1u66lH51De5kb/S0
8B3bxPpZBgd8vlA/4X/sD0/0qyztvT+zQ+ALhowpqIq/L+XYK+He9T1KDwnAzpYgmNeJzQKXIixN
YDb47wdsrmN91z7nkqwKNY2Q2Agm9LihESggqNdhY/eOOe/KccizBohJL/AwSyFYbitMzkoEyq41
m0znJDq9/qCF+g38q+3u6NLRkLgLbWhWlnrBvV9mGkMzLdauvS7yEBcqW2qgppedu0dFVehXJsCr
KoWpg0eNJ5Y/Kq72H+p+zG3AL4xXpvWlDsahhE0KQX4lDfZ0QJR4idPlutMUaypi2Frt5T2x5fHj
XzCNNq1SqZEIK5gp2Jk6avyVmzKSGzLDG+1MjsevsouQaxle8k8Ks0EvoD/hOJuS+y/kBp6ti6IL
hRyvvhYG0MIg3HWDpEl5TThJ9KC5N2E6yrxRs38wV8cwmGNLe6qfYX70wyFsmnHHCppOwVISyMx9
BRHqewZE7IWDGRcO3itpJhDqbpaBxvizMIUeZUjH815Ch7MM1kVuAutF8IsdYWzfo8FW+jcD6Q/+
SW1ax3zkMe/LHxPrat5rZMLyZ1wixK0cZjFn9IUJoMzVYvRk1eg4GEcTv/J3qkVDgf2oE/wDatTK
Dmf3EpGCsl3SfJq590MOp+K39mtO4LXA9RSTeJxnCO7506e5rApTVVAsCQhfx7eQ+sCpLpl+edEb
w14HCF5p0WehCNkxjIOEtHarrtUGBJjYi4mSzs00LC6luuS5DozBHjxybBB6H8MXpXOfMRgnw9MQ
pBEYbET1Cou6ylJCdIikaDCDzzhInxU73ODfFWdt7b0CIyTRzNYZCQzEymXlWUQkW4U/WH0Z6dS9
KLS4odOBfd55Qn45/sFqh4N9eKLg/l4wDsNVmqhNPpUUPJlmlQx87Ni0a7kY8+ohYJ/HlCnWXm2N
UHnK5Ah/TPduCc1Rmu5MfqeyxVewpeW+YyoahtiEUNiNoOMexnZ+qO473X8hLiHxz3NGtvGY17E1
UFypTS9H9piXRIgPF3GUq4hcq/Octij+Hsl7ak3hfARvRwv6HnR/+llMTYhZKnRc6LXYof6X4JBV
uwinish2xk6j7yTMCk8c+NE8avNaYrB3aSZP6yQalRxq68Oam6hCJExUyfE9SYCk+d0am1brCm9A
OTKXNkC3bzWFdb/qVhwzujaJmGbO6lIUpSQ2P/hcWZ8yrcUjwCV0ua/or1let15MhmOczA6Qth9V
wmcJhKm8ObeHCf1c5nWt1HN7DG9NyqZHkbxFA4ajS6akFQ2IZVvV9EtuGrW4kVIGpB0HzMLZRhdu
9aP9dlBJlJBOR9sYmL7Jb1bt4dLrJ/SEXyBLlXFh0EzGc6uUneIJbMmYT0eKQGfWcXp7gLeuakv/
EaBGfS+/vhKAMhfFMrN4jwzwjSgpbeYgZv2+P/0e9OCqKqQxR0m1gAP1fiHD74xfekaRCHfjmyyl
cUuJdnJPvZP0PFevkdkBXTmfjt/p+kEim28/hDhYMRr3K7gc0L67vPZ6WzQZcc+SYYqWoann+YW0
a7Wy1AEH1HRTuGnNVefip4wlDHkTZvTFOko6WcxN1VE87jIvjtk6wqKuZbG2qD5yml4zkBZ4wylW
4Prnx4WHDjK9nNTz2HCtf5jIDYCKpKYo2QRJJRhdFNapke90Zzjar2JRgz2XwQCNtxqlq2BjGmkX
zL8WMZXwhuLFiKgu+mNoQU0ljtdN3lv9TFToUabhY6bqp1sLlNalWKTD1UB5ketTY8EW35R8bWpw
lqnLqvKHZX9N91TLM5BPHywBoYCHQyzetJoKh4LoCFRmaDIv180aVPhJe+h91HVep1j5rCu1AWLL
+ob6idBGl3HMiL092iVKFoedfodWan7m/o2VPSoS743id2BY8uKfymoHN7EMXGquTBnlvXQDQZ7m
yUe5gzIxrWDVopvnjSmiUYr3BHR86FSvN7CNUXTqy24yEz8ylnWT9d4PVonRfS/z3bs20pVpfZmz
3b08grxcaDjNsRGaYUstLyfTLsOQKGLGs8Yqn551dQ0bzg4QIZ3kBjvt1e7Xw5L5qVHmg3jUuTgW
HFHTzx69/dvDiaTVzYPDLAtfiBkPMzAeWV4ZpKPh5yT+i6AGJOaJzJH/+Xjd/Am5pFRUHuGqrIMr
YLdOAwe3DFSAaiHZGG4Q/YXKX3tsPx1nxBiBlZiMUpHDD0pzUndHxttzeto8lnIbL+vT77uDxdJy
ptMFtNIe2d4c8wuFX2o+JBWRhTJDXFyhsFgvz5eQe/DbiZ1GYSjMRcv1rZrFbcHBcySsL0N1w3eU
WRt27p8DLz6jfdQjboE8hm7uP4nY9EpLnakz4LeAUbOeexO1l4evRcDkpFnpp5Lt99l2hvROKdEp
nN8ZpBbT68MbcGj5spbEgYFLfDXi8x5oKoh36KS40d1O0zELGxAue2XG4daP0D38FdXuBDcNxwgx
jvIRGpsrMLb9AA69mnklZ+LalHQ+vXB1zq0ocgfUQjV3SHeRidOMoVTxM7CLM23OD6SCQMYyViqy
fG6S4QhaxTMubdcqo5IQCLXDtb7OhUCzUDG/kVjSBmS85/mzF27C+ofrKXM5sxOeibFBBSbN5mCU
VwqWtUMD0SlymA/llZiNdXxEhPQnKZhgQIjZIGeny9b+jshEdNttKOQO9u+MpfWLqN4AFltCgNnT
sTsjErX9IRWYK4PPBrYBaF0SsogmIgjzcf1rRbjbhUGCGGKfv85DySpBoQeBK69Fc8sJtVFcE7HW
RHHiQcZtGNJm/59b4diLhY7ZmSUGwgz8jzdFGm7QYR1LlcjXaU/lomHfZC/mYcMZTdhaurdpcKlr
bYGOHQOMOWI2HjGQ7hgwAhxufailPd+Cm7APnSGMiYccTLIiVjnS6XtORt+yiu0Iyshs1vf88aJV
jDoGApBK2Cck3SuP/k0vAxxLgnknBq8s5byVtb/K/LIOjdjmMfPTVI51934r8qDv15B+SRj2QXmb
HGFsNdleC4Clu/TcbL/THdr3U58Js9V2PoDAcl356syw3xr7Db530O7GQ9D+MDLzM0uABRztbOkq
qY9SvACajOI55mAVC0JK4G5bDT4zvKrjkjkU2R+VWjhlnoQeZ6dXz3Sh+nn05WlQ+4N6+0l5as3/
CE61Enph8iWPL60iEwU8jfjqjqYM5BsOWgNZEjU6SnN1LuTOGGp9+EfS4zwQZdqxTCE6OZnP/8lY
tWf7m2tAuhhv3zQVEm12q60vVJAi+3Y93NjP7LOaweAv+4jK3lP1HQFHI1suUQcK/XuIo0rov3HT
yS2DVZGeepTpI3k4NPlqRE79aoZYoB1Syd2bA751KO49bGV1uECRJ63HzlsnhHkxlCFka5UvhUTh
jSf7JhY2Qa/lUk3W45Jlks0bmQRTUSXfnFa8/CR1t5jGBNpn6NjonjJCwecbhysKQwa89/kCokd8
XijGJhkBdU7rMDNY25krwZFXpGgKAkf8I6pZmOABXgaG1KjNTYFEM7Tv2CnvV5/k7AmaBqQ4y2L5
/UJ7XSa6f3KRQlqmVQ2kjuLZvr2Wl1hurqpt02HCt+whX61z7/R6LeMRdJAxj1nxtBZYBw1YczEM
ouUw6NHI1bIUdYzsnsK8f8Gsc1yOPWLFn2/PCJDh5GnDRHbpd9XV+AhiSIDU7ba7s6gfOPhi5vbG
KMusZIh/MS7xRdWEogJKfIr+JYsCSJfZEeBn1nc/sztL4TznsmIxhsDYi4KZafHQAqq1y2ecPxCs
7AEExkFW5yKrqUBm6i9HVyN2NvyQAERchp/+NpoztRpMpkqpwDDpXqEHvGTyOfrGvcrufnGTRenV
qWoRjja3WawbR5aPz6+z0F+RkD4Z8Un7u2YdVFtavcqvebJeO5mKg8/EiGa6fQsPhR2mv+xqWugr
n/bdaNKtHFRefgWoQ5OUGuHANQdMVxD8j/5ZZri2VIvEMXcRhprEmkUtQZkm06KU9jLCkBmg2b87
g8GH+i+o1VvsbNqZTqTGU+eDQs8oUAVHjYXtcOtTOKWy+OUW5hzBUjaFbxSTUu7LHYDuSZHA1uVT
w3yVif6GOiHdCBi4l8tbRuYpEzIRgpeYjWplJTggE/eLEmfoNBLYc8kpL0BDHriCIRvQKHOZB64c
MsBmYHzwVICeFlE8B6Yth3HCWZUmkd6ITG1Ksv2hHAfrBJy8MnfvZa/nIsJRMtbXZFfUvjX/MeJx
OyRdKDvIe0VzlYk089xxaaGrhAfviTPU6RWgymAK1WZrCtMYIOKLMc/doIZzAXA6KtfJeBwzq4R3
264WWXdafLUzWs3l11EPoug3ii0qTYTBmssxUKvs6HtD9u8MGImk2x1hm3YCkxkX8caZ9kNlmHLE
awbn4ScdlQH9oU5oZKk74MFm17cJv6A+iuHKBJznhROghOYnjA7HkCiBV1QT6X1Cr0osyxPvoTRZ
zcfcag4Rm1qU7XUrSt1rVqAf5EUP4j1bbqYbhIAESFD7NBpjPBNImPk/eRjEr9CxMTjtF/qlDrPs
gisivqNlBRpRpqAWDPtqd/tjV+SNbgHnfrl8TmQGIIwILr9oXn0Tr2ilUALWElj6DPMGJxkupIaM
RTUnFteDui5Cu6Fs2bHcJQdgeyWkMfigt+fL6vLf3JQOLvrpMCbA63W9GseopGXzOrEiTbaRUW4c
OLySrcBvUUHT6qCEgYHJMCzJeBWrw5A5AGINIqFtTgX1DhcAcrSvHn3e4FkiJIRGPF/VwjWEDTFG
j/hQHA8trmbpSwxUqQ2cXDQX5fEZiNWol+8DjtuoapNN97Xd8JXJ0qjw0FryC0uSHiYbALbf7eMx
nix4WBq4IcXgo1F84Hjfo2EgjNGRGsC0I7d3zrucm62ziVM6CHTHs0CXxev8s26+5A1UTkiwQqGv
TyJfasUR0WLgK8GLqjsWIJgSUd7UyKVtDL8GbI3VdlBFs3uBrBBNBQujpBQmG00kZr97M0MfOLdt
ubklcsPWicalKmd9St9V85IXaZMt3YHK+Q+OrFy4U2yhKVhlgIbV7EYKXZoUxVoGAMqUQOUhVyNv
KjpHggdEwc0W70eJWIhWERGe/H+5RFAlE7trKeiqE2NtQZFnt3llToCdSHTcJlaLz5+54QyaVXlf
2bK/iobkgo9OWAn8IPgADLYOEmHCVJwg5snURV/1awDJb0UhkobkeusNp/kO2Wun14SPQ47fl7he
T5WdjozoOrQOMwdFx64+iU/VOZKUoeFN5WwcHD+NjodjVsdaof8zbpTETvG/irayemnsWUAg9vYD
hsFdncdnKjtKFlfeRa9IGK43tcCmudJtAQK/Y4cla2McleM/xsyrUIwYZt1GGUnIwU0MSNE7F1F/
JyRyi2pkWBjT/VvuGSCv+JKDb8P2ca9GCI8FEvsmxbLpVw85dKUzWT6WGjdNLCDug2zcOGqZo3n6
CtRtSl+NVnj9i1P/agth7wF/2hIF4WF26FZZ9lsqHLDGsGWSNTgCpPA4d/B/k1NlQyG2XyMVs+Rp
O6OkH+nOib/+MJhRE/Md18qoHL+PjiD+LeaP1F86KinFvfi9vxpJ72KKdaoTc51NZWLSY8xGJb2q
VnXFrWAnxKtknuR10QPtqojY/cAL3YEEip3fLLv1bd4il3btu3sMYOikPbDRrt5NEqZX0vHBlYUQ
65tHgPLwdmgF9Od8ThxZ3w9pFGopLghRcRXBdFQinnGbymyKWjluchjIScTyZtBNiUeVhNyVYFFc
bQeBA6YCvmq4kj3gezWsYphcMNKU5cIS9oC0jN6BhdC8vRzkY9hM8PhcNrtjgKCXNqHCfyLUqZre
0UCFMJMALHv8zOh9/hSqzz/VuJm1eiLw6Q63n7fDgDMtUVEORn1arXplx0sJhyKxzFY6mQ+KYQ0o
nK4LY1qI0Kg8ya1JrXX5Q1aC4OrEk+lrCe5wzy8YLpBYimphkwH+/v7CA7Lm8tD3HyRy7sJoPmc9
jqZgqxirsjCe+5MXL3ekXsqEIW/z0tNGnuQh6rubADZvTaCACFjseI8O9N9lZaXk3RTMiZM+mGXs
RxI0WdE58H2k+7qMdjXhEu8dKFujfd1NF8oLRPsZqCq4JMPa6CCmwMDOUYeN8/zi/hvw7jL8wCjv
3ExTGn26KI3nnaXasQp3nNii1W/kzDhnj+YZXYae0UnA5HNkXGWfbxCNJxHZWipg+55tjTobyn5Q
jofvgmCitVLpnhTBmo6j+tXBsAyV8F7967gImZBKF3ldVdgvxgy3Zpnsc9/zKe9PwN9sCtGOvQEK
QNqeUiPpd0fT2BszvzcCalvdLC3C0dwH6S3QxDSgEpFGnztrHm9Lv8L5DZVp24nXF1TXHTt/tBE+
mq7THUIamRopc58QuHc4Fl+7xJLaBTwM/xLjS06nZNTD+RitcGZtouFWsP9LYtng8LJof+cNblkD
bi+bXWV5C9l9Dk41xRcz4h1+I1JTAe6g9iOF09ArAqZjKtMpKwLzo485Qc7Fe262+w4lP8jllraP
ncYLpB87cktUysF+Ks/atyHS0HcdYNUaVL/Otckj/I+orXzxxVYzzlKHosbPAEpELzTJTDbJgsuY
/TWlcfFFexIir6OTmk2J3AsVelB9HjA1/1u0Yt5cz6nNyzXgkjBZ2+GOtaAuSxs3gUW6OVuHrFTg
ZR1UNW8MrK3RSQZ3pcIJv2Pg1BForzFYCoCZ1vvu8w+JFqxZyi9OECxUjm+3S2Jx+WlapqWe4ZgL
gdgJwkgS7r+kNe+95ndHZxaozidQ3nbxmAbscSl1ti80JWyZG3Yo4CORb8yjlLw+0MKDGaBlwphh
pQsup7W7dWsjgk+xbSQJYUAFN7tR/3Z/Ie7g5SCiJoBj9Qjcs8buTQP/oOt3SHk5w80YtePgGSi4
9g7PyBm0ZIqeI/kRO6Id6zFiFSOOdXyCjQhO51HqWkQL5Iof8EWaO4uS4Sn7QsVsYey3+kYf2ls+
3FBdyosGXFQ3bA1E30LvHB0XPIlKOPt3tPG9cs6fngsK3gikTloxRxsw6Ix7dLrxNomn9h21mq4h
1CCXdomRFWzNx9/HboidRaX8OzSPi7T3EFmm/QUPoSLNjx+bEr0RmifZLJ/2/EpWNIfrVi5SPcvA
PsfgRt2uIjFz6BaVYYEttD8I9bSt2KLISKyQHRggHYrDEjt2YHks6s6N+vDoUlekDiVFtRLWuVoN
8jB4kRXZUo4vuzSrkF/fv1wwHiqp2Uxsw8CfjKlL/saP0aH52KIffKJ8XlOc/bWkkMgDFCj3hSo1
YOi1pV1l1gStbO9dqLvnvnUTaibTkM6zYGoYjD1EJ2AE6M8u8w4R94f3OksSOqIwmHU0kwOC32vH
OTp2YVkgzX3pK8BQ0GUgnkgBItn5gjHjvr9Uvw5kOuf+0DxboeQYTraGE779W9yGRpCHUVzXGz6i
qUNYH6eslJUKP5HN1zR1CKtC0ls+ujDonL4QG0EJFdc6/4w7XWZH/Lmq+PvHLpYeFb0qBGqZJ2x2
IXYlZA77eYRhjF1TuGT040xKk5amLIVBoNAZMHl4lT4A2XpgTLqrLgq4Y1/G86FplRuZYhc6s4H3
IecX/wbTSpFngDKN3rsdKoXmmqrme/jxCIY1XkZpzv/YbJucNTfL+szgSOx0UnFlDGDUzGNSpHJl
VT7TpiScujWF8Jo4Au6wdjvgHEIQf0BOh3XTaWNxGzU9q+x/ligGY8pF9u7kmdfGCsIEyIz3IEoK
oz9L0T5S0HEU0AY4P0MHbGE0hVgsOM2518tG5ixww0KvAJu7fI7YmVviQFCca3ajQSX4AA/iJvyh
4YPlacSaTuuBn/RUDOEVdhFuPnqzAEKpAApZN6BonT785IV/G1iq7vBtAo8q4MFmj4Iti76MGU/P
UxshdfXemiRUhiSBKe1RTgzsl3HNGjk9v8GZxGRAS6roq1/8xUE3rWsmwV9uwjtgIUns5eO1O8pC
Rv7kXM7OYhp15JV09rUNoRG/VlKDLs9HNCEh/i3FkWMh/NBo3AA0rEzw0wduTUvsFEgoS7iQpmAo
sE0TqQFmbXyNMc0vcSIYtmruStN1O1IzmwypZoG5ZzBs2/1antZr5w7qY6s8xeavKPt17ikMkW07
XSGpDH67TfuW3izHP2d59Aq/nvza85b5NaxyUP131AeHivFltKkLGK8/fBPUI1jmvBwzbOEWm22+
/6sR0Te68+/JEKAur8wODV6EQdBInNQWIbnppzKOEAGTfXoO6wI5n6N0yuUVmNK5+gghz6X1S+iu
ljhE6G/mxRqfsUeqoyTbaJQSBjqgmHwy959OEQXBs3jPWZTbjRKErHM2KQE2QR2T9KIiMSXkgX0i
F/FKtgN4jIb6JDVteXtdwWrbvDV6Kv/S6HtmPu70G3/atSjJHt2/mMzo3XVSTsO8X7Ydz/4J0tpN
G51hjgc+S1nh9lR4D03JeFJsrZfsF6CsUlIa/OfxiwTtimddSFIVupZO/FJnLrfQBHEYPgZxuVjH
fdVzyAHwri/ZN8ylLpuU6X78Fv+IY6PlIhgHD2//R/ygRTOJJcDlz9J6CtkVPtZfc8gB+4gLgzMu
g3PlVTGJS8GIE+3XvaHA+iwBV7EqOSysZyLpAkR5rtqzgw7LcDeVQDDfswTDYLMT/6EwbitiC4Lc
r+B6qZwYvP1j+UfnCTM3By07sNsV2tKSxhLyTeU0hNC1wZOuGgCGUPAmcLmPL8y+wi7TfCd/zryc
6j7bpndcN4hhf/yIhaB5IqWmM0+6rkg+Hf4hnhDNDMUofUP7Qjt2Lr1ZoFhzpO7ZRRWnFeOIuHiV
JCUsHXbb1K7p2Yh/EpIFole1ENZoYNXu5vcEMh0cOgXJnXwLVUSwQtmEjCWqR5t95CxuXuTtZV7E
l7t8pTHMk4N8SR44w0q8kcW7sIgIjvUYVhhEQfOMOCp9I0l3RoYICdOPZ55KMF4cLPRGcj4MeEKM
42QEvRf6XhleZS+05rtUfTaUhh4ctLLYk17d2F9vdzefd6/jvFQZOe/a/Rd8Dme8nxTYPDYpzbHi
UXEPCjzIFxF5Yca0+LI7nqdlvTb/cUp7AwvRYEQJtnRK+bOP0F122RC7TkwTBZRh93wGNPdS9z0P
vfW59iER3bzns2Xk4xUfFhZLzmSLhKZIRwClyHg1C6gV0shEvQ0lvwhAEzvQ2WfWaZCYCdQ0tVmr
X2uzuV9hcD6Vg/NOKH1SIHNqwmjzkkbp5yOv8bjiw3/gn9zcku0cfbK7NgWfIbBriPraNcgCI7tB
j+8J4G17D+Wx9u5MrZzRDD33kcZkA8Na6s0Bttd/Q7FDqwBDMTcUO7eLANp54RcVa2vzHzxAQBQM
+gAjIas34It/8BnYVwhmSelKf7T1nIS3o2QRaUokUo57cRXgCJYi6oRnEwDMXmKnYUIGo2dlcVUt
GPIxhzPi+Q8VXnTiYTD0VvtwcMun0EwUwUD+UBJA5Z2bZJE7oKZApWWo67agNX5vhNRF7g0ToOoB
xB53sB5V69N7wcP9qgyGPmRjtXkg12N5ft7xX9VWuSyx+AwvQzZXig7EhrgUmAbnaqhI2PWcpY1+
IXSlj8jBusgNItela3nVVVd/C/4M9uoclY2ZXlXCTXhFcU53WdsZYsmM+IhRPYJXv/de3rhQx8U5
V1CWfDVXmCRwNoyTcJUvmfDQY7YBXEvjyE9JfWYLwi+3YUrRXSMQMRFbVj56lqr6IuHsTptPutIq
rXe/AgpvJDAvvmzL0TOcDn12UNtydXahxaYekZowdcss8naaKJchjcjfoIh7r9xXmF7OK4Lxt7H0
fQylTpcwTNO7XtAJsrIepNBgPavjK/Lh3BL8z76qcutxTbItTDtBVzl6qu7QfP9GrzXZxYtyeuHC
BJ4IlmELz7hfswpTsCXoxn25Ko3L2JZJf7LtwI/n+B/uyq56Fi0jDXhr4JlQrzgRmvaq3mIMpOjh
O68iVfKca7WWJsj50cUmo2wwPivbt02ZhEaKUXgwPTk8PYLt1GKzBRjblDproy4KEG4xUHRCpPn9
nqd0wcp3oMp7QuJucOLWOKPyOwaYglmuldot0PaONrEvm3tpPDAzf5mVlc6d3K4eBQsn9i/xxRwQ
J+0n2j0T1O0jHohBGq5LbNCOPlF83IFjNIMy9MucALfc5d6FS04Y9bWXnA1PsFIC0NrKCDlm6qc3
WZqx20YZl3ZYvssd8rRejihHr6Wj9NUR9p2xT1xyn/QYTNBsvKigg/qhA65aaJylsX/1SvqFGj9T
57AiIsRd6DxGX2F4EaqrIc3dD99pGSTpaePlLeomxRT0VS3BIheN4JDU1gSOvdFcTcID8AuvUEY2
dgES+dfSbH39MUdIDdVQprqbomBKPR/fvTmU7iyBhHjpudxXpCwubMlCMDw3XT5VDdgtykOJ60FI
vMa1WEOwxj4Bs4uje5ZuRM7xUV53zAeihy174NIWrosouhhcX+nluntQPyXoGlWChFm574iGd6ZF
Vt4B8bV1SXH+jnujf8wA0Yp1BNzNl2PCgPqbV0i7yfZeLDtc3OXdD/yPj7mMFqyI5nV/1OQfEf2k
b0BnGWTpq3Nf36L4xwFDLXIEpQRfjIV6ZAc/xmeU7zTy5lYY3i0ZsiG1RMRq2JTN7aYm9hKvAXwy
JRExAE6R6LCdNSEpX7XI1zhg/JwJAqan+b8mAsw0s6QaDU11GXTkVh+BM1J8PgJCj8qZmXQO0KT9
6jmWWJJQ9Usfd1pnW8o0g60Sc5ra3ZBLXauMrM1qPBtppCZPAt//GHX26UHvKz++6NxTOzhQTp8y
FVGD7XtFBi0fjxPKHKlWDHlqAm7rGFKmVEU/6CQobnrVP0oz4n1bFLxhJTcr8fpeVrGOufbn/dtY
P1RLGw1HiWvOwz0DEBYE40pbZepFJtsO8+mrmjOxEqvAXXkIOiSvC5xcVj180j4q6fMtOKHDjemf
cH3F4hvgbPZ5URsdbocSZ1UGKoGsqgjDB89yWZknZ1EAfUY6ho9LB88VWIjpoYcegxrtgzdmDviN
H7hznGUuiemhaCS8OVsD4ea2wnAjhoXZnRnp9dTYb7EX6jsCfPz7TMboRPTUSV4PfuEEszlCk4si
BymoTulGdByUrbesh4pL6dwPy02xhTukgUtgDtUQU5yyMaVbO9vEPWInKRHiTehyjsyQPNM0SMEh
SJq/VYfNox0Mg+78XLpk3Rh8OENFNKBwtZXZdjY5IKMFVyZSL/+l9MnR68xkJhJjSiAkgj4VVC6r
gz+uwFFC/BuRGQ5vIqy94+gUJp8eP2g/OaINbD+rRn6cs89ShHuL8SDWnJSRENJ12vc9Y28u10I1
Vc/WBS6r/VqVClOauPkCV3GUmr3adZUDrHcaAJcR7fnY0iOCdkJV1aPCW6yxtFroGoEUSF/dYjWS
i03xD3eObvSKB5B8UyR7PTVn2lFBUKYKrkXzpUQYGK7+OUdTxXzskc0WegvKXPZrzJ4NH3FZvEI5
TSb9JZ8ZjTM8x7wrsun4nZULwvSHEGrzHDYlLtV5oimk3nB6gVu9pWIzoG2DX9Mg3tOpC+BGIrzA
Ms+zv3/NTdlCdxHADtO9zMniM1rUrRvraHPTgD9djKPhjFcXGzVfJZPpOkCceqJTvIfClS7r9QJy
ZQCs9tgsm4Cy1QA6fMe0jsnU2O3yKI3ZP/O5GHj9cAuf8JyfU5q8Ng8TvR0Ty+ISr5+vKlYmpLll
w1jUjDttid9I7pTB73qc9EQZwxPv3RpmkMcgtGqI8vpPoXtz51Q+iTNrjp+/wCF3Jgl5Bhst3eWX
mYN5b4ESQmT1eHXSXSYtGKPkky0GzPHqT+ro9AzP9fcmOAZMvYE8dLz3gDguOcBRFBJrEyg7QrPr
/0ac/BxiqGAxcLUKRDA1/XDOcwJ1mBiguqN1ro9S2mj+pAR3wuZKIjR8aELCbxlDqNva/TzBN1WJ
7QR7zl0u4KgwM44+j1uw8PJ+XzC7na4p/WGjdk0dDjg9ENXaqxRdid1cYZ5GMAmmC8cgDLMCsYJk
GokPt6a1YMTrMStFjviJHRUEfjVQvbbcaRBuTffP2BpZ18ETlKphy0rx1I8mwsP0vJUqL4F6ZrGR
Qqk0ibgtbTtWuB891ALHI9Eu/VIreU2HDrxZ9/uOzkSoYuQaYTC9HkMoaS2pfVQQT25das3uqa1P
iwDmpxZsS2XSBYas9SE3GjKGY3oXja1PZopcuWIL1Dj7s4nNJ7VZRxqQobIBjXtuJa6u88u56uDm
smOnnq28QosgA2FQKrqB0CEyWu9/ywGDF3H+fNpDRuNXEz/csypiC6sJdP8ghawIxw+kKQmeqPk2
/+HUw0UeQp9saezRXpE+XWCzzsbAhNdizNJuofRnHZUcy3gLfSYTVlY/UxHjn+p1qyG4/WOr5t4t
oi0b9iK1NhjM1ISxSjuBP9VvQO6u7d0dsbHtBeBFKAcSb0iAbm4CHDKogu1zWpgVqe4y/OMLFwgs
aqOukWeclp3SXklQbw7L9MDRDwg14jZHsWHJlkx/C40xj+wkyE9WD/w69UitnLQOhamm/bjKN9V7
6Zl4vnizkgZzaIU9/PtkLmUy5WVDAjzCBvvCivKtfD9ayaxF4QigruHjxgJH6O4FF4Ro8SwTwS7C
zdmQMeq6z3AgmLujhXy33TFVrPHkXfvIntecfLeuQUDonPV6AYC8yXjzG+34DkYwGUIi7QwCmGjX
RX+NaycPQoiPv4t4Sq6/IyxWGggKDih1OP4bDY0PGEk3dbT/QG61jqmXsuv7PtMBX4dk9LsAsc4T
3P0ROZk1mRURtB3iH3UZrY34C0O1FNu43z8oYoUFOJL8rkgjmoYBHQzWvyv/PFEUrUDGLkWNtJXA
r7DfAex6+CDhEvjYlXpJqM6OGqgfrHS1RzceAwZ9Md1wqGro9zY0TEjXtvKQcFvp7mQvYCRbr1ET
Lkofg+Qcriq6lRlkCnMqsNr+fmOQ2zTRuqFb96vftfJkJc0eVR0xrpLfRvBhRdSmau4XQqShW0j5
U4uCef5QdrouIiZ8BHF4r5P2u9b07MB/IwTgyAjVwS/LBfUsxkuUO3VkBFKzS+TQ5tRV3zerq1e9
6SA28AOgZtbt0Xt/URTmDVvmGaTBjImDMCAyKiT+ozVtChTPtdBY/LRgOX+t5RpBZP4gnJQqikw0
r5lWJ1DA4VDNKeYQFUyQVF9YaT0BwEtpQf97QON5bKnTtZZwKZRRDzK3G6qZUqTWGm2qhIwqkY0V
06dVQXnBpfhdqi1dlOEBpfpW/1Uy06/8le3o9wcxsZ9OvWme/mbsq3JmPn0mxkItyUqSe7NCJNKx
jLS9fu0YZ19oBWq62y0hmJHeBkZcLHA/wqVC6Faa77cm4zl2Ad7PgpJOav2GtpH/DxO3Fi7dosj8
QDg7WGKHP43dHDaWJQv/WoCPWI/DY2w2yiVaC7bRFfSpI+Idv49DCxZ98e3Om9j2A9qxeqLUKfTk
ICuLr5GzpFBA1cuj1dfTrW/nhDn7x/u9pki5ssk4aXV9FNrpeFRxWMioLW9fuObtP9u+ME+i+dKI
i+d1ogO4JvtmBpsV3IPVyRCbE4z4tstksy26S22K0KLN4VSVMMTd/kbmEbgWPe6IE/aQ7ZR5qwd3
w6h3E1qYTONR5q5AykAFB4q6BC5oi0jjntCduoLe+QM7v5TtvS5K+6ceBmNU443vAQGbKzYkr3wm
Ih6TPu2wfK08n4ln3BMXa/782ScuGbFUPouVHWeo7uRbnX/3Qxg5QyBeS5zI7DwNZbcZjeDOI6F/
bvTJwu9r7d5kj1Mu1ynskAc1maouk5e1xGoWcKZf7FF5iz5OOYCpxWI4bhWqmWrprPQU55+jYVcS
quJzKZ4iB5Y1GFgMmkDk40zoRwDNcGj7CDviymorU0/42V7vrLnIn2cEt7UVnfBCLErGKOCC6yXH
rIbHnHkS8Pjv4QhbgJBP6qrG6pkv6J0lKIQ8LvQXip9md8crW+Xa/KGd08iRJRjrEjCOLN2Swn73
s3ouUIPxekEaPHzKH6AIVX5cbWRZSbPDyNFNpwQBzZoKvyq2NYANwbGsMoD8tRZR5BS92TRwUQ5Y
iJQqKjY0iQb+DdKkzfqaRwNYwy53qM083DzV81CsHBDY92fkSBvljaWZR4VaqD8Ka4aOpzhMCYPs
YBKhAy33oDuoQx7dMJMRr+dNK4Stvv+OKDrUTppVQ1lNoSmavdRmD/5M9JHcfaqeiX81BqUO0jA4
VYYsDOAeM7UB761JhcIHJXmQJvFgyxcHBItOxadmdLE+PS1E0X5FL9gfeeFZuUTv9s0ErA4KCVu4
qAqQHOYHAKyzWr/qP4uT+o2dTmF2PfmI5Gwif0yUNJCgNlK/8p1APTsAY8PSPJhg67i9bflc6v46
NA/MJD1T3tL1hmYSVdUt5mKIcJqGS2hN7rYM4pKh5OLkQhNXBTFJcFghaGkqQ+zSCqJE0HeS572D
pTKxN51lY8le29lxl2q87gonrfv38NSx8AraJf08Sampj040cC7UiL/2FrUl7Yu6tSFfumb/pNkb
4jCmspdDqDggjbuvoZICpGbGXGsbDDr188UgXSoZjwvz56HZpWO/VGFguQMcCJ2zV7YtDSm8miqB
vtqIroEuTv/YbMQJgpCG93XvvDa8ks2jKsopAJWT94GGMyBpozY6xsj6ah5HDHM3u8DrucRpJVTS
VDs9B+zedX5Xrtc7T9S+9/WHnUfNhLksDxr9ks7vecO2/BtZhIp/rUqcjrbVXcz+pLlxjKkMfqST
1bVtixdJSa+UsX3d0gfcC5EVRTNUiPykLxG3C+LSJA01EwQ6q68BCRi+1yjKV9FEPEjSDTLCck22
jC6XW3FuJzAmu5/E7HDmD5kpX/s6eEOnWzaghG2lLu36BRMFYj+yV2N0QrtIgD++WdGgxG9uFDPi
7zEkh9SmmyJKbbuP9qzDqcRRa24qoRHxKsj2m876ggws5a02LV2Tivbd6piD5ei+M/f0hl724JQv
rDvjIbEgl3J6nUA5CpForHB7Rmz0Pp4UcWN7Kbw1mzITmUjxG4mAw7tdrNEklijh09yn+mfZ3rbi
fVPuQAWITN82g8znGDv9zjKEcitcVLaI6rn9J8cii2h/gWvMw4IeQK00xEqvNAAwYTFiXvF+jA+Q
T+wlcHYp49WWcDQUwouZgHoEmowlAIhEbdJhGgozNv/3Jme1caRb0afaN1zBG5piwirFnTq2t1NR
N5NwlwZA9hy/1kyi/aW2NlOsDx4ZCXW3C+mu9uITCPzR6c91Alh3e27LSA51usWM33PNBSIdmhmg
8lqGRQnr7FNgUK6tKY5+vh9kLf7XGNvbg6VbQH8QL9Al66ebTjCjw8/3SeB9leZ+LnHfNAKnEjSn
nakua+KIEmbF4O1WP3dFHgkt27eJ3kxJWK25zBC4byCslFKM5NRnLCh49zPLPBb6SxOj8ts7JJ2F
JjtrA8a6l7C2k+JsCRk6sPdkz99GLMX0MvK8CeUzBXbmPPg+lOB3kw4fPCJTiHmdJX72ChWYqgmC
bF55hG6zrRfQLwWhrvOUtJC7Vmqjb02n/ibFN85BfjdAiN0anu0lXxC6gUFZVSq/m/mwUbzjQ2C7
yrQxN2TYOeVYEpNUe/vJ8aLJtrrO3QCfrJ1Brc41mpE6WnVPHoU3en883hhv2XvxJS1DHFS462Vw
1osRJ56FXMKCradcgbRgzFiTi8WJXWb6otKikM63unZQGBNmABLkcQ3VLVzeIUVD0VoqrpU0xO48
2FgovSjJBc+aLHQuO8LxIFKAihSfuc1kZDzfIh78jtWSyphIeEG1tqjnkYn8yvqowsw/HHEUMSNr
p0OFnsJJeTu97u3zl3w5lkSjfEm7YZjci2UhS50zzZfFXQ6sBN3ObveqcQfskEK0l/yTp/SMbhxz
ENTl83ygH9mYsIz73/1w3FPkBZdRTOLnIIbyIGo48+2FzTKZdZZr8fi/JdinRx7pqS/ZKfPaEpGx
r19kJwAL+o0ljtYTaH7Hq3+o5XfsiFq836uPBmTYmeUJeKwhm0OtrZT/6N4eI809PSZqhUO+5Vbg
fgER14KtAi5bgV/me1keflQTVnq4anx/Bb9/2So3ke8HNTqccC8Fi412wO5mJ77zo0XJB+O+5gRB
V17u1N1rA4Jp0H1c8KV7Ds/SnLNw4XwmgjD+bygR1srTK21ucFNdtHrber2k6GtqVct1TFAUaarL
uXBKWl7RIYdCvk+rhQINH6hVXl1iWhZBLLdBAZgVP+gfiYVnuVoVtkTsGg+TFMIagTdfDEXe4HrI
CEhbD+iDu4wNJqOkCEyCn/pk/ZO951pX62Ue5BUIhPORhO+309CYE072eSQUgjBsFwjhMnX6nfNW
F/CYwMBvxcpS4IuEeqw082BZUMSZTk2hBaPouND1f7RgnR3W8CNt7sqZaqQVHCZ0uPBYfT+Nw67U
1vRXMwxGLP0bA9uxmz6Cu4XDnWuTXUWgofKwu32oSrAiTu8SPmptd54KOU0GwJ2I38P0ru4auCbl
S+TZvAaeBrhWJyOCeWt3icfLFrXJdkOAqCCKHcumSquf0nriKbN/VrSDQIJokaH0CUVTDku5jtgc
QWPP8Lp5df7J3qLJEnOdYvMdyxsZ9m6y2kiXQLwW4OyKjccZK9LpuIX5E3Q127Tohb/d6qigJb5y
5O9eFwj6kyW2MmzBBPfcsjdWbJgdxCQ2nRKn5MO+t9W7tM8LJxJ0EkpeCF3OTCPIfldF4rt4jzA5
OdbgKyw02Dak5WWxdV38BFBRgbBoBhhMZFGxVvLddx8QriWrxtJ7qfH/VWdvADGhy+kho55cG2rL
hZymi4FgHA8YqibjZWoBmlqFgPga4VtO6d51+zmKosUAYUh1pOtD/eYgtFRJLVZatI3Dbjlt4kmb
4vlVKSovzKu4RkJgYUmqo7+ZVv0HHRrFa+q9BkUIl3zRi2UhS4Y9LMnth9qzYEoNTgrIq8iPT1cy
l23VQ/ndVuVmyILpOj5o08W4K83skojednQ0jDnvMeNM7jYeR4cu/kARK1Kr6JR41Y0ohM64ITcp
uJI1Ds0dBwbi6U4yUP3m7Vtvujs03VmsVpi2py+J+dKRnYGE1lAve0zq1T2YyEJv4I8BLmrL08cd
jyLWQp8Mk2DJEyeouLSAG0atb/HDo6B+P2S5K2/EAvFo9wHtQZxNdQKhrMNqImOkVLWoOZb+vASB
e+P9DtxE7zk69iPU/VR4O9XEKHMmY842MWxld3la3hGCp3Is/3v6XhiOmm7yNsWnmH6oEnP1Ad3O
5ZNyFF7rYmhyjSjnxjkWkLjZSUnvTnoBG0SBbTfBDRus7+NsflD4t+xEeaJH/X94Hj8losucZun9
asWnobcFVP8lRb1ocuqoloZqG+g85bHCkb/g9q1pU6LJg97WGxSBE1XQ/Is+VgS5eheaCd1qrgcS
ZlkNWOSNasGu53LcYmeN/N2rZqfFmlQ1ZFTbQMETMPIr/2jyI4Td1hdSXFQEZdrbWRf28ttNjH8Y
/FZx8T9vru2S2SjyqaAD37T7bDkd9u9RsXQBO7chHD+oPUzxtrtsON0fxwuQloX10tWlf6evig9y
/TfqurTSBM8odT3kKOE8lTChyqdxNfy44VZi+kPegO0aqEGmcFAw2VBe96hAf1v9d7+KyTCX+AD3
WX6Qc9GeFP/1egfVUcdQopWuiNx8Gh6QxcwkFrwQEQRjnM8xNLvFd9rdpFYdEvvhZCji3dVDRqBg
i22JxGN2Rv2B2c3b4/XM1M0s4uVChPKjhJ03zu/skULY72NKwMQzLMK7qOB0o9jUr1O/LQ8SKIka
NL1R/aU/Qo59NClIXzfoY3RFcHMe3MVtmzq6jdMKF4nieUVfhKhBb81PROSvlCo7QzRPIu60m9Q3
fb9e3CTXyn3v3FrHsJ+WjZji/xoyfRlz+fId4Uj3NiCTWOgEO4fpdWpV8GLrXBDJPvgZuhvcJ2fx
TjJnJSkT6hmTkAQSCczgbE6xK/SxmTyH4KopAlUi2cSd0a9wCkuthc4DMj/+DvQMm2SmhEHYW7Eq
IkGzv3HcTdNzRjHgf5mXBJ91GywjqAaltVp6T0yxLdV3OKSj0Clv+V9BJom36YCCkdDUqNTph++1
P5GLVt3Eqeb7MlKwGh0cPy6c9qtFnqhi8q4E+v3wsG64WkWd8DYnuOcEklFdPlHFSgfMjD+mOWq0
ytYMfWYIYhM1V5bWDOV3IMm24LqXUnzHkBd29bBQHfOf0YZ5w9fH8JRaiEjnRWKfBlKPByuvywqf
2uNdSAB0tTGPMlCfdrkUz+gXiPcFobzzC8CFuepcfq3aYsHBhgY39NhqJ6KUTPqBvVlb2gdBR8QZ
GWd+q2CpORAhqxAl1oaOt9Fbhv6NHLQBBxA5T7jrDQERir0XhH1rH8WsJjV/ot2SKKURWfP+ar6C
U4U6gNxUo6zzx4DdP8i9VOvw2vtZnVd67yirZqcyyQhiRnrFBhX+7YP9XeqUo5zvBAprxA6+8B7r
ZQHr9NcHxx4LtngOuM5kiSijISBw0MGQcFQBpWhWw+KLpaRowBRlVInos1a2+sJjSdniPcvjaiBU
pIBioYtlOKJpYEund2XYYhFdxBRvTeVqiYeJTkpyi0ShiRGPOk8mc/+NajTqgae/DfyyfOCO2WK5
gzfKV80GiYm0YViZE0mlUZWHPwZO5NiJl6JSWyrNQBDJQl7yj5OE+QDNT8gf5Lfpq+aNEHChQR2A
d6pDdKrJ/bMZmoQrbAz2FBn/RiMs43CJbdv0Vai7Kz2H9ei+3pTq9md4z9GZz2fvvvycsTI8d8sG
5WaILuQbN3cJDjSBjbSZXIVXuXB2ADK1qWPwLPuQ7ufNBd9grjCfHFsIrfF4wwg/MXZ76tHXOoC/
7Tznwiuyikh3G7LbzugUVTfRx1rKX5J9h3mUCslThagLKvPCsC5YK+aJ7oqkbaTycn2toPonVJ14
67RC2lwMVWIvP8YA36fmarYCsR54Hz8AOzCs6bSlaK7UeUJUu6ArDTuab7adiYmD+F+aUb5QaghG
brFwTQiRH5wRHbjvV4m8HaHRiDA2AnilWcFr1a7G+MnvnJYE49EGsTncgYQY9ZWa1EqWHwslxrLf
52WjVAgNgrxiZ0nYrHGeKWcH1LDMXSOuMcePbeAur9ps/GnIT4wLtPZ7zQo8NhhFt7hj15WGfgqa
p46sLc6OQ0MjXbTGQn9lDpOw/DYAhRspMM/UlZwD/gxstmrSs+PhBj9ONewz1YfWsSA0CGKn1a13
JPoZZce/s+AL4HUJcboI1mf3ytUSvVejBUldP8fYnVhxRwGMiMBftf0G701Pw0VQU6OcbFt0hGEF
l4EmfElA/HWkGwJte6OWT2kuXDNSmQYz12rMgxVG4XbtlihpA/HMChwYRdsfM0xI/6gLPiqdsB+I
2OyMy26Q3nU3A7lbxh4elZVnTudL/CCIuDGRHkvrFoioW2TfYm2lmj6SJOT/kScnZOF8hBZ8v5qE
QcRpxIR/TPh5YcDSO6IGagCWGuXjhu8J5377B4bNMxQtdAfC4UK2+8+aSsXIuceyp6g9mH5Rqqb2
2KK80QpfwFv6p7Yi2zfKwjw0rCWdXkgciSFAzNvYNMOGSNF7m6LcVSx4F5AlE2RhYFpSy3OCRNIY
OEa1f1N7k08WnswUuLsa5brtSbhtUMko12Rg8YYTd38/e4Yi9woDpVISfJUU7L9N4dJZ75iD4Qut
VwpTSvrtEqSKZFBtrDVYe4gHZNSTCAi1SdfGflOyW2Y8DIOb9RerwIctfV0Htq3FTUxlmpflVZq4
v44LpxJTzBuqA3MNYSljAISPCAXqI3NLnXGq7f6tQ5Z0tOPZGPqt15NpDurqCIm4kdl22i92fU8g
Bi74YCPxTaS1J+4MLLH/xGbq3zXyditSuzlLsJNdqCX4yrS+/0C5uPU9qoq5ewylVzUOBkiMti5R
BPXuB3DcWeQppdEfJffUoQ5W0VBoPR77K3pegW7YNh9FkaP3oDfw/s3FU94LBC1BpYV6Q3n2TkMn
HJ+maeAkjNT57AK5TAj3Y8hRLR9uCWe4dwXdmo1HuDmFmwSVhNOji3S63vFoUxl3BaqKvEMQB0PA
JVO6oX+9BHQ3zYk8wkLgVbiJwbMwg7RaKI72J/FGw7ueFA2eo5xezQcddJ3cC+WN+i0r2/tWKp7j
X6en+KJp10swrLhtkDShgesGO42tzwHYULJPKDjVFJ1C1O6Q77YVJ/gmCL89+F019p4SGvndp3wB
vI0bo+VPXZp7qjpUFeAX7UX2O72KsiH/oRP0DsUPB1SIQOixc6EQlpA+oc9IByQJCSKF7qYF4W56
u7cONei1L5XqqcgQ0+OQcT12RW4/T9PYAROSyzGTzIQJ+4MvluIUize+cAMPvjeS54ea/o7adQzK
vBfh8vhGyIztXn43q5RgA74qpSbzoxtQN8cN2AA5VkC+dXxlbMUqPlSD1BltwnthNVgNREhEke+/
mNSRYAV+zKSUO62Tpd9ZBG/ci5q892XlemVlwOirAHCLfhMdZCcC1ShNpu20KafcsVb1NmWYOdFO
G8SVCtcqBw47Wd3y4+0X7/9z31DH5TOJjK2A+CwHLJ2xYzHHpO9M3jM+Mpyc78snvGtd37urCiWX
Br2Z57CZoMZY6WrCJ/4r5LyI3h7cJutfrZAU0MDzsTI3qUgjbg/Su0Rxsq8JSFbyUVfoqUyX2SN3
Xg5E82Xn8G6EyEi3I8iy8j7zxSaFHvlvEVF+Ppo06lYP7O6Lj+n9M/aPEt4h9hot/eU8lro41pXo
zarfMt0ZPlY3XBSdi9UrpHDl0BdiYIyBBeyj/MdwnzLzwpoXEIGNDB2Cw8Ve+aLGsw5g7uBjdS80
KjeDDz+YgRW/PLA44d7MV4bletGkvlAJWe62mdnMk91jxGiXL0vRltqH79JkVZmTuaoekvejTxnD
s8vnO0dFt6MdMusttWJaywDwVkYvFpGcx9RwKNbqf6NPmIW5PMA4s8yeHJyyLVFu3kV1wNlHfZqa
YyvB5E9wa+4ZOIODlmlatxLPBDrTqFx2hTorIvkiXtlnQ8bYm09WTCShsRu1OLc3Rbj3xnsx6AAZ
nXeRTyK0Y/YBUplHzk0uTg7A8+44PIxrfk4/AX+MMISVNbFth/7n2AMOK/dxETULXUAtoIPELCwi
erFPU/FitWHojYvhX4G4xZPZ7Y2GWB3qso4OTmIKB1guLSnXSGS1fnrs1GpIWGGkDAG5wRLZiCiB
2110J2ur0RfQNw1Q+RX+5pDrfrkXxbeagJEMeo1sGXz/ZXsETobCSO9IIpxWRGAK0bTkB4PmZUh+
RN8/eI/enpCVgwnYIBvA1rM+sW74ViLDJS2PV2Ra3xcm7KclsrSgnpy/1LawHflUnH2xvrSKMbZC
hZkQKm+Th/mjpEtF424ut45E0XbhTIohbB97hjgRSVCOJRCgLNK4XSM3m71b26DS8sBT1wEF/q3P
duRJZaPXqAj0Mzi9xLs/9hAxxO7JJ+G1/N2Gsx4VC4Q7jm9Y7reH2MVi/nBr7LnytIKcv5rhJwKF
dvSjBTf5DaM8Xp7ekxxMUfo8lP++yAGPE28oLoH1OTy5hRtnzYjL5l8CrC58/EZhtRQ6BRY9sZhF
RIlCoXubLuKtSJTSYuk8OqLKeutOzaTCeOs9yfFOHB2p4DZLqC5EPLJ9tII0xS5r7dpYzLZOUcKJ
mHQJRsObws8IPQahpYYCLZGaM2oCzgd15WFMmd8pRjNUNlO3/DI90XW+T2ZLabLqtVmfYltEMntc
0F6CqXXXzdqbEhfh1DcTiLGgmeIa9T2AhwWutzPQECxQNl8G3iexC2pguBePQP8pGchzm8wtNuJn
Nwc9omaJeH8VlsFynRklq2ybvcXTegDJnyazAZ6AXCGSBzJQS4488WbpLBgcAfgscIyUnvvLcEio
J9JsMyxQcVYkan/IUs+V+2RF0I9djZdM/h1SeiaNybfDc+/TJy0cH2iaugMqUN77IcJ3myk/CiVQ
uD4qbZfFRbkahxUhbxA0uPxNNcpLmSvkgbjTlfVK/tstxT+3DaQckLdtPq8FugQa4Ya/jocmf576
qLTebFhRm+SPwr0OLUII9dUePYMEwN33zSQWcKb0MHM7NOjKreof0C6h3tJ6gNZcwVnsrPITbTZC
vu8Gv4ciX3PuT+bZGBKqEvAu8RDp1PEcpctRe3OfR7JgwLxxdsyamexufEDAt/+Ms9zTz2fYjEda
pMDv/LiGah0Kq5Eds093GxArnHWvFUuxcg1C4OPi/46/8nSIbmotoVPQ9s1mSGBiwgaabd1EmAIz
zJu3NBC635+TDWIxaT70BIyV2FyWeVmEFqiH7yoKxknbbxZqDwxtxobMoKk8mjzibeiS4Xj3bofR
WoRzBKN3au1eUCAHtP3sD6RZVq0a3mbSJkpeyLq04e3viO8R0ZFIM9cDnyk/u6yuENc9gyXiWnze
UYaKSpUTr+Xs+8LZIf6pzhRAv3TOABna4TtYeIly1ZATdAtyuHHFhI4iQBftBoPY9k4JmztSIBR9
o2YnwO3iXGrs6bHxRtb21bodTwIrL9+W9TJE7gGdaODXWN4lR8gGARJrCV0vd70qTZ+7KR+jw/FB
ICqE8qegG1HjcEWlkglr+i/GIMbVLU+ASjaJela3KkYcP25G78HHRx8VlXJdd6zhgDbiFTVoyumy
Pr2O9dSMtEt60iJAo+G85YiCaagXRLA0U9r3kUFv048KwJvHhffsHmz4udFJOSLbxPXYj1DcfS2T
JJUXAv8pPCtNFAmtUYsNeUfw7nrbNjUcggbc/rpkHzLXMFXsPmSNYIV4jG4NTFwWUGzR9s4/Ay8x
1JKzN25tZ1DOxMeRfsf4q472E4tOfY7t65ImrVZMg7eALWsH0lYmTwRX7gxtiSwhZJnWMM1+JiUx
3fsLXvMqS2WHGl1i78mLP/ozYd+nV1lulIIFsI2U4l1SYNcnOCIIJB9MNknMsIVnqO778pi9vGcc
MF9FRkLCCSfEsxuFCiaBPmRP8InxfYyjdgcWUfKU6AeGu5NBfr4NQ3kA1TG4bg/oHbAqv4Uu8p/K
5oCsq17lgPee86jHhMZWwYPTAoMh4B6VsByh1vnZYR0utteUnjpFZ4xMWCNCm1IjcRuld9eazBwL
yJJ04MQ26Iu9o8wi3OCOchS4OnVGKsnGLoSrYTf2uhXq1J7tTCrtcs4MKbZ6xEvIAcI5Ntmv+G3U
BLjZFPZGO6997D7dnaLEaZATy1YxzCFhiJv1Szlsv93if4622zgSHghV2gnV5HhR3FlGI6vF5mCV
qWyJFwy0gPcRivra9IZoOukKWwihEYT+kb4KOQlqgU3RX01pMXfhuTQkTRaUlHkwT8cfEqosHEfC
ZFqZpqDNSg8trdhtEdxknhdCn62jukcLy0T962gamA6M29tODv0ziQJ89joNfrVXTlpZGxkrpBpI
BFQTYhxlBeci/nDnb+ug5W5dQv6BDCBzok7/YG4MAqjmFKhat9wlpbBDFJjxcRd6tTy5CW3biK0h
WnKdpskhhYMYS9kHijOh0rjROrXHVi/+nFf2o3fMZN4vb+VZL2iMV4XnTZKiwA9bRrlBz/YFvy5V
uOL3JSYeyPQ0JHCd4Sq18+HQyBEQHp+Y+P/QtxsnjT71nECgNF5w9WMoz/Y1xoUjQBnAGpeHNrb+
9wzJKAyfU9ToJASGrM/mKZdKMcFX18leCALwRDPIIhJuPEevZj/yqV5j21N6j2h7tTQWPu/c3lpq
ZAIjYRVYBD4NgSZI9cxWipenbdOvF/pkSDhTywdSsANe8XUP+keuDAZPWtsBHr4+70wGFljotDCW
xY9DjHy2Y9OHLketUSx8PXH27TjT3rxrecukkFh9yxc1dxRdBmfpKU7jfhyAtMascxivlD5lPgen
jn86AgdwppGKLdCdMjYneabSBg7efTJU1UXXAZaDYf/P8k8ByZ7D63tRmaz0whsCcyBdi+osFe6o
Db4TDlgEmaavrz7Qv0l8Xeqh5dcI+i3YoStAwa4AFfqX4EGXO1V0YbxzIjAoA3hRTd/TPAwWYSHv
ntYASwFg298YhnWKxd82W1PIwR1T8c2hRxOTZmBoG1FYMjeRQwpc2/ANJ58qcA9GO+MwkcDKd6aD
Wpo7/WYU42EE7CwgXaE4oAKUczNKt6VOORZlft1Qt+ZOundHiWmY/TJRAbV4RarL7Zkf9YG7cqk7
5ZdUAcGLlAaBNvoA/z5FRxouk9RLut6vdOV6k6EDQi4Xy5c2QForak4d+pi/pt3KeSU7xze+Ss2Q
aJ+aBia5I9FQUV9ISNg0Hhvle/d+NHdPa8HvL8JxOqYeoJuYADSWNFTGgAuY5ZV/2zQblBbw7jCk
pdfP/KfLtN5KCebXgxiiOUjdoD7+X9ZFYX2yw6m/jHCYAOXZi/oIZk7OaT1hwkt09yNzZOM/XITy
g6buJKqVnl0Qb3RpZyitbdr3MvwetiW5gsBR91hwACggfBA6W3JMA4uu6irpNG5BaFskUj+A1ule
FT9UsRRgJHFfQpli3tnOd276Otq+G5DO/N853AkClTj+gp/6pP3hK1nXD8l6Gb1dm34lBfUdwjpP
QqYCVVW7FiB5yOrHFr/RxTmvy8pOvvfiMMz/P8iWKymT+YnzMb6bK6ZMvMkN4gaZx46OVp6Ke6Fp
ASMUIJb5YtOKPSFFaLywgCA+/n9Cw9bUPZOZeqr9QEXYxoflkPHUG/y+IEqGpcWzoujOF8e4ZUyK
leguv8/uv7x/93xu3wGFFGhDQAtRiaeSABgycoKjyE3HovXA7wr6RRdPRrh5qwrg44Qy5TtukTAV
KfX4ZmIkofX3xVtGJno3yPOYUnIS/faLvzZkmziIIGoUVNqNUo0J9PpppcIdQN5J+Oy2Mm17BRVQ
R/DCAwOABjR0M1sTECdYUXPKNa8rmU/lf1Mb2K5ZWrI5G+qdwqDSzCIGgKfUdZRHmOgF0SmbUJOj
orZ7YwoN7lFmca0gHTrLr+WEXrVIKw/sohM1PsifWrqhryHD9eKXz5zWyQYYQ4et7+CMUUxClhxn
zpLykCDZ3TIB/VPk/wbp80mpGKLQ3nZ11nqGq+PODPTK73jU7obBQj6lNeWABuQYp5gC8dswmKE3
/M9GDU7WFjUET98CXB4qoYmz+FlKV9lLUxNsQHgK2bqaxiKHIVg5liOz5SmV2YfmnNsXU3wkhTZk
jzL14ijFpIJ1ZEgDkY6W5ahxVk9GiYd9llwbJzOEpKFjsloRkFKZwEPCVMk32YGHQXPmj+GEC31i
kGzMDqgsQZ2PsUQKKfGowYPMMUSoUfSxKMlYzzyxX43U9nVbDQZztd7aYtNXbkmJtKgDFcrHbQql
KjRWHgSGVsDZBi/AJn+b3BMHvMa1K4uhhtPB0xFDS3Yf1BnFx3sBGbqRbCgz53AB/Ug9K91nnco6
MC1y6i4IvzEkoZ+QF011rpDqCjKLainP4TOKOUEO5+/RJnDYV21Sn1RoPTZoRFMXFXfnI11nEI27
XZzQCNB3PuhXmYEcDlOhHUkxPuN8r7pBKbjq+ORXjNZ/y9T2NeEQx8Zo8p6FeUF2R224rLmiKJz+
Z8Uyz85VoD4o7WYd6WHMoG8L62hnIKJFgYAM5uXDlS+qB3+U9DbEkqpeCgrmcBmMjtrUBoZHGDPJ
B/ZPMWRu3RCCzvcgVoCIIPmn2RT7bZ075+3BuzS/dy/hX4EXDE2VKlAT0OZWI7cS8mZDl7ygsm70
9gttdQ6QczBKyeILyqhXDS0Y5VVnUsfB/b3NVr3MmUpBxQ3bSdM7nhoPD4Er+v4NK8kBRJ79Hb1R
wpW3yr3ECOn8YvNyxakBZlnzHU2S2YN9nCiE2r9d1EC7QYjhy4cvzCmYwUAhyezr6DdQgBT23IDv
3JoQJEon7Zr8bdLEdC2zi7z1psBv8hifPpRwbEBRsXiCvrybwGWanhOmUyOozhG0XGstFwd9bTKo
a4pgVMCHRWBRNxBvFW1NW16vbq3/JJgPA9S6DzysqjPq9VoF1iBgOuEf9Vzd+oz6IytYVzH8CQYm
AV5U9r7nX84QmBoDshmexmxviHhXu4n9nI7azbgIZb9412CO50URVlPVo7Q4I3Sf6yOgiSdmQv4/
J1CfjRffHWz/D+Z2CrKCXRmq7EXWsYKhnxn6pDencdoIvkZEnjHRmGCR0O38r1VodOhrVDv+3H0d
7WsQzsuJNbOPhE9MaZm3HI9mzJ9OzLEYYJh+vGEGQ4rpcdJfBK/34ryD1rgoKrzGr2/mBzxISCgR
GZs9XCZKNW6DEGMUMQc97wn8S9PvwxLHu6RSEoJnG43tk54/kZQon2xNkrUIdzk370tDl17LdVBv
kdc+AeXdhf01XbGeUBu+nC3/Iif7WqCHw5X7oRf+4Qg3Hmla5B54dw1tskYJDfybivT8UoQY7nHb
Z61b/JNqHbZUK/zc86T0T+AMEW0tAcaI7rSIMqjTQFfHtM/IIs0hp5IITsGCbeY5BPbHm9TAutKY
e2Jc/xpTNu2LL1mNTOy26M4WFO5W93oCHQHCTCpa/D393TKOZupfVnknxObux+AAgl7p1BbFvqrf
B5Xtej1RdKSUNxmPkrAZg8fYTN61OcTap7/xSqQX5gkdQ8EWYFvJZm8QC1CZ2vS5+ozrRvcM5EbK
KVB5GAnz4Mzi7UPhhkAnKCUJvVpVVj44Bx7jBT1XtOxf4/GCZQw1uPlpX4aodcvqwieROa/mGXDC
HdnPKDOdMPBxgfgU0BL3HLqrMJdC8tmI84CWZEVC/gaYlso6yep3yYi11zPD/Jwdu8K8yPHApLWQ
JLrJcj2LXoPPs2z65/SQLbGjWHDAjf/z/c9phhf5ws9j2PXSXxNWYzndEpfOuoAOqk5nv4cyw+VB
GuU+ZhJFeMa4TXDJCxWBco1UMZZPOCnvQK/EcSEgX3Zj+i0RVWlf/NjEcdlBCtPlgnjYXGhRu8O+
wSLFbDoqBNbqEpJAZeBFfODpY6LUfq81ShUz9YJ5L7PzUHjup2NC7VUtE2ioJMzsKHcEdTQAxFhF
K2S95szvaIQwJwvqj9+BU5ir/cLt4gulgdH0JPWZfLGK+uYLU/6T3KTiDestnlw2l4t1z2zsURuN
ea/qqflZB4R+btD58guiNmJMHr8b5ny+qE/JRaDv03BiJnwoeXtIfHAKjAmCchBHEzPHzQiXfJp8
EA/RRNhpYvVMakfivaN8lA5ErU+eiWCUcIKfPU2I7QjQtfxNVrbE6+E4EfKzulkMvn5S8G9XWd8L
5lOU9wQ9QS82NKRctXXNit+4jA1ZJrymZIZlHAWGTPuBDmzilXKOny14hZiklmjtuZuUfxO9dGYp
vGR19NNNr83B1SiLFIP7DaXtcqLr3ySV8eTz2MTJosNpOXaEmfonzprG0d26W87OHVsETfflqg+8
rHbowP2nx5KMKRuPGFYVg1Wq8Da0eexTsGjPLU2So5l2ZqsO0oEqcd6obgdJIHtpZ0zADsx0brbr
Wf5uNAK9d8ipUIGCR5CK6KFN5upOj9FTGFu3/jAf243nVhKpEwEScD3qFurTDsxK7Ccv/YtoCMBH
rzTC9ZE+q8BfC0HveEyR9JQQhONmvB/haT3QVBVvKLc5ZpARVCUEWQiz6tL39Un36yLuGeEwN6IQ
2fck5DfFu2tqLQfZQeI2nGpVCev2CvhBK+h9M5fKPyQ4vS3xdlU8S5oP49eMQOFMNpjtUYqoWjbF
CKkaQYLmmMZFmKT2Lkt7I0dPcXWXr1vB9kpsBCuamOlhJMNg3hh9bmjBS4FXq+IC59gL8NQm0M+v
hIqRHKGRg429HApiw+lcdz0VGw1cGVV46FbCgaYGXiPc6qkLZDKepLWm6rme4gMsgIAzQ4nCVWNs
9Le6u5ip9BeUB1jfNqC7DVa1TiL/q6vSZXoMWWm3fSl9xtBP0iVMlu8KyoF7XKAw4gamTZmZ3Jv4
n+Jnnph2C62iiXP08QZ8vRznvmaVO0hykdW34tF7sjk59b+gyfylQbRqoNWtbJUE02rDiXus/s6o
SQ8xpfptbdjI/v5a00NO6Wq+LwFT8WhP/sYo26d+K3M4N5+jUXW2LcccYM4dIBOKCnWyvPJaHhf/
AwsBMJRAAjtV1V7ouaMGH+exVt2K0uBHYuO/SR6hY781gAfGJzQqrvZvyR2u0SRbJm9hTL4ojdvI
lMg97h1OyKfcNAJP1U3f7DwDHNiFh/Ei6Jg+3OFFcABcdzr2pVxTpF7xqdOVnUFll9iH1eLyMJbY
zToeMMfeWCaBxwaLUpYLUzFWE/0r20471XAcBQCLyzx1w9obF4dsk59N2h6QQTPZXcolVN8Jxvsr
qf0GHg79SRgv2ewTNte275/o3HQ8ZWBEhgkAg2VZ7tizWqgpo/T/4MG1K2KndU7xD548lpDRIo6q
F0XPYgyrf/plAxgk3pVJusATIQfaVSpU6arnfNtySNsBqeT+RFXgRJJAmGmDtF06mnVNjnjFyxw+
g3dzVa3mY/XhQLu6JVnVo/ymuNMwMVyUnK0oizz1QiMS5vlLfz4P3XwZU9SrpB7grcic46Hk/KX0
uLTxeml5jI2AOay3RYGvDNOLlAlRgIerhc5lGF7h7lu9g+EMQ5dfmt4wa5z3giU+To2QuQ0ajIWx
7pgGziZqz51qxFK4gB+L3PKlEKZSAs3blGg1dtlSOJVv0bBdT+hQAHT0Gmzn+kgKfk8Qw8nvnS2C
/l7z9hFP7GiMq8tIVE5repQJmxgqANJq4CR7lZI4EXeLN+bq1ssgob52gy3lXQYZW/yiURX6pCVm
P2g8AzLsyMTAQXR5+YZmoy7I/xvYKrPVKjQ+6hESldqQWtdLHEcn59QO5ilrHRigSPtJFamIeRSX
XJnnM3WJeR+i2uI0S7GnfBFql3Z54Zsw8RRwwb+BOSWRVKn4n/dekWReBiZ1vgMrhO0l5xGuuODu
IuZR+ZncvT+o58kd7zXL4VUVTwsuOIE7suYIuJJH4g/PTOgMeX7HQtnZ/auY/kpCYOWoAH4cPPqA
x+idDaxzI/zhggxxBpKWcgC4ZUZ9bC+J8+tlUro2FsoklQ9rpybBV1bIsGg7ge8naIgDmL0Ykfgf
lm+6Ry+TrvHQUJsX4BxER03W5lu2MM3MFf/l6g1/IqEsNYbJQS8QPnIqipMrHiRojEF4aoEe4msK
uxDUgT3V3RlD2H+t4b+vGCYRx/8cWySG97xLP11W+TSbONIafZKj//TI9Mq+Qbr63Q+QxLN6Q/fs
JSq3Qx7LI9619EZOggldjO5OcETXmUjTtAFg5IjikRMq9OmVnaTZzWiz7pIL4jS9CIG2+6uDjBGc
tmPVaC4jtckmeacYOKbPuGkX1oOuFoa9vvdYSzWSzT1eLj4jIEfblNbsSPqWihT/xIj6aAa2WrZ8
3OPQZypEAEumQZcaBcJBQ/GXnxvJHbuiqVx/nQZ6ESERigwv4pG31S//VHgAqjUVvmhK2L5zcAbU
TMpaQhZHJSN5HDuNbGQ5Is7x81/txGfzTmHmk6kSGk335eFO3zuzv964sZHa6LWS0MTAwxP30mlb
5GOjxNNNuFtdwXM5zJ7L0McfSLlFU6nEiL0wAPOifL+fRU7lu75844IIg/RqCrxbW3esucRNVGXm
fhese2UoZhx2i1Ivq8hXwtf10X/nJrhxPDvfhgwJ59X1Kzb6mJJQZ2s459J4KBgbPA1XD99/co/a
H77ZNZpxYJxVxlyrmeYWwEBzJEGb2VjJKjRh/i00u9aJi8YIffAAWB6vqnb6unkQ/Wd9jc64HMDr
1Q95p/dNUUeRBvyyXaX9Rk1tUlfeKpdwDlXvmIVEyIToMtiDB3++K5vDQMZ2ZqKjSp+S/eWX1Z6h
eRyhi5X8xzFAK9CPjlxip6SYQfWDjPPuQZsK2QQqf2kYVVgacyWNRMx74DTH0tvpoKpqxGhhHCEA
kejCQtNS8kCYsijGzzRDE4SJorMnvcIeeH/uFAv4qZFI0cRkCZTUW5kuLSvHJ7yRGDrule92ugzn
LQgi6q/+GZxLIuLEEXtRsCp0uE9eedZH8Y0+nps3IMAt2/DkZ4q4dKBxb87Z+TsfEPKp+Qn6ZM38
3CC/QtBIo3TKoL2Nsrh5nIIQMxH6WBi1y3545tTpUd/HcYYz5kLk4wdeKBQqQgf53E1SbzzZrfdW
pONbFibj4o3978s5aR3KAgeJvDYToBNno/0BjT89yECxHts1NmhhALcV6Zfe2rqcohdXMU2iM5fy
Kov2sEFqiwmmwFzjbFOIbErDH9z18LVum/1s1RQFXMjDhPYcUWC68wlvDZx9hSlC2YTCR9Pq0COJ
qm4Rf4c0V+dwRfdMb0KGjRsgkfX+R1JXvy0TO+dzhyrCrANssSZUHndtXF83839iTRzGKCsy6512
39A2AQ+FIzz7Oi3WW6F+FpWIJ513rzTH1HwFOGEs4g6PCPaZWrJJlLiVFCx7eNps/QYwghymW2aS
GbfQ4z+rm95WuQBytyGm9rMXTeRCzOIqklU3SC1XuRbpRRtE9IiqkEsB2uwSPTRjq4QegIN+Zr/B
6JTgmBGap2W34xa+fh7DZYVtPc3pkA9171CNWJtAn9FmVN/vkwG3nMQrX7lOT5Jz2OCobcFpaSAe
HzZe8vi3a99UE73qoa9OqptM7AhHOtWRD14XCIR/oE9rjqpD6RqfxCFnh7d8iVXB26NsUcQcF9D7
wGfgVSUfznCeRHwX8a4heLYceN0YdCbBTxjRafTQUMcSP+VPBhUEm461HC08QiIbnJkoYNzw3cTc
yNAP48cBIauVWSjRnGMi716C3A4ZStqjogCNnwT+Ma3Jtxy5VtSAUHUCSiSKnwWsOpsbNoJ6Fp5J
KqIfbGrV4obzqJE8hxRmlwGesUjJyXKoBMyOyHyvqG0LgD0nYXaN7mJM+yOTvmdq5p6tc+PkMlGL
5IdC8QwNmEtL7/kbJ6kb3/XH8f6JYViliiXlDn/q9AlH7sa8veYV9bs1ZseLnH/oMhqMV5QOSqUJ
WqOQD8cLBYh2SOAjnXJzWh1u9XhBXJrNhpTfd2uNrroczqJSAbCuIPA52eIneP505J/dLAmE4jfy
0c3dwnn2IxEEVxpd7EVIcVCGQj80a9qTrv7gFhva68MLH5XX+eIufWwpG7nylL2QA41McNj2m8H7
aB0lNEexrzMTKVdv6uh8w505pbwtZDFxKSakBmqQ00vAZk60yQ7YQmyRN8b91oXdI6XpAMPcA/g3
qNlGTlAu+uKjB0ski2z2fj27c9S1hqnRx5TvvRzp8rfg9djKOjv7IMNmA9jONIBQWr/ejeudrrCN
/y2xQ2yyO2B1uTfwyGZt/eYD5/xRefU/lDTCLMB/htsxll52VuJJNy1TdKEjfqfcYsv/wU8fVKmO
3tzv9lvxhzjXZ1ouDdcPpwJ1RbkTLTo2PEXIE1CKgSlWJCHDC3JF1jNPcW3yEzGiWxULWdKl/Eb0
CMICqpZCmSh12e9jKYIHA8bbYFALW5/GmIKEl3F1h4Szs/C95loU4ilBDj59hPIXg2wMBCjwsiic
XuFHnW/ncnYeToj6fdMUg4qJ/dT3P0QNdJCNwVHMXQIBC5qASu6Wkb1bNHw5+lSZvQVvjK7dKJqE
10Xb45sJjmXBLuZl+/6grMYusf4mm0b8c2y4VMmCjkKFfgsYwR6Thvxgi0+xzeZ4ES/VlL+VFDuv
GpFtFrF5QexRBG1OX0TdRZZcGHwAaCNTw5nUv1bAfUJKuNuQROOHnkyI10MxkXVxFB1/2sT4wahk
05I0eG/wRedMa56dGUuKE5Y4Szya66jg2DCcq5BmbVT5iA5hqdVT7Tnm4DeJ0Rq2ls3UchjNOqys
amqD+PRcC598wPEeSn2K2iX7NGlnmoIIfHbOaQCEnl/i5ORxLbdVJxEX+mnmEuAm72t4Q9qJ41Ee
crVbPDsMJHUKZ37O8aZc0EuupUufMd8/1mketKTAYnRrWDIvOy5prniZ7Tn5OmdlWbNYGdMyqABA
PrWT8rP3DsseLJEqG0iDfOe9d42MyiwdzXp5/SftLzGBe5N4/pyPJhPrCkOA6TxjG6AQr/RybhCf
DRlE9jtweM8N7iurBjKuR6iQAQupO0vFg5O5xL8akbUhdAYzhyno19jq4UaAC82CfeHzmkR6iHqF
xSrNUot650fNkzJyD1Jh0D/nKvYnGXkaOR6ra+ZTuMuuSm9rGfRxsXHqvVaSRJonhe24LtKhHCAM
9MlzA017mgV2+JrFwK7dMBzsR9QI895NCNnjzaXItZLSO3jxo3gqb5y1J3LjWfm8Yr2mkR8LjMAF
iZ6yvhRdYbE/sMBJTeBEczDqvvUS6eKjRRmXiyB7uIboVrk+EHjfrQ/BRxb1eFoQppjyFLt42aQM
byfLR0nRTuFcjM2IhYOMMqIOu4T0Mjlr5jbnuhVV2URZm9ACVN1auYUrf0YmdfTiGyfqP0XK+HtB
E37DCUfd+A0VqHAfWp3Nt+STLjHJfA4csZt51IusnbDqLx1baX+sDraTPc0WnQhpRNXt/RkTCOCI
Yx7Ix8nfivPs5Ds+ViaqqDsyepQ8Pl6bzoP9O2HO7ntjDUz05FzTHCMSo6ubZDxrjqG6JFvTZPtF
hpOwA+E4ZPlQKx4dhCvz5gJdDwqY0Nwy/9fi9d/1j8vW5H9clXiRtJmKsUlYq/IHD4NBO5q1xUnD
M1IiDksp14Y24lhtD6iaSOGWH1D/1Q5qGMUJbF+Qs7Q0WI6m+11UTjEYa6wGeuL5HcZLcztGlyyn
GmJSgPRshHj0e8fMpi0aazLEY+UUu27HSgn9QR1Jx7qDu8On//hhEepkOsZfNlCtXCsL30B7J9rD
Qr1C4dmCNTj2E7IutEY5bn4d16A8wdRVUDgnHEoOQxUBSx+PrM1AGnSSh39MVX5IocdcY1klxylM
jIHL+JDtqRqfLl4daJdqNvAzC82AHcMv+zUob4m2QXQwISeGN88yFSWk0UwlpTx8K+yoG5u2F8EJ
XQJshsVM3+KxMgzW+Ib2ycesGu+OMqsfm+oU0TxogBpvpY/976vdMUIjIEQxPOequKkzreWu331N
WhNsiCcS9EaEq7hUP8v85649gAQYp0LCaaug+chx8V+THZfo4z8s9aTvAZzAjBXejV/iiornp7Uq
s2lS/ZnCUKgxu6sD8LhaQd1AZo/3MmtOXekSVJasHAlAw7oKSs9EikCNQvEWxMjZey4KT8bwsxVX
7UYgBTOzp38R62aiGOcsf8JotsCS8y00Ig240wtQo9S77Lgp//9Zlp2C2jYDsGkcwZd6AxbJXXtP
kMmokDDSBV6uEfr3t4sErUWUK9eeBMNXSbbCFT43FzgRKFsVTycJg+D+E767yOKbiZHUq2r/TjmT
aaT+CBRm9TTiD6hXyfs7zLTLB7IOSo1xJxbvShfOIfP4ZfOIZSLRQOjSLzy9t7b4OuxmvwLYVkaP
qzLHzyZIVgqVcIwNhqTWdXitO3ZBgcIko5LApuUFR89wU6dSL8XX1kIQkjgKg580QgrvYcwGeYyJ
EgDcAzPvLflxi+RkCTwkvtzt2kTXgdHpd/9OCHQqtNUEWWjJmPBgdLSRWRCKEHRsZntVWHf1YwLF
70DVpH0Q9xUXcYIq9MJR/WA6C31JwZj3x3Rv2YY44ny1R9jsOprKmXq+LNaCj7fTAtpbnQ65tF+L
nfXTgtGB9mqflCQaR8q9G3VVty1Bel2MFN7CMKZ7OQ7mdV+WkbE2dCD4bp3mXuFetLNimgOXLuyK
hjysG57eDlvk4w3Cohp0gQA1xiu5DcqXx9dkTZZXu/kgbRs81gGaCc/+/l6D4ubsruM1RKQ2+uoI
idvfwKW/Jd/hTojZkOTd30y6WMCx6Z3GF4E2ovh7i886n2OM2sd4o78SQqwFo4BWr+PHXKZn0jmy
Pt4JIZDfEi9D46VP1rZo8gXYQcd0M8wdwHLPiMMZklBKwvIXVrMoqOYh5B2O59RjMa2c7dWxcmZ/
5E8Z+/dgd8r2/DPQuhXP0ljDlGYmuGuvk4yyHHUQUY8tV44nfPyZze7kMeOk2BedwDF4PZtErK58
7+ZDYEAQHCAK193iVyOFJvSlnfv2HxtDkmaSeFiimxiuEnlc/nk+krn7IA6wQ/9HVsWkoFwKVgZn
oo148+v74NMKKYRM17UZDbov25p0Y9RiWELj9FQQJpuAlwxnLSPVtVfLwp3aE3IYKfYVa3s01Lzl
+fGWkbhOQhPcKtVRtEsCCA1pS6VwxcUfhffjgH22CwWra+GiwZIPytnlanleNmGr0iUjQUyoWgQG
Yy/Z3SknkA66XA3feOpiKD0C/9QPFOT0N/87CTxodbySKXmH6hzu+ygsfKK6gfEn9jYgLeE92tRa
RRDPC41H+Sd2gxOPVEXNiOURf6tCrF5sxfo76x4oN8tFCrBa+YvcU10KV71hXebweEW0UBCQ/Aw+
kCxMP2ikBDG2UQ8PPl87Y+g61j8piwSD/v2kKtRyJFn9fwdkS7TWpdTNXg4za7v/idKxLmpb5mD8
yy4o4x+Z7Hgp/5vaiYfU/Z4bmhkDx4naNpYH0D6hU7/7khdN2ySNmVz4Eq4bsjPFumQwNKGi/Ntm
TDuVwOZ7BTvpPG2SXhYkRXAxJpYvLOnX3iJncgZKAb1ky2TGT9iNFO2/O4D+bu0KTf6stzq1zpd4
MkGTjLDtMe+03IcOJNTh9Z0IQ6UD21RK8DrR8OMQoXTxEiERACHN5ePlxPsM7rZ651RP5GcPQgAF
FCKw5Obfqzo2fFeXXnAwnYMxQH6gQG/pngyfN9Nx9DLNuBrpbGXMFVr3KMZb9xqkbDk8/LgjFYVB
QNT5252WQc74mXoSjTninHDgBah/rZpC4GyhcFoTOWfVREyb9dkV76QI4Iuwo1hyCazELwXKjKLQ
D20loe+UoDON1+tdOAoqtqJR5HJCjF9RFb4yd2ZGdUjcVtLJgbwzrHGpmEPtiBQMUf5lrmDYP/TP
M1reyDKBnhL2YhcLuGGGiI8mFBn9QM1S+oIEhynLkbl9krT0kKLJV8jEPFhrLLGwP1T6N+st57Sf
voGh41as/uFuVcB7NC0QtDMfp6FNy6MJ/pX0YQ6dVwfXJLNHaK9rVlhas36jL+f1v/AQ+zMlV8pI
2WGHNz1vjyWDeFqNGJqFY6Jc4ifrDgLAlaAAM06Pq+00NB26BbvLikzehEIhOEfW+3Rd+xZykRtz
uT4fbSXKtJtTLuMQvpc7BfIKqda19BC4HwZF6uKnKOCe4ADuBsIQEhEMJW435WVkVlO/h3OnvAs0
S3GL4kjku6Ed63peAw6PJk2vNQq8mB2cXQdmyQi8n1wge2kmGrYB5o9HRbFWQVTAEdgCXflTF8Al
00+VSdLD4+puUMyqts9hXSEGuIWeozXCWOl/tzpN84gEsFhygxwV8J07gFYkzPs9soRq89P4ew6c
A41ON9pfq3XJiFm0uI/PmZsKxCoikdBe96WV06X5kVChDhmjYaC/Il6hb3ukTbo3LL07hNM2Kz2K
vnaxuLLkGkuFUCTusmZaGN3U3d+Wx97ROWQkgRIk35YalvAdzK6/gQN+GAPgqpJpipOLxb3KFqb4
2Z6xGoi4RpCj8MeJABWjwXDWzHzX9mnoSaq9i2TLcboz8ZXyd9xnPg8UC3lKD4/pLSnjJ1X/D78c
BRz0pbx+HMcUu3Wv8d3mDPgqs4LmBPp8K+VyzY7ayuXXbaiCiBS5KNKloijIN2HpaQJ0ZVF+L5c5
M2Xg1rmys1Fm1t3U6KZnPui9TQJKt7WhCgjfdxExu88oqYsbWklxfAT884hwSDmL8OEnv8m02GmO
w4GuAz4C4slF8/8ImHTtyFNEeLAY5O/DnXvK4v0vXJrsGXH9meZB0TbJnlUuPj1rzVIyZVS8q4gx
eYPNKwvJmeeXDuuiqcOfVBIxEwa1xMOGjuXKq/Q+w8NQ1z3Fu+k4h1RAD9YF6Y/+WguFQ44pj90M
eTvIIfClifZyFY3+Z5xrxf5R6QMtyE73I+a1bI2bfbSaMkmp89Dd+sd7t3/Cr1WzdwduRJmTPd7/
BacU1V9nl8xHe4XKXBApYSWotbpz2e4aa6763YOsxyFGbwMsv5l91RcpBqSL5rt4u5EPyoUMyIAl
JMEufrLe0ibxdskywR67eQH/prSv8NG18G4jAueNe0URKBdeUbDY48OcxP6BqxEWqZ7lPCHHzlvf
5dL4doYP4ZVWg3JyGiXtteuVEGs39Ex+5884TDTeR8QnWD/IYqCP2vEzoXIblDrRHF84K0IRYH7r
vZVeiELnH3UEIicANJbOsw27+67ndAyHtT/KUiLDKl4NWRjtnB2OJZRyN6vYsVH+TNmKWxKTAwNV
rb1te9/ySq+7WpIUgPgVvrHnRnDMI7CwJb4/j+z3EkPHxq7+Ux611LaVkigb34KB7dz5JjigH+5V
pE0yl1VOe5e4DfLJ0/5L49PUdNp+aPNza93zjumqu+ixN1PVQPPR1yWu7fK08S8XhWDGLgh0L84g
hwDxm+PQLtkd3vbtnBRIC2W4hwPvpwhkEh4RYhBI7kWMbDrp6q8fA338Dmj51Bw1QhcSA76vITWy
T3JRctl2PyYo+EhsFGyenG9NJCIxdX8ASOsKQCmUGuOBykq2xjxZhY5Rgi6bVzmqDyxMDjmj5/5Q
e6vDgKOEghet3hcUf13s//r/RkrwOw22taL+b0NqS2dMhpkxa5JilfZpKIKKBFhNVk152GMVdglS
mjhv8dRespk3nYaA+f9o+b7XISPlphpq5wb0LwsDcYDcBAZPpk8FAZmwBUNRDFyWpDOWWuHMCzes
zzwCqp0QO0Do3tp4vtLoouyB3Ww+6WeippBOCbH/JB4k5/dzKqGn9mMx3HotVpPYqfHZgsfCdGGY
U5qFrJMP3dWW5WuHfN95S3wGyKuMgnowh7Ey6Gxi0tpegVhSuXsTykKPPlKyTLNuWzoZRp1HtTku
SxNTKMf8GFbURR7mIFe65bd82/+GCLjfeDb6/iHLTXDDxZiDLMXbHNsxUHZ0VGDrGlGACqdOdaIb
KpMMn/cz3GMA1t9asuWbL+IN14tifAicRWrWwVRxi1bwpEE4D+QG2msAUktpMnNbPqu4c3Z7QSIy
ppaq1TSiWxdTXsrQNLaOATpdcObEwJJ2hH55/K6kt31HNP9oifSQQ0M9gOkPQqkK89F/NY7E8+r9
8K+c8IX+HlUdzTVH9BB3IbtDtyaA//60Wez6o9jd2iWInrcSHr1avKxaPOK1FXOm5j39gn9K1vmu
FH9Ow00uhOQDjRPSpXlEr1GRhbJ3gljNRwgQ1qKjElbLdRCOszoozVVvRw56+Yma9fALhnzuWQJC
3Rxe1Mmu5SWp2XnuLFfOD5HuqbMcJ/Gq3m9Y6jG9Ke3QzCscTt54jqIBXX0Bzovg0BFYXWmgBfYr
lXIcQfV0bUFXIBUVvTPBNVqoE3nsaLGKGaiWZs6AK4J69iCnQ/XO9rKpNUZfnDTwFIyD0Q0SDeog
sL5ZG8oxQEBsQ9/RamN1KdztXNXCn3pje8dzQRL24G2zRIMN8TwSDxpc28Lw/JDnb9dHLsHHhhae
X4h0fzk5iSTamj1shiysfgCPiHM6Mve8LQTMsnd8FTJsjUL+xSja4Dvd1meIcXgMtjyUQcKRemhi
KjYiuXDQ85aQPQyXK+n9wUa56K4PJ/fE+uoo7bfRT238F3GuK9iFK7X64IqzTqdw9ShUrfuzZBVg
WSS2ZNCdcwAbwfK3XJ5wnfsrGnFcSGPUaVH2YChfVmV5Y53qKq2MYC2qTmA5uIhbPBTO6PQwqCOQ
PRCI8jTdj2cyRhb2XGM+lKJQjzw2xpSfHknL6H5SOi+mWABIRjxwnTQ/MokQq4VOlJu0A4JcjOdj
Ut7CRO0Ery5FF28m5bc3s5SMNn9nm6edLLOwnJ1XZgEB0TX038CJH9S3eMXZg9WnF0088tkRzHrx
fEvR7JZ83StIwWifKObLxempqpGgn6Huj9mkWS1QNRUMhjYevvejf0zbnDXLn1IbKJV5DLbbxoxm
a8Kn6mfVgkq4F6mthqx3njnoJHRuR/1KAv5ijC6g2CrhpQefGQixt6Gqwa30QZGxjWcMay8EAkj3
8FqAveFVWB4v/ZH+tynjyn/eqM3uBT4vLVBmeDyGuhEYBsLve6+tLoAO7F/k3hpwPD+FCdWfJakr
31sCGUVdBjJXwSaHiaDHGFvER4/mPsKP48QawBE6Eq1zQRuT3fzJheBKJKFVTd2yKUpLhjpEZL5S
B2Hho9+PX77RYFl2twL3xLS0dyRulQuf/kEhjAjiz4KNeIGwIyzTCEVQxJaEK8Xtaw8gGMfqufW1
55ziM+VFDGRO8FHOXHX9CKug2mCxRLjYxvzHDVyFEghp0Ofjfnd9/rGyE991RW0xJbz3WAml3Zu+
axQ5/mdK/arIr3ysRUjL+23Sc+BrkFihMUNel50yqtdKroZ0UoF1lElqNAu6F35ep8bNiU5IO1ah
rZGqrG5/351i98cInbsHJ6gDCDctn27+H6nRdTZqcrauDH297xhd9u0v7S4KF5BK6mMgRRftkT8A
RSLhhq2q9gPq2KInAHEGCoVvBANN4C12pvYw20zSrYvmWTsIgJRIeJUkqO4RdJVpLSjs2VAKl/dp
4BzhQ2CTHzxQC8vV7S5eFBM6VP7PNa8PYhP9zihHXVjlwTYow6yHapW2ijrOwSOka0Oh4K57j9xk
1o3AC+qpNZEsSzTaaXDFOmagqBRCp5A8nRFkxBhoGTs9rP3NJlK8Vg2tUfSkxtiLqQVKkEW8BN5f
/jqI/OJvNcg0LUS7251Bplswwk3Pr+QkwADWcF3dXBqRBhiP0FeJ1g6TsFOVqeXz69NAXTM4zJgn
dkNqphbDy8NGe0i4cqhyP6ujH9okld4IZ6UD4EEvKgXjqt8YN52R3mHnBu5nZ9c4QB/9Sy0r2+nl
hu/wUscEyWMbLhIb2b590dNh88CdHXkIUdiygWwgDG+xWQUuBcVq9seDBBiDGPJikV6Cxxn9aco1
+Yg3iwDN22UKctKY2Os6qWKjxT4CxdamI20E3yDJnOTrICl/2lB4eh3jhvAu09JdGx5rOPpu7s0u
vjRVn5ehcH02OWCAOU5sms1yXwi0DW1M1js0LVe7Urz7i9mtXyYONJLUjie+Hae3+s+cTyq+2fm1
Lqal8fE54prdwHQCVuUk3Zl+vWsNW8kZrpBu2eeeEaIwvcRZJE4Er+VOJp47P8+9xx4LX4EG9ytw
fQZFV9dlk8YTQgZPHoHIaivxkCZw+2wV6qnofURgQRM5qK865P8B/YLlQP+16fn0oU5+uczLiLVw
Kck3sVe8Hlt6+fmz622/RfzdoA3AZmevX329/YAFdYrzYCgUy64hI6QbUjH69kZT9oZG8U5u6vfK
LcbzEiagpVwMhK3MPjefTyyw35tPdc17L3iqqKzPiszta/inzfIGyXFA2dq6mgQKIZaN1C7gI0Jf
Sx0/+O1YgBniWGbTQrtG23t+mZwmaRsdhAxfpXf5wOmpG23GomAA4DuaC7zseSgvOD8bfwdRB9nD
DN7nBxMblQ4JZQznFFw94TFNR0m7TK4o/R7G6Q6cDWmyxqEz0fGkYHHbjfYXOwLMeTeoplxk726E
mI4OP/DtOSUAVubvZ6WBXMU8sZ0SUoPi3oJin9Gf/niDMBCqIaUHG0gZMyF/2zKiNgtTVOql2lOR
uBGFf6ArgjTe3Lik2+7Zt1X8NNNDQFikbvPmy72rKjGcJ9IscsvyLVwgoHRge5g0oEaqzvkWy+DX
okimWkrDb9Y/zywwfCUxvNbIlXzxTNNkhN89OtKjJo9iz/enuQjAO6wZfYawVjrZi0PtSJeFZTaZ
st4pNGT+g7jsG/PGLC4Js6Ax4YAtlU0AeM6iA+lvLjrcf/7hcWwhGn8MwbX/RNY+udekshLQSG0h
K5cJ4/P1Q/0IK+ytfiTHon/T3Lj45Kmy8aG2zu35zuZ+nd0xscC1nRQZi0lYzOqdaeDNE2V47q9G
kUjSP2ZdZ8T18+4kX5VzlP+fwq5UV7MV/z2GSnDSSlB6fWFVze67IJpPVL/1opkeUOE/wQCE81hv
seu/NIl9TCNMIMWB/gt/vajhgXlYKLaqB1Tj99qiyj9ACT9VnO0tw3CGXIkfHgSgL8iiWISSYWFF
5BCPAzrzJVmVlGsvDS8u68pxSeh7xBs1tx1JOsbOVKT130ARBQJoHgMi2PmuTGwHG+kwY9+Eo+iv
BxgbPHyqGVNnjRum1031xiKidcM3DSpO0GdqlIGmHNkMg1sUoMTp9Z+hXQ2OC9jlmaxJASceiKiq
JypYG1o+vOO/32nU6ARKrxNMqeU8y/KZwOnhvilZeJSgMJbOtSBwZ0kKIXbUqjsX+ek/lqHGtZPY
JFjHd9XANH49D2zCrT7pxZW59MvUlg5Mfn3KYYvhXAHTSxgZiYik59XwsGXQ2rtjHELTm2EIkCms
A775v599gBgP1mKlYp4byPPAIcFNSXhyKh19mtx3HFETC3b6bTz1p7tMzfZ9bzh20j7xHTX2ceNT
y2PkONyNFV54+WiDUu+guAB21p09b+97SbgsxrZy//j8/eX/lBG1cc3mp47rEeFXqKPIndrMbxZG
X2F9wMwVi+TB58WpoysyMAt9lR3pCGyeeXF5yFFLNDgz0XFqoxvrvs1MPhQLGnFPhd/3gFO0Ix0B
fzuTwnrzVJlSUYDAhtlXcvjex5OB/sRQ0yKNqf0BQV1GVMdvvUWhpEbgtFidT41bgFx6st3rve5C
m5EF9MQknC6psr4t+htnI0MuHFETIZN+f7SFcDnk7NhYLSZdM6PDf3XLLsRL0zNF4Ivaneyt9dMu
H0FFfeTXcQl1trhNq+JSo5udTkjqi+p31Zszb+9RAaSQbvw3oILqCxjEVL2CkPyoyzR4/oqbSp8w
qGWZI0c/E34GaVj6zPsFimYBkfPccjr/Ct5XW/aP4XbOc/t156lHOODGkvlpzgo49VJq2n4WkuRl
Xt7tiF/BPoGaec6nIW8V2nNCw3o0bFonlk2p5Jr7Q37fzsnzEJs7vOMYEZiytjHZidZ9bEDHb36x
zHzyccLqcko7hPVfNuZ6Sjer8G5RL3rWjpWdaBvU2LE4gArIko6spa5GYXxAxWS9Quxoae4txcmB
50DnKidp5gqccQxvPDXH+4NbZvXlmTddUVt6T1La5mhztiOJFJINDmPuP3ccLvQOAISmekz2D1Jn
Hw6onD5wDC7k9eQ/SIWhJEyQ9DWgZC7RCxAce2893A0FoaWjcytrZS05ZcteRbMUYPGQKgl8rd0v
AuXAf+kJeuEa/yYOvaVafxhoFXM8rF++w5AzenQ1w22xaEkgC35WrBndvRwr7dl7HPCNq6F14455
i6aPS033IZl77KILr+kZrugCS5im704WGf8DbL4od9zcDJtruq6Jrv+iJHh4vd9/uqlXMoM3DCRM
/x+4SW9WGhJhJJs8COuGrKljAylEiM4xw7p/w67FQ3CcYCn3WxZKo9bPOxj47NfeLz9haD6u/6Up
BZzKQzYuBcxryHaNMiUJ1k75zOTPCJIrJzGO5L3pxAiO9dMSC5l0cRnBr9g9psf6lpWm2wr47eYT
HUqxAzDShbQznU6KaVLfbGrNj4vJZ61dMm+Gi6x2iR7rmI3rs+Z3tOhUitvU34x4BxqxAY6QDhVx
hB4ZOSLRJmLUFCQTY8+o7Hgjucy0KHw07nnmhQIJ/B4P0X/cLkQSsYVRwMUvEVVFzwofarFS5yf8
0SkLF57UFSE5Sy2sDC7QZIVJ3Egu2VXPGD88oqjZOKIvczzzrTtmW3dHcujvk3JT2dY62TZLPmzk
l/GHT3eHudKg0ygUIwNOLAf+3QBXUaSRRIfyOK2LDabfhxbAIWjb0X7R0PaSiPhgip7tO5OqIB2D
gH6ffLbubSqKlk2HybNxi2JEg0UL79g/QfCgi3pm/ItTz8iNFe/DArit31Ix8daFKHUyHMBN5Gk6
f7N3qqt5abo+m78Qh6xCC6gClvPlSiWr/+DH5oaI3vDAoAs9AYVCSMQJWrwYTXIyNuXUC8mmMuED
PZvhMVyO7pHMQVVVH1NFBbtKIkC8jzNd1m8wM64Pt2LpIrI2QGnipbhwArd6KjBweuJl1lEdr7C2
jsw3B9zDKBLSyTkj7yqavULcP1JPMDFbyilPftQ+xt2rF5zubsYatFBrYdjowAwOsBCGA4c/SWcD
KaykSGWzzmEWdcjPJaOfhk8cE77i8kGaE/vfK2QPLg1qI6PbfJHSv7HyaZwnSMQo8FfxTNwWUvdQ
XR4red9H1eHVhvv7k19ihdVk6pkh6zZznCF/FiD1x4pxIfyCMHk85yxXnw2A7COfNxKn0bpwsrPR
H2zzdIf7duSPYxQ3HFAbQIO9DZEK2eOQNfQfrWpGE59rX8WRN0+Z2V5nvfpQsEuyqEregyERqK7i
WLCd0X66yFKDv5up3VxP8Y75d8X4n7Wo05Pzi/CwfmrLC65s2ahhupRjiMgXSXC9t2x87njL6yUM
WKYCtypx+ASHqr6TbntN/VKarwr14VZeLxnxFh+faqhsMMQUUXWWBCfHrECUCxk8SS0dMes0gmtN
sH/HqC+0AUaSQOlqIS1CTzkjZT3UJmerw5KBl1NsyN5QcFBn8Y5SCjo4Ms4lpskudVljutQErdyi
VP0O6BNRXoHYzx9eNI7xSQx3TTWYiniOucyOaGFZATdFtkLyK5fbyBKHJIurQXOMbn5LsIiu5eW0
Fe6s06mfjB5sgM1qIuI0p40/91uTaM4ZT/HiWFCH2knWRan8LUzNxEJLebDMpiyz+I/I23YQolYX
ne9Z6DfyLP2WVGZx6bs3AiBsKndZKYDqUilgMnbIJTmZan5nBY+wWpt3erOEHSQOuOufSUOwpTRV
4j3WVi5BOntTH9Z4b/tlHruJp4o2f3351m3epZSMUFc95N6xDw0DEIVhjMljweWk2BWMFDQkusir
afho7FbSml2TTfCkPuJjILspoyAjjglkXjZ6y4FR1yWakCzGvkWzG5gYLBcuTGFmwqqDYeU9h9kn
dW/tvvSgPbupsx1kAcAgsaItF1okdjXupWtRDxCOwN7hjttcpP89Nae+h84inhoqjpz1v5O3zdHc
0XfZRbJpSEd4QuPHG0jlbCqrqis6i0UUFMAx9KscxK98JNkky4afCSngP7DFqG04ggRskLxGDm+Z
mWQKRoM1JFm0V/aLgIj0vC9XduYcIqKaYKRJtAEiYBcpgAzObFaN9/MgSWkDmHCJ44UNOrXwZtPX
o52QYrPbeZ2rwAvbjqgUuxTrex+nF1U90btOEUo4I6Ol0DWnU3noS72481s9R/QuJ0aDKcPVk9lP
XTB0mxbtNEY0MX74fonTV6PaM45lMVfcojkJZ+8d4wgHr/QjjTyM9+vnBiunauRthVeFnrOdiI66
sh3kk1hYjf/c1eyZ87W4DgDz3zhxW8W7I+eoN1FDOfsbn+W1c4/p4zwH2+zz9JUiHBVoR7j0v8qX
uOkiXPr6rw4YjyW+Oy22G5Us/JWn9t1JcgoO+jNcR7oPFVyvJK+DssveE2ojq1bmUJ8VpTBSU9ji
BFnYeNERVlSb+yHlneaX18SalvvJ2q0ezt5Zenq658rdTSOu14LTA0XOCymKK5VJEZFVJXpH7kCc
WLfaG9JpdWSnVZmw33m9i9w58NeeWV1HtiMrMjiS4b2Swiz3ZbRWDQL3m6ZaUEw9AGbiF+LvzeDN
zggBWmBJEgiFQRpiA/hwp95ERViQ+22mugfdQEscQPIr4NSyUsUoiRuATYVrdmzcU/Z/C2s5+0VS
6xoEXZNBDCUH5ahZk9j1/DacrrMwGcLR9W+TGMQxa2794nKnr7SDvSXO7UOfIxykEnl1E9LN4VT7
s79hZNZGy8Py8do00Cwzg/q42XrSPTTZTSAdYWUDKkbLkDFMKi4wxygjk2grrGI3rO7LsLo0o0ix
LosQtoozTWiTeAXzAVXKwIgCZRU6OL6QyeDGLYeAP265J9Wk3DmmIhNsBJPpSw7qRYd0w+zBcZ71
MicNEprPRs6epFJHuSzZTHyHR4bVesAjgnEdl8UuSueFeKErVdhjK89SfIe7k8+1Yk6e3qwvf4pu
e0CDBtV2iXGfRr1P7CE6hwQtUVmoBI6puhrJ7mIwLrvFrIHOqe+zZx/mgqvDjiGVdywXHt6ns2gh
rHANtqE9LPiFlh7RsIPxKAmae7OHSu5+dAon4Y4UHzjJ/VciylylDh7dkveRc9s37kIRf2wY6cHc
xptG3xuCTXsBLqIiahA61zxNLfXl549DFGhHxH04snIgvWjmxFkgeZJ3bBR8KH3CvjnZTx7xjmXH
tNvn/WEpN2kwg1x9iQc/uqvrqUFfVjl1iZ8TtnSNRZnIKZX+dPJMeGvqgIW32dRDodl7lFa6wY4m
XHV6nxgkGkVYjNS/HxAq4WwA055gPwzERJK+5l16rwYkULKpeV7jYZSIFSelP6cksiO9C47e8LgK
nSJrIC+lfDZBIGDc8+YEkNE62O3kj4NmT3JSStaYGYADxRFW2Wjq5Yl7xod4xdaEc1g8VoGfdYgc
2DAsgSmn4BjRhSFn3TG/0HUWDROLqXB5vtA9w+4cNHsA+pm6VSGfjjpqbRGC8Y22dywI2pkiGPn0
o43m3CFVciOj+VgdL6s3LaZ22gHrmtZUDhxNeqwJXGoADUQHFUhm0Z2kTFsCfYGekuaZZFE+55l9
CH+XLmgt2+ihaguHYd9+/8h9lnJegjM6NZgUttg2vQcOG4BbTfSbxDnU1dow5d3N27gfvUE7nHFi
Gx3zqW52mTwpXn95upjIjq0VRkAm4ERb7PWtEhEoATY+pwntzxKI9GXv7mnOJ/rAUmCBRQ86jviM
DVWinM699+UqhK7Qin2jSGDRSZ/6BD2riNFNkzJwz+PRasQTk8NSu8hpIDbd58dZK+Wob6UwDvsO
6a0TsuRS8VD8tER50bMDj7ELpdIaNrHyLyJKnO5A998keB7ISVTPnarvdaCPrsI54rbxNNyKK9ln
4noiDrehYJYtvmwTU3imJIWxi8pMq2v1NKEZwxAiH9vSSzUx7QSNHli+h8TCxAQFlRKj+0Jq/dTv
Hs9z/dLzG9m8h5S7WmG9pKAPCUZnpj7RTJS99G+DoZoYHZ7mQX03sJnkNtZo+C1G9omTVa9jttzA
xn9R7qPnDq7JD1/Wkqv0Z0AQR7yIKh3b+y51DTPj0jBEZ9lNr/hFZr/NTCW/7n1/1KEQsegOQEek
R0y4rhi+5+8SvAtMonQkKiyh9slZkRTCEFiZ3drRNfi9swuac94UL/rFkJ62796IiycVs51kJZBF
A/4qaxdCMpR0N62b8A2AqGT6YDL1UjomWUy/t01xjkfDUjswRYHQQulA34DeR/K7e67PrYzHeKsF
9901KBZYFTiaMa3mOBTiWCK6Zfe4XeZkbf6vCJ/OnueeFWqwDdIUF4/LoOZlWiVGiL4ayNMpbIJn
y/8UvtpDSNtuWISR9UK6MFhmZGgymZ9ryIYDmrtSVNuITt2XgW1TeZZ3Y5Qk5WdLflU+ZKgt5sxz
NjxYzMm9YIyU6utBPO1T9ml6PUtHlnrJSyY2o7R6G/qZX6RSULbs/y/Ot4Mpru6o4LxqSejZOQ74
2AtpW/YydMAANrC9kxWZEOkCsOmbNj9g8xmrkG01B143sNuIXvV4Hh6Y3QiyY/+hrQLTRy2Pxv3h
P7l6EAo09I0MqvAhKloZOD90U4pW53fkkDYSWJC7QPhqb6v2mBByMRDnUJ5sZWSfCoRzeNSYwtKD
Qdjd8PGChC7V7MpwzYk5KOtar5QHste7D3XkHC1J0Sp7+EUSXzp1VQLhwjLyEghFL5Oz2e4S0X9H
KOydcZApWEckaOVKGTQ61AdFU+tUTzcEwpkvq6TtRB3sbmoZeoZW+QLmIRmOc0JtSxxHJc/w1MXJ
fVHX9QpkoxkpwO3yZsbVa2TuQrdDKfnVlpdA3jVi7SotIGa2uEVvN4mZvT9tbrMmbqApg9fcZRzT
y3nfKRK5xV9/pEIWmvUCuEear/qZfoT1m8g6/8UBYi6hbgCJSuRzmOhSKG+6xD59ZKaa0baH/UNZ
PyepJ1UIJxKKGjtzQEweJMfiLnPOhoAuORaoxKKnseLK8s3f19mWtQDaYINjH1ZmJrMwLiL5UN9M
pNm5qWaGHDBNjrecF1P/1H2PASDjRH31zR8cnuADHiZDA8iE5jEvUJ7Jh+iOR9bJBqyz2TpWIRuD
XYz+y6D/dQSvoJNJpiU7tlXsOHl+VUu7r3D5r0QBlHIm/JwSuUDJivjdn510f7vGAPwIdU1J5Z7k
4Lv35oARwuBi4+fgoBZ7a959r/kiIjD3sIqxLSaldwQBb8GevXKp19+z2xdQvjftN4PMxGQVB/cx
T6QYFJ241WMx7ICD8wev6DNYLsW64Dk1SnWy+t4Q1XDJXUSu0nCW7H5tlDxJ3lK3itei0XbUrTJJ
7eEtkTp7STzLE0T5vLINPoh56FdidmgT+xo7klguJ+rNsnIjzd5RFp5K7V8kLwOeW0k79VYN8PHq
64bknHkf3UqEUfWgtiEqzrDEqibleZCyhunTFaA0M0wcejkakKmrwxlM+G6CGQyX0sv/PP9uuLMg
YGQjw1t0iSJLnV4lt9n35KdEYlP3lnQLr9LrjeBoefpyWoGGZ6W41yUkZLjnITT18ADh2r1oQL0Q
fetW7IahGywU2Xv/3Rp1YLtNxD88cH+ABtMJ3MXtpIBgu+tGyt2V7mv4uycjBpfXiWvoa0LmhxEH
blDPZK0KUHFT+9Lmm0GDqCaMTjubfkzkV1P43oAL8qYggjvos/Sp90hRtkbZQVp8s1EIi4neLZ5K
A0Qlp58q8+gQEbBQnanl+NUphbvMbIvdGCWmvZbokOsiLGVyrmlE2EtXPYmL79nn3rndiaQuLQBz
CP3nzFP99Qyjqh2+WMAtTdLK7DnKsviB9bYD2Frgxbb/IgOYe8fGZWJohOYPqL6Z4hu/RInOODjz
feN8Uit6bps9UTdMUkLAfhCtCOa1/nL5I61WP375So38zFrYOUtwHeSNacLEutvoW7ZnDbEDnjdw
/eWYaS7DSxXPWBVZ5bSUTf1Pbb0nrNzfB07VMEEmSD+e8xPamynsTjXD94t0EzDH4ffYriFjBVaW
mY6zWhhnt81HlI5KR1XDu7jRi+teY7sUng0sGwM++yJhLw5Zx6b0Tp+g8nuze7ztxmW/hLl3A1mf
sCc+5s2gymbC9zbAPrwdrUciJeRo3scNK9S/6YIREhrPpGN99pfOM5bVzKAoJukN+rD8XZrVkN34
kNhwrgVxPUwzTn0qlyj+NDwVhC64yXw/VK2gt0fb9Jo3Fm+4VI1CdHJjVFjalBhdlprZ4uo9mijP
Tr+RdwVGDr8nkVqMCE+0Fsy9LldiSRN46vXAMFvkBKgLPCzkvpGclholke/B+8lQvbtwljI7go+m
orFTLJVsi8A9Xr40H8XBAEqcovHK8pPlg1R8kP0Oo4Ky6tFaFCAf2R68tsOHh4VZ/9LLcIchPxB6
s0dEESLAsVILMaVAYtRMQYTPkoJzUIb2VqLzpaP4PvVcHTNsta0clC5iBZxxe5vlsThi1+0SGZ9Z
FvhTeILV0B6aMxmChJtYtxnsHUfeQTQigR/fScvPfjaH0qPic9PfTyrPCN4msNcRXAKtxflkH13H
XFh4m0k6xMXOgeJBcImFC+D91XlGKuP4/BGIepukulz9LvHxUq8tceGRlz/6fJQnJgGtXkIXDOSf
LoYLNkhfVNvJd5SCa4VCSsg1BYhiA7gkWyV6dTz20Vh0ou0uSwZWBOyO5s9f4Wk5+QlapDvsGEiI
8cnv+6DokUB6iieK0+atY37lyUYHqe7WsOFIZCJILUVx7n1BLT7upw92MTKanjdslkkKQtkslzmt
U7CTyf0IkliGWsEkmMKUiNZxAjEcpnfL3r/i8GgTGSOWrwjaHKB59JYfTk9OG8qzfTlkctix2WF7
743KgzG2lanHsUjzkvwlGsNrZ5EsrsE6wzAE2RbdN7gw26PXEHAR0B6RK3cZ15hHUDWavw3zBaWT
Oexish6muSreoTnIEXGZcAsVyB/FWexjEqXrCYNEFG1ktq/AsCkpu86EU3CG9Hf8S3ZSSkfDLE/8
Q6MkFUdKHEJh2DfqBIVwFL57/X0SwpbK+RCRppLcwTVXAYWgjA5VoGNm2N9p6cmcuZyG6f1P47vA
vPoFCex7zr6AM6IesvH0wdfQw1qIXzyDNMQDYHdx8pCxZYdtR40AKQevyl+lvTiksXKpz+Vu9MnZ
SpaVGRFt5DNFX5rtpx6uTSTWyaikcsqkdgTxGBJ5OjCLIPKdLjm9cBHtqlQrmAPi2EBOkngkela4
Z5c8fVPCSvUa0phm46HLF++RC4CsSOlkPnRStDHlQDmyZW5YQlH4k2clOhx6L5/g/l72v+p47OPD
t51bzPy34PlckvnWmBFhExXErbsjbAtm6KgDQpNU0HOx1vi7ctzHmvuMvRKt/ZPXA32eOTVQKZur
8niSfPMRsD3Th1Y4qExCtYUjyVhvTPRvQSWGQ2jkR158Hs7+D4GgqduxW6ht/7liRDc1483JqaPF
Gt14L+kIZJJosLNV415QczuxnL/bBylIpS5Tp2FJSmYovjYqt1OD+e7B9gI/1g4RePhPgbrI5Sp2
I+rU1dmiPgpAsFmD0O03A/n0kcaoqWLiRuWQSfQyocFStBBX6gZWTrQaQLzWeKiuSO8WH9UaryoU
a/ZLqkuhCnykJBn+ERyJTl7CFBMUbXAaA02VRjbQVM+FLyfoJvACoZzD6QhX0JVbhiwg0l4EbHjx
eJ6i2HKUr8Wjtm5tbSG0GXwhc87QkrguPNGeyNW73Lrnz2K8g0WVdNyHgtkeMV/iQCaOyPzfRWtW
mOe2f7ovXUQ1xvnbjPFqLXyKEYPSUPbJzl+77sIpBB/ttmwt4qfr5flprpPwlUvTgxecPk1+4SwS
CaS9NkaZ/gW8ZWE72apfyLlVSewIFsRi/N1Yvpvbfn6pbur0ome1LecBCyzLavXuqojEgqBXa1+r
ff+0yDyqVdNK7hG9txVYsFapuvpV2HPiuofd04frytuAD7HTwYLz9Q6L9VB4Rq6fwHDqJOSd3ud3
CZxgd0wZuj0zDGDrHJoTfuf10SilGjwr0TWlLP9O3JrA/jfp67QXDifKDKOdRzq5eqtr0VSaK5z6
/JfWvLsAVo5iKqCOvU+IibrRc9aZ1NC7TcAqMhNM4Ln+Q5ovbpLInWLu1ai6doBtZLNxjZkXDxRw
WKpt6q+Vy10mYvXFicDPrLuutdpW8yCq9YqL4+wC++QmvIxIMAM6C//9Zql+5THT2jIFqqDCFqO9
KwMxTp7OntbBAZvCSkveWLz+19pGlbuSpRh8rNEjP5toV4kL/bdrRS3YL8I0fN5gygK1OSCQLnv3
jcmj2+Kp9IbAHgSruRE0v2xvM8Zw3Kx1iq0yrrmp7fFKulhKW03pWm196azkCx1r6uaXmlqw/maL
k/IDk5VES4UQVtHU+l/7OpZMCNdzezlbZo224lQLHK5kNf1u8yFz42vFYgqeb0whlSCxVWDMPBog
c7PdfMBnHbjOnrJHyiQeNP6pdGm3aIr0s9pKpag00XU2KveG3MyFiSivZt+L6aIJ1YruFJPuYHRJ
C2idI6ohFjdUQICuRkJNLOjrSlLvbbq9ST8BNP4tQ0JzwTy26Kt0nDqisRGz0CxOzksXX40LZEjn
CMJmArNaWLFR3WECs1rk5ZjH7zPXBj3EEKHyj1cWLe0vouGuBxk92wYV0bpeJWc+pRM2s3qAR4ec
aV/SWATfnO2jt4PhMPS5+FrhYEbPx8XpVIaDqAcoY6jRgl1J5Jzl2A7FGid8SYTSvbBJ4lfTnO4+
H9J4cm9BhCTJVmcWSJ5yQ8O1+4YL0zVGkYfVsP/pWcHnChMnir4Irl5UXim3frHireL/qMx/Ho2p
C1bx1w3GovVxOe2EOoa2pJd6FP9Ui3z9JwoQA+e1f9OCdkB8zGCqu9h6bZrqPpDEW9eOJ2pDLmkU
a8XWP+SIs3NmR3uz71cVS4fptQoZgwa6fbE8OAQRiE/+stCGy1yB9RnXJmp012y/DZk7eVW4Z5Yy
2RFmxZqTTeeb8t9/1G4D6q73UoYTcPOkJrq5HUdHnraa82BCFYHX7tmMxI5Yv8mcpU02G+PeZBPv
LYdrIpjZuGob2tI8MPXR77/tIHgBP3V2tXtJ7Om1FgVIYJvZIEanlW5snH5izCwO+T003V/Z8EfT
jRuQQ/1SWJXB82EZjphJP1/xkxRiXtVlATY4y0j+dot/7F1SFqup9JgRpJcdLNM+9MCHt/oNwGLl
xqj81u9sNmGXeehpj9tOlWGQMY8LutukUSFRB3jSr+b+RixrV7HbNPnAiP7FMcRCfQdMbOGdK2EA
lDyXsWALk72FItNdJQJZIcGw2wN8vSr3qd90bk7oxBGty57HB/bn+dTGtvJROxOyJxwmx+RPLvpS
fHS7fzYA406AxkZDTJqQcKv2idLkHyr7S/SrnYMpI324XuQVXDy9n88OiCIWpC3B/VzCvr4oT8Vc
nUfPlJC3GMO1x0GyfozkoG+7Hyt1X8FdDVgYF2YA7gtSPFgPCuJ6cZxpJuN5i8h4hLiYlQOCJvHk
Mwye1OosUC4avasoyYO1pfiylScIsAQP5wPKL/UoPVIdH6E8ad/kySy16ESz7DzzuvZxOVWuHKYd
fplEFKdxQ7tsPmcpbF40km7g6/bxkcq5iWRkZSirgdalhLct5KhckMgvU0WhRZXVcLhZPSyQ2gak
y/wNOxQPreP347lqKj01IRJhUVdXjIWc2fvuBqieXJhi2skyOCogLBLHD3OqK/gOWcL6uITkcd2o
j+Xrq0CvOii+6gbPsUY+Era1bzj+UlwA1M21X3IBbSQHoAPXDGIRMN6IPyn+RgrdqyacTLQAAjvF
ihI7tHNx31yPOV1IR6Hr98dlZiHLu7tV9be6h/6608FTcuX9HyVD3A82tVtBVWv2LQpBZrcspv18
7bU3B8LRe32OE1wgbvlsxk2Qi4uu1oW28/dukV9Z4rM3R8TOsY6AGWNLTYO4/X3ymIyn2/RJ7qpD
sQv/xtQjtQdFTkTI8Y09zZdiMQbUOajng6onI/Yy9f/1OXuUHSwnd72Wi3o00rxFwbi+xa8+0mjQ
Rg5dAL4Lpp5EQWYvUv7S7MmUtNmeRAfGxB+/1Lt+V6rLs254qpGWlVuBFrSMwIlSxOb9q6I3S4B2
lHuRrjZU1i30MhnbvWHsV/1173z43ipo/A64rbpykqYc52K5PBkpV43pc2v2MPfe3oIC6bpkK+Wd
2x4WlVO876gnbbz9RmjncaQ6/UGySs4jVehlVB2ZVRgn77TkfA1FVNSwu2gzC1x4PczvZvDAhaKu
0ek8awDqD1EQnnGHu+b99AupsDbYkGk5qhNwYYj7TXzZ4BAawPg/GNHFvr3QPQwTnHmuql3UzdnE
Ejwc1wi+n3H2xbTy11uTzU5m5bo7vdocXezaq3oFX7G8LSjXMP31ZqUsQnJzzqlBTvDZjk+X0C/L
ApMoQ2rTWIE/pbzwBOu+HOIUWajPEcTiABJHj99B8OlS5p4UUcs9wj3ObTQXe5nCR8n62w0Cjm2B
BErNyV9tIA3nsTVECCnd0wwLRV0gD58soqB9xReQQXFpg5b4CTv2a2jfkCzp9bbiLdeLeGLy4oUg
melR7W2PRYrgG7kC2WBQDfBmkYjnKpR90lTyU5bzI1feyYSAOwxA46/FkXKOul82q1sZIRZQXLFX
Ge3agfghR3K5apRzCER/F7SYymiKQwa4XlAFZg5QiuOk2Ptx0uY4u9hnHKJzsClRMXgJnr2QIy1G
OvF/aLmpcf21k3xdjTcGyZdUEhoDxiLqUo6QJ3daq/UiLb8l83wVAgIDvMTMz1zPFzLVcVGpALEp
iy4nuPvIBvAei5fnEfHQNhiqopyoAnSG+lAcUMCY42gkIJoMLxsECqClVQ50kCAw2IfhH9bJYmDC
OXx0rL98p3WS5xAQYh+ygbLG+smkTDXYDZoE3mMw58JEwj1BpqIhrR88TBX2ClGWW+88P+oE8g/G
c/+kZvTuVye+jCJRmqICpnVBbbyFcrmGGkJVj/vkcqMcSPyQzV/fRHbp8AR9GHesRUUJjiDjwXKd
JmoD5C8fgWyeOwjxIdu9MEnxwkVPvQ/ZNwex8obu+5s/Q3WfhCkBBv/Y+PUzmV/FVVOkYkx1+r7v
Plvro1M2yFlx7KXPTyn26+/SC+2aOU8wV1ovapG3++E1Kk0ZkqacRK7bI68ioVnZ+IXy+iBcTXRg
jVNpcIoiDgAr0tJk1Xesqqsfk5AYq4MXqkIIkHqw1hq58ZFscrHANMt5p1K0PpuAbFjjO7nxzgHn
txS/JlGDf7AyexkocYDmO4H/a6G45nuYDn1a0Iv8oiHyWJ/nPCOWYtcMIkoAbw9iPRYufYRLBJOk
QbEwoJRJzXKMInH2TnABtLJQV5YRIYHb7RR93EHzPyxCLmc0vJ+XBbdU+DNgVo+E+IpUw3LhtbTX
q5nGsNT9v+Llv8CXyoH7fY3mSGsGhW9vciA/8ZYSg4c2I9U8Q6sXrJhi3tptgchNKDlB4n91dv3m
6VpbClzhxVONXD5fN4+yb3fY9eFKBvBDTtD3ADwJQkPglLmdTefOyuP+IkBi7kJBhAqwRR5NhVCT
i5hJ/Butt2/g2fyh7EB0Gew4hmStyjtPq9ZipyA58MuptRpgFfgoVskDcf7ywH1wFnr4aM4p7CHY
LpX/LTXiWF6vIzrkaFarDWp8A6a+lg/2pvrfkEgWWBp4YmdYfalD9GUbh4P8wCMn6yXh4SFibcho
mx5d+4HNqDHwuIvxs5nWE7klbuCWDEgZc+YZPzehu3OVdmaECdtvQ0W4E0zz/1HQ3NEJniFbQP+E
l+X++YMhTPMKpbg7q0REDCGj2paecL9FUQDxwPkTxqLoX0Tl125A+96fbdntZFhbTaXIfrF/eUek
m4PiJ3gkrMjdQ+mW2gF85wWJTloFQFwqGGJeYB8ff//U8iNaEg2x/L0xN2v39nSU4Q1F0meDpW2/
bU/3noqmtgk/mXaLP5QCJ34xaxQ9qD8A3g0hcDoKL84Zu/cgOLqGlW0KOZl7KzuZH9LwrZlUhrGx
OQDgODVzLPLe8gsxuLLACbMQQvpVXb00yQ8URXYT8O2U8N+rVLpturnSmNRRTMEsnXRmRTR1YJhu
Ik3GCYOhua/B65MrrTcMoqmIzhOpXFg8BrKavKXdcGjMjTFO1qavNX6ZSh8mWmzJAra0na97eOtz
38SvBaovE+p5GAZMNAu90ImVrLYAqVvJdIm+ozxNN6SBfZudXIMy1uEm2OyHrJKNuhOAgk2citWY
NZioziJ5fUvVMDpSF0ZhflhkEXcseImcn3IzYigD+dIhLCwZpQKEuW5azLB8IsfhH6Y3hJdJoq8k
p0tZVGxSb9pslsDBTH56/O/f7XofZOsVDPrEjlcAduy3yXcEGwSDJ6cAx8hBde+0C13xZGYWge/F
oc5O53w3yov9gs4zqSnC/vc2ejydXpi6yDf6htu1sawG5fQ1UxmUt0/CNfHpaqLwaxmK5sMMPkCd
4cMEkyA4TSKsunwtbK1KQIhVpQSJZi18UdOpfHc9UkUDUIP2k8h722dBMAV4YeHj42wTllGzLbp+
5w9Bhtv8/OYnOxjVmQRbJ1jDSGnvO/O9CDzLzB3bFyNOYgYRZ9z2OuNJuRVM3GVyIqSLyRFKMU0o
32Lt9Dd0m03duFHjTzTwdQfd63AWNtD96ZHrzw+Uj8hRJgn4KHrYpT0B9XzpakDJRoKFaEfKHe6S
iCsVAi18WlTSdyS+a9SO9y6P4mKJJ9JDckL3N2VWKnBIang6vCG3Df0kcp3rolTH7a4jdXfLZt1C
1MG29+PCCCFZwBBfsdDqa/gXFZkZzv29qo/ol2MCp2O4C96+CO6VvLJdhXYWWM5HRAlT00E9dyI8
VDsZ6GIKf3pp53EIHuXYvuXqz7WC/IhX1VSUwe8v39F+SZvBsRgK39aILojOtl/TAOxil8RMZGd7
Padf9O+fa7r0hQQPuJ9JQfKz/fMPHrb+W2ONElLqUkCdqmx8QUlVjgWQrupuADIlVICSJoelHppi
gsZeKKV4nOpTeKoMrpXxbKa8sEt7Ptzt7GyPGq8wDOkxzFHADYjSSm3OnXIoTYVWPO1XJof5IPSf
ExqOsiMiTILzbGGuhIHtyhzMtyYtn9vg3iHmEpR/lUZLlS38afkS97MQFG3DyshxWBPE/EPH1qY5
PuRaDrOxvbmui4/kL2vTxgy+d7coL3QcY15kty9Mtwjqmbxrp0/77PXz+IvN/E624q3ACbZ2BcHE
tftfzlPim/pnEsdI2ooTQe7usZOyDwsmZEmMQZlzJRq5joYk4NqeZ4aKa4exouBJMx/6kwpDZq81
VncVfc1J+TIJDF0mxXZhuxkrMSBfZBEHr/4671Smn02aY3tw4KxVOcub5k/RBNToGmnJ7Fwd2YSh
/A+FEi3NYs941jenO/p/bDbLdML4qHxR877sfI709qrCaSbB6ursw2yudD2jnKKYf+AUfkD+xp+L
DhCEArSLxNuZRpFBLcsAreDN+vOklJTcZ36JY8nXwvVHSgPU5+gGcHizUR8i+dlX3PTnEJqjf9O5
eg2eOw2fGHTwppMx4EsHlcDquOxflzhoCTUosoMtL5kHOMr6+pBbR98T19a+TY7JwZkP4RmRMLRX
SYZLAZ4H0GPvulMzt9yJTMiJS7SWgwBl5K9CkMpGgNd+GZXwouW8MNVN5pMj0P172U0ipBp3TEQ8
l0N5DhmRIm1pkSX/u1GuDZLIIAdtfEQrXSBzYjr0spBxvMj/Dww/F5AMUNY7Fg7ezXtmU95TqbM4
eq0nvuTBQkLGRyqG09g3Cr1WGdRvboE5cWU0jxGvAVRdBpJV+JAajOW4FMiYQURa1iMMiU4iJeu0
B1zKaOy6y5QjMYnszqDuVukV9+rn1QmnvczPbpdUPLyKgX8YiuFGuEG7pUi2GzliOJkOeO3Fnm0A
1yWtrBCJGAgx0Qz9F1d0ZpE/dnNhSQtclwChEyKsRcXPlWQRUROBpxWeKCiDY83k8L6Zi4hc38U9
sl5W0jojchQcq4Uqi3UuIJElwciDVfc+6+w7xIkeiGTTTroX7D7hcPjDA1cBq7bTmDbx9zTMzDEu
TjJInh9tATK1yLRloIbVWNBly4D7R51pfAtYPTQ1nao7C99MkL1VnMQubnqW7UE5tVmAdd5BqaDY
9u4zV3ZqclBpoQjqM1yQAb0k5c+XRybEbTIF5AAiJr9HZ3A9uO+mv7hUwDAzVKHrJ0JF4SvxCuhW
TcXS3vU7Fk+7/hM8yje3tuS11pPkRnZcY3ltzNQX1NWQPDLqBNR94YDDB2pLv2a5vo/pnp9OnHP6
thLoHBCPzjgjnL5YqAv4De9iJl+kKjHng6Yl3nPvLCwW8717SSGIfIOlMlrSsKVYKgnExFMdTkDC
OjCzOfNvt9O/IwUGAjvlOxZIQXxWp5mlasKIEYST5ml4hB6UgA4YMBf96elBzEDkPxir6dE8gi7N
arOYRGrhC8SRAQgSaRw7DuXxZ/tZUsKQF0xFeXtD24MvfEhbSz2Euwsob2udit590SArQgvA+ZnP
D18HSNVer7pDHjGtOw0coSO7lIgbePgTA4QtA3+XmO6DQvyiWrioG0anlxFZNT+uyMTkuwDd7LHD
nG68kzahHPzo3ui2+T8vRSMFzO+j0wkmsCgGv5dFYCtkU36IyUQ0KyisvMaCEREj82TWmkkekZpW
SSGMlp6DOVe6S9VLBt7drdJiFVwI5EF0aqdV6rHrU9jzYNfYgPj2XoTvcwwyMBI1zJz0EsVKlXmo
q8ncqutUrKv90duxV5qWaQOIclKxofCms8nNjSZkdxVutKCWk0HOPlxAcIf45ss9qBhuUzZGH7uL
e1vvg7YdADHCJmsiEPLLEcifynfUBSYQ7oLIeeGGPGLfsuct5Zh1sbBOZZrk9AzgHlejHm67E0AM
CEOgWavHyTYlx7OLMGIdJr8jc2mZUW5YyLvUEoVjatZ+q2p2Zmw+h0vZhjXarxndXlAXIO1T7Te+
SPi1+cHHxVIcEcV0GJftkMvG4wCLaanAFRdnneCQI/r2vu1kaT4HlSwO6hkHosKGDm53IOSIYOJi
rxOqRBf9KocuP9yqKa2x1ONUGMHspKYAQ9X0p4W5lfYOo4SGxM1Fi3xeLplYAI19ACXbG2utTW36
hgd5/zzJBZ0M0iOaL/b0MaH4mUWCFBpLGkdbOtMRZah5oNgcdOU8dBlmjH2zOJ1EFTPE5ReHC6V4
ElDKfZ+zEG2EKiTZAzM0XZutRtSbU4J3Yav8qm5ABPiKRaBAHF7IDb87cfAUNJKvNI3f/8ai9FV2
Ob4WjZVfY13Wf79cwZ7ujXmLn4zXH2wGyijeLfjMTRvdUtSH3vvGAq/p3AWoyudtEcblZzn1lNQ3
gSXjfXF3ic/EZl6pGR/lXaKB6/hgFd9uH7ZqGfWY6nB1sNq14JSho8noqjnZRkhirjg3dhAki9aO
KoLnxCw5r+Jy4Wt9PUcU/uY2+4+gyTNYiTg+B0MFb4/pbtKsBtOd6Cf8BMtSxysZJy7rcJEiqt66
dtCBTUBAhooVpFqZ8xrsDGIPD5x5m9f907rthhZfKcaL1Fh8FcZcOm5oKQmhYeqKDDhTNrlMPqcB
2ZpBLu85vbxWohQl9pj0i2lO40PDapgmjR0MG5JSnxyLFaPqDYhBFX3AUxHJ6U0WKz1xYXemifwQ
WErV+jlCtXIBnMo1KbVcE/KoujP9TCd8W9CwF+AbQhVclDSqAXhWiB9HVB288bqVoNlmHVbLcHFP
4v/B8dH5k8+PsN0qakAARs3GPd0YqtjORIhpOl9HktYNUN52Y+KB6PF7Bm4cOQVI9TpCgTA1jnmn
059qN4p8orZU259A4EFijkUP5VY9VYf12CyuUegnSgoH3y8ZaORP8lN+48UhbB/MqKg9TNpUWNwZ
zyVtNNecrhYqLJ3sH3wX5H3I9VvksVgxnMKjKeAJbsxxpIk4YTl73I8lNI82YCC1PIN0ByK+d8Ff
Lrl7g1teP3701H46GpaARtrYYWSO5iRT+n5Q1y75uTCCNBuigC9Q0sbnrwbfViPPOrjFp0aT4BYc
JVoj3T3ET+fd840C6d66s1e1cqGb6ml8oyGdxhYaSrswx86CxBta5Wq7+qopVgTA9xx20BAhSYq2
ZSK6+JVW6Sk8HosqKD0UEF9duIcTedEPG5Ey9b3rhngTuex7B8MBM8JYL3DjJ5yxMnpEWGk8vjyl
Yn5Jgt8uyMPQIbTfsapHi/2lK8nq4Cis/shvezBXUvQOU89MUBw1ZC9rcXaC1+wJt5hkBqRUggFb
lgTqVoqF85i5rN1/rcakB+df1lyv92W5WdlIetYxRF9YAyqlpqoL7uXetKQhXHAy7M0c+gvBDMaC
I1W3RpHcZKrrQf5VC8uHVOU4E4MrpAcu/+rz/yzcJQRn6BJrH9VzIVxuLT/J1ApJNMi52swXjpFy
5aCXa9RO9o4kbhYFJOdteKrOZAb1lNiWXRd4nlr7cq5Lh4r2TsCrghRrzZW2i96nEuzywo2fr1FF
1rDj1IPMuOuZI/KXbIEP+p/s4ujmA0qj2s7fLEzcwyjMp/pjIKSp8pBthzN41Oa/zdU5Zv1Mxozh
nlXabqpGlDlcKKVbmgfb2lndGJOyACiqkXyuGFKqCObV5BOr5BBA12DTGg+N3iGiKVWLJOEK559j
TciHuY7j4pM6Z9T/RW7gmiwq8syCdsqACcOLNo4RkOYjSkrFDhtEcqlF6pHu+DpU3xl0FgjuImBs
e87gN3A4u1P2KXS594HkML58eCPQsx8vJaf+8grHEHOwQXXK1iHsU7eE9sl2k+dl0mkGDss5s23t
2p2N6YtVllnu4gqwvc4ZGlADiZniwPAsueH9zz/cj3l6EYg0fBI/aOdMdFvFLewml2vI6Rr3cbFD
f8/e9JGMC4ys285/p25yWmeLtN2lqUQs0aTb29c6u+2hb+gpmxv5TOyHkqs4xcDnzPHZrzfAuc+c
qg8/n0ekxU2uzXALp2EUkHUtQzi6YKLLn2Cb39HTI+BIH6aATyvSvBcJlqnV8wpLtsnMTudoC9mv
CDxZqFFNRX9DpEvtzL0Wj7/ZnJk7mgFvNL1A4ora2KZydBEWgt+rm21bhh7OwEV2Nfd/aInYnmBg
2ZmhvE21oxVKeWyTGEBMHHKaQXiPeJ8GjsUlu4eJWsKgiqlXffsmSWtsVCfdwkD5zUtXiHnXoOY/
vFVrv8/EAkVGz13NNtGKPy47VQAjSVLNYToAIqjMwvSGMXh/YaeWHZ8SpdrFrizHdyXsq6JPZv2e
BcVeuHEH3NPlC6SNYEeWz+ROGroCZRJFBAcYdbPfGwH8ZnN7KKdWPuAeJhCqltlQxZZ53ZmhN0Fx
u0yPFkKBOzaQuURpZ5RXuMwlenOR9ko+PaYl9+b6hHd6o+LgSETB+gRfi5DTVjHc9qnZDs3EQ5Yf
S66nwUXK8kDcvkLsTXoG2hjBevEI8iM+Dk4KYKi60TP5U2Sq1Tv8eKAA9MUEwjFoPZb8mcXlnGev
PO4evneMlPKB9jDTrmE7ARo7KBOhGpUonSTMeG8QIkRRNgNEAY9lkHxRVfOJTAJ7aDvt6W9m3/SE
hdURQyBG5wjBmpR37mnS1Zsr6g+c9TXFltA/3LRSFIxfk7C9n70dpZH97TRJw83OR80PeEdiuRvH
8FwC1SLZ0iD7kjQKS+oKhVsws/FMatjU9BE5qvw0wE2LmdXDyKmJAEWltuAO1RdWq/fxn+FDPZcz
ZQUSkYLqGPZX/wHc94NQ4kZg+BanBd10F1I65avs6wRdllQKjp7o/DUPmTFxlS58VZV3+NMbgKCN
4gL6IRjv3om8XtXGNuuThhauCAtNj2VSFtwoOd8tyGGB35XYLol7/tRceIo6zcJW4C0QSGfXTUCl
4/TekF+fvH/4776YI37BnbAO3ckMNMsPc6JaEF25QhdvTtH1zsj2akSq4xnf4oYmfyorOnzYPRYy
Ct1+yc3cer7YSO28VmcWR/o/kQofFihH5pKA4633X7N8Yvb5gc3rcAhCcTLFvkiRDcxs805cVpd9
qj0q1Fux2l4UImWC5k8QAfSO6LTVFOhbS9fenA7I4R02LV/oUp2LJVngKeEd/wih9NVz3dl3aREv
EfaWdI5jCbWvS4R8qZcltbBRg1Oz980L2Wq1SuARjv+jWtM1Famb2UDbqw4xZA6XjG8asZ1yc+b6
tkEfKyCGUvzfFUWqJ3x6v+4OE+y8hLCcN2h6pxpBUUxwq8WkdLuAxoKj8hnQGVBUWuyXgwvUkS96
bMPlh+dOxgHs5nUQjDCryNNOwUYal2+5vhX+DAMKtz3CPFuIaI2IcSrRNKVIkB2aIlw4TndHmaOH
cyMwWvNHwpn8Ct7YKjiJHSdPP9aeOYLWrZMxTH5m/MlucyDxdrbEBiApp+HKozHJnmXVqe7qVUmx
tAQKI5iJsri2+LFYOh48mImcVydIyATHPSA0WlGsSZhQe0E70Oq7AD7PO1IUqq/73t1K8Wz/Sfxb
vBIrWxNMQhJV8ued/ExurY+PBNbvac1zEs3u4PCms7xByBIa4kjW7NLW23xiSOdzClXCzJcjLukp
BVsfJvlDUMMafA6YMtG0VBwCVCl81nCavFCG6kfCH+MjDzB+imio72SeWWNXmAQlIFt/uPQbzcpD
/uZVBEiuxO+FXQH8scdnjm9DuWndzgeOaDOtqRgLT0Mu0C9iuyK7MZGDd+mvcwskGqr+TWWy85MZ
0v+VNJjiCfD0NR7OmJ63dA+VDk2c9AJ57L8zKy20F9jNWAKXxKx0yRcB3hQh1y0zdqgSw0gmDH6M
PjdFLTiDQ+TY/dIozeGnG6Dc/jDoVL4coCvTa8nnIxSh/fRvL3cNbRYFtFQ1OOvTisLnsZiZG4OU
p2er1RRW++dGl/3GG5uYdeJHU+Lt0AS7qLEoT2UtgZcCOzYBCqJwjM6I9Nhf+MINRBe2pLTJ4CGX
7t5zvuRi4ETeBqDpVlZIOxth6w4/UKN6SJlKWF82Anld0gjWzGBcNbeSbtYw2PtRPTD0GOcL/kYD
uKkPwHkcfIeF4koiyFYl4uqsnNt3zDzGbqyjzQOjCd8XE3jx6UjTKBdmLZVuztKt7ScuckL1ur1A
/dQ0wKqzSY004HklB9OgTA7oL8v3Sl3Y8jlw5GgoQNm6Zp95UIEyWAPd9O1fwnCb285ULK5HmW3c
D2zyZxsfy1nWDpBFekHyteHGJc+uX7WlqgSOxZW9f8LdRF3CKM+m8XJ0NS41ZXyjrFWLaJUS2yqR
nXRpAqusMml0Cn11WhJAQd8aOD4hdCMoChhnWfoHe87CMkldnArvHSG7zYwXJg6yGC0EA3+UJBvY
FLaY/KMXq3X4ykeasLL2z/E5/r3F3i8bl/SZLajewAfGchlw5tbAV9XOtXjJuEbV1I1oltWruAA2
DwL72tWOIQczjes5/W1rVcJtCy8BexdKr3kpept2WAu9hatmjtMdnylyMcVPPhLpsYAXAfY5Q5nf
stelrGcuBbF+MshZJD2HpHAzeh6q+fbD2/SoSK1IcN18zp8OEmyZeBFWR5xrp+cOm/1eHlpVTU8Q
ryVVGVlMsoAKOfWVigknKd5sOMh9P54r85B6ia8sbNQyJki430K7YphzQ9bei322sOlNyCo+vJRJ
q8ZRY+DJpKPp1arAI3ApfWnBEf/hnMVsQC0cFvQEbRa16R07vMJ0sr7DZ1VWgi+zkArJjpZoqQk5
WymX2+0XdxQNGHRGCHGhveNMzaUhEHZc8ZqyS0F5AnqZH63cCfyBjaFLC+gopoy7r2P3Ackg5JXv
zaQVxBZt1tR+3T4E3GhpKDp+AncofugAVlUbm5QbIyoJOeMHYazOa+SzqG+oyNdrgNW6Y+67B+GW
yV2cs8ptVqgxu+9W1DtpHO1uMYzoscji9pA36fOID7EdWP35Yx8bSo1GHrbl4GfOWjkp/HJkQKsw
bRPwP6cobukwJ+Y6ysYLwo3TJgBYlUwjFF0RC6+/kA9pGSuy7hwQM+FrLzNqmKQ66exi5z8y10D8
KMR3mDE1sOFVmpbZEa65O3B5r/NH8N54tWxXZ7Le59BF9jzq6PYLr7V+7wA1prH84TFtaKbAf8NK
ISiGnPwyp8MJN/ajvrh5ek+ESi8ZUXhgcxSxu6bwrxtFFLhqXi4tLeLUpB7Oz0Hi2AJBh9k3KK0h
Unb3z18rEHVR/S2jR8bsA33lGjsTm8XtZCcdcgCFcXdff5t6k3lebZGEmXg2VW8XmoT9TEUWmNTO
sjnBbgfyOZvkaUozP3bfhifkel4fiNtAIsW0jDzwUtg0kVu6ghIXA61MMxAP9kXWmAgM3+U0rJL6
MwvhuPj2x2cHiXNCbwYJMQONrwrca+7gQJEtTh9T6EGOwsxDqHM4AUzj4/ugOJ3VmO6jLAEIEqxu
c6EZ1OZ1ukxB87VyHlO61DV3W4KGfz3dx+pgaE8OpwUJdLCv2EWpGwwpErK2rOkJPQPyN95OT8sV
0w7e+uXxnCpUUwtAZCExh+lQNhGK4UZ0FntHH4E6JUj1clO7EYg4o0rbCSW9gzZBdibwZN8T1m25
EYBGCHM6LFMO5n77A8WBzns6C0SuZRIwaWqYEp34vD6AI9h/8MBbu8u7zsma1LNgvsxEWDOwZ3NZ
Sj8yO5J2YADnT/yxJQFpe3yRHMvB4vAs03anQZucMlhD3XbfIsGiP9JsC3gTdIFoOEDxj0uTfUTu
mFt5eIXIICWzkSYmqTvcz5nXUKpBEITWt0Zd4lg3m8j/6X8P8xvbSFEVpKtoRJzFngZyXZXCk4QS
KrlpzJlA2Lq2zrwY9My4LZd1xW8DLeeMK+HoPc2fj3gpXerkd4NLab8zUgGdxEWSS4oqAAa33+uZ
k1wH5xxj4dT/GM/LbO7SuAvvvAs4n4hoYs8NXPU339w2DXmKifkBt0CRYKmmc0bOY8EycVmjJx3M
ZEmcAnIZ5pMqmCBNpe2b9/9Tk7dwRBzX6U45UR5N3iuf1YSgCc8QqBVk8u293aiPtql1JfAAxWdf
BP+Elj0M9otEHEn3BoGApAT+alvVDnqrwQBFc4JlEiEAZehZEUlZXqt5aWDfjxQ4lszvjo32HuYT
+lzJUPeDkQc+1WUvWe6keWGuz2fCcJV8tRwzY84VMDHC0inBzp2Aq1regMSJ0ardNJBTOV1LDkGi
AgiFWyHaNp+qLyrVOimNAQiitGD3UqCm0VvxzAYQtHr9yP1KrCSU4LohDR6rJdk67RvolYCnffOE
fxdmjAq9PHyiQvbgVYm5dFBJSet0Oga2tK/tnVdtbIVJQ/Gv8duiAbUdVVSSH3Fk+z493JvJJUKR
1CQbM8smv36l2gZlrhRC/t1R4MHYc3Q8tQkJl/bhyYxiiGuxfaSKw2zt1f1yTBEHEd7Mc9fqgozv
xFigDJYiNFrlhgeRD0bI/9cshVdXWAPfVyJDs6G2OBCNgtZzZiXiLZRG4QB+fnSE3vJ74hCluzKr
UPOASJbnQ9NQQK9AoDKmw2vPtNvx+vYr6CuWuqr/I9M8zcx2fexPMtN7S/Dv2jcsikjbUokSA3bn
0sz2zGEkctjJi2WlEkS+olWOHejdYpOTqwVXZhvvlxcVgueJVlnGALo6fCN1qAfAWl8ysIKLUtcb
vi7yRsfSa61sa38zf+tthpCYtMr+2ibO5ZUQ1bN/5hkTEOIMPxHWtkE1+f4GN0Md6aJ0+ZEg2Yva
oOlaXYxlohS0W4/YbeFiQIlf8bc9fRizOgbyXicCeCiSfY5TY/55us3QpzQf5wOKsU2btSMRrT9Y
sPwn5Scr+d8vCrl7ng/2r4cLZRTa/DoMEjETVclKXnN8/q2yXSW0frAFC+0AhiW8MthIyznjRd1s
pBjYmxjO3VYrCfjyFZwsgHjrYjzNeWkwcPCZ8Y9uup20+4WDhBMmCwdyVZV3IHlG8t2oN2xsVw4y
W4FGvZ5GNfY0vgLBXrVTlsvCpNwaLVLdMFmuJhp9fDI0ssErF8oGL7GUrST8RsH8PdovN4xab2wI
a7oA26TalV/PlLUGSA8Dzbgmxp/DwJkmmBqGB8xELh7nIsLAnclEJlesrHe4UAJXk6GGzG0kFTGA
A3ScIERHUdxdP5YsUYlyPwd6yiVCTfvTO7L5Oy6eo7TS+qWm0PA+a8l8U2+2z1MkbjisBjx85AhI
gXhUM056wTEwFzIdAM4Dz/ck/N2fGEUlehl289di3xdR/DXas6m8VRk7BxUxYaGJ549EslSmTOYF
CXBQlUJGvfKS8kWsjNmojZW+uvUpIxPjZBAEg44TNM3GrKGDYAq66A5UA6RZFjb3+Y+1h9nORPPN
Q6Sg9MgmkC5rECyoCEiENo7zY/KL4VlvQp/pHuIa3Sq2U5fMA0JhUguVZW5qk0KsKnM+6I6VEOpC
k9av76ApJ9SvUGc6j5cU//ug8cGHehQpvnKGEFBw0bGbqN3nvwe/CLbOtIzEZ09fLy0CkxgFt9f4
KuAxlLdBbZkS2vGR2Jp9U/vYwPvcy7EN0lascAQuZM/44GLfEBMs6GTpQ0JH4iWIG0et1B9TAtq3
YNRV9xdchTZvCcBmtW8emcKbF3IDto6aUnnCRYwmit/qU9oMXDVpNDuY2tAEHOZo8Eny7w4F6nqi
itMP1GgFYGV/z3phDBqCOf062QESe9sieuAlLNaeH83JPhLwGx7Ca0VZGswlrmljaVqrPtyrcj5I
RXV1lJnyGdHHTyJroG6Brbp1UAjgT2Oz+9nZmao8cAHO9Q8z2yKiLJ8p51v5rI69W0ZEl/3E7jLO
k6UDtjxZvqlGa050JkBEetgLE5agQne6T4OOmeb8wE+fWnymjB9shGBAMAjATugFU+AfxqEpmeJ0
ndnbYAF9OjncqhIhxLkhkW6TzQ4KG5bPrs3ZBYk9OzI3VitGKKOkAlFpdlyOtIhVenuGMdLJ+E8N
dCDxvG4Q7YEaJb4gqRDyiKslxghN6hum1Ox9CsW7CR60I9fvbyuEAFB9Y6+L50RqNWYDJv4psNjk
ccdzV484gZK+RojFkxfhf4MHkRyKjHWEBsNWnNuvKmEd/EjSAZ/VeqnLPBdFFkF9E0wgwwAV1/U4
6ERLn1RlzaPET11aDbjixYS7gaNZGSuUdpDDex7E6WhSmymZLjss1r3G62ZdE+5CBIAYKd7IDcbm
dLwULIPrMO9sx3bgil2nDskd90MhuEFjhj2vp8YcnRHDle8ptSMtu7rRvWATskfrtP97IqDe5kEP
0S1u5i7icf2bapYUQ5w0Z9dAhU+Cfl7borIMuq8oBSqxiOZFOe/bdigbELRMgQy7h+uEMm2QJb3H
m5E0icYxH9B7zKa1Hv/m/lnUuj1VjlRJ9xycp38wuw1uHGoPFCOCXVlAoKysV/O3+6bC4TwJOgzo
eOYhDleWNXdVDbOnvgRwVHOTAdIX3lD/5D21CjbWqgdO6/zEH5gAtWDQwgp0I8gMk23e1iaMOzzl
KAph9y3bPjKhXzJnRZ6vpvOh/DPSFHWJEYG3VuAOtYiEyQbFEbC/oymljddgKfCljZSdcGHvo5tU
9dae1fICWIOV8EQNl/wENEP45R0Zp3ZpCGQlZcF1lU73Jaf8uKsEgCMujMb2qCDDHvPE8YlYDMt0
DRMP8um7UA5tawONbt0kCILqPTCzea1y9nJg/ixK/SUxrgBd2z/Us4pWyLNYKAihToZIEizubVpq
BCUEY7bd36W8IF/P80Bpale1rZcBaxZguDVSOlynJeLbTrrWMi6oL4Uk9PO9CJJgjsg68upBJsls
9wwri+3goh87ZsFIXEd/uy/B0JAAAvzTFkIU+Qx1ZZiq5G42/TLfnshGvf377Da2+KMXH83E/eEb
Z+f20gjcb2104V2cIb3OeRy/KLaraRD63AZrOx/nZHH2wLtIIbV8jtFeeOOoZGOLEq6I1rJA6uGn
lAlGyDtTaE84tyRhM4QVxEwikHqA8sEM0X7pIcpnDO+tv6fC6f1WeN7w8/6BPv8af6RfhRRuM4mp
rqGGyapP/E5JDQb3+lOJzDSXv5h4yBrM/8TrmaNZxqALX/qUGphQyr7AK4ixohC8gTalyiYWI5qs
ng1UVQsnrySJzVfqSDIOZlH3yGyqFE5UoYc3icaqgTLkRA1gd5tnc8eJYFiU2iAZsVpuaBFSFNuJ
yH6DhtfwoK4SKGGPssq1pb8zGbVSZaKsMTsSUhJowzF54rn52zaiYfnfoufssY1dfxRcWwRac7gg
/FeV+rxQR1/L18yvBoc0HDvYy0r4/yaYMu4o0QrckJWXfQE7JdStpWShvA3s3e9p7iPA7cc8oyax
Wq9iQ9GBW+uVStSmoMDoYSC7Vg6olOihhiq+O28DkrD9tACyPEYBdp8nEPp8bM/1+6fJ2rH9rUlZ
ivN4x9TgZplKWnFjY2V0zsVSeZB875/OeRYcVDmhX0bmdH/+UtWagNhsXLQR+DKCdgf9ZgQGOBmt
INaNPkYp79FC1jvn4mk/H5RCuXQg7T+/GS2YxF0OdBoLdj/XpV4nvPMbg1ivz+3LXEA0Rv2ZcxyZ
HZqElXMkvTpxLfGx5xBPAK5cvtLF42gKwaGa5XD1my2rm0d1FuYYxXCGUVWYJW0lER5saWldd5Hm
MKdd9tpa9GYAVC9a/sayNVYSHkf85jRjhlHuMSlJJl9yrocrQkMB8z3oqkqBDcCxqUc79FPgwU+r
skX6+4XBf/R/cKb402i5Ylc3jaSMaeSzgwczMnztBx8vL2cRlZrPL4r5RjkFpTQGoUqBTKHkNrnW
SqcqSvBJ49fydwZTgFzTi8VakIN+o8oesUVjxnqyj94rubA8AB6wFWEcMo0W5Q5jVSMA1t6VPSzL
Vy5ZS8pzCZ5c31WYxZAjwvJn3w8EiHw/yFAtpEiZPXrqQXwx6GkTJCmHcBsBykbeiHXRsz4Xmt5o
HBks+lsYtbqAOv0b9LK0+eqfCrp6TFlD89ajqKx41F7tshRNKmYTLHLyFsQbKbsHm42Piu0/OHyv
DfpBSKIH8yqS/dy+gp+Z6aic2AdU3nvhezUjDKfA9peGcMndNBnJBj2C+DhR7MGsjItTs5hxfLwk
ZNvZ7BJUManYd5N46KEibdIRmx+KJulsaDEfoEO97uDRi4NQvwGBtQ1E6JjDSQ/hlC84JT1DNKPT
T7FvlwjwkhDznkXgoMjvQkem8r2SiQCoUVcYb0JN8Zjwceuz3ivSqhwB/jN5wfGW5ZxTQzbp0Zpu
RhDsK+DF1oqtfHvfAWSKhomkiaU195txh2iC/rs6LaAcYmk1j+ja+Fi65WzCuFH3Cm0mULMl6W/T
npoAw04r6C0Q0xBicdOBs1WIbMGs8uF5bmegsCFsGrg1icmIZEgTPFMa1kutr1ln0LbmTn5uyJJL
QqKbb2LMT8SkBpAJHcaVTJB3ECePmHgxHEqudz2YB/gX7orHDbOA8GGgC+kYb+GZyzjYKgRDFyJO
AeBdrp99Acw8EH+cJYSnozsMbOFs2qTxeauXNePqmahksiu8Y2Z6/B9Xqz8w6HAh+JJx2lhJwhsu
fgAuco4NxgvJTsM0u4p3GfBG594l1kj2oXneY9JpZK1X6Lc9BHf50BNvM08etjXS02pdd61NIVk7
jafsO9MOfGlVX3e9UhryGGOPiH4MLfSpWJBWGKJKwhFxoUS1JoyzYqJEV2MXHKVo6U9AWEkCehVb
QE2uTu2/AJw10wC+6Q9hP8ffEXlaRuUeqV4cabZLHfwj2FvVlOU0If+7mT9rIT3GLbsKmjkwbma9
Dua8pdOP06xs87f10VSdUn3XkKeTnStv2WXFGHniRkD4Ia8rneDBI9D3HHuf6r6RGGvthf3slkBr
808Wxf4Lji6mPQrYFcVfIOoPbCGNVSWrX8UANuXq5iviYjAVh5hvFOnIlF8wXjFegayuefSE7YOW
mXulAAc8AtS8UUCNQlqXHQGR66sQvXHTu93jLrC/bAKbXoumoUp9EV2bs81zKT+zyMqjkP21ECbn
pGt6upyZFAOL4fG1vfZpoG9O4fpR7CqmW1kA8533HufV2eJHFrk9K84FQJETN+DsPYhwVgTMU6s6
jOc6GFK3k7MVjgQLWzMlVRsuAMyRQ7+LYX8Y7njs15fmHPFbdPlh8aWKRRXu/Ea02r9GCxAORGHX
MtDQ3/Beu8VHbQT1gsKUbPMCPm/65id6CMlB50jDEzj69KrcbIGlKkME5Lp/6Xl2/WrhV3EK9UM2
UO2w+ekxXdJll/vNuk5bEcfYANJtHZhyE9+h7NTj+QMlorHC+w3aJvpkZ01xgqZi+C2rAjsFQB2q
vtp35yJbw+1aJ1xyEkq6ZAag1sX7nXi2jfUuSgK9cOizsKudFCv80UoKygH2NzF6xctiLno3suTJ
MeoadFcwPfyaj/xW9QMEkc0uVeTkRS6aNZ8BKxBZzF0A6jC2veGR+snsVzUxwvRh4tLiJmWFLoim
uRH/DL8INkd8Ag6bt3MVndSZIFB0Qwz+LLL9oMUYyC0j/QbrAK0D8n6pl6lt9HZ1YlXciElekPkN
CCakdahm7g7lhM74pOApSzpnVhIf7ojWL9GiRBJ0FuM2Qk/agkXRLejYtCPqHPa5ALQzDr2nrxnb
IUAz2wwn6fjYZpTLFVkctpMajA5E6KiMoXMmMOUULczluq0YOfqVOdq38i+otOJjKvaJslkG18AG
zwLTBQewJnVBlRWQaFGFwLzr6crdyExU+kwUGJO3JolEdp1qpICbVzNjNsiL14sfcyFMmt9yzUzT
q0uhiihxGTtzLaRGa5GE0E6sBTuAq943RAHoBCBA+Ch26woklvtBipJgtpZBBPhImNgfybQZpQvR
mkD3miQD2Roe6lANm6Kb5G12xC80wC/J0NkPJ8x7o1jn5g3CmgHQyJ7GmWHF2hGYX1er5zBo55Gc
RCt7pR3Arr03lxC0iNjkB6Np/9nPG/K/C9MDOdEt6dhoS52PtbhB+/gf+CZlslGauG/1+MHOIULB
b3R48+sV6t9sI/k30/3ojBh/37rthiTo/rFOn3QzkwV/JdLBvk5qeJvKeRxmolxUjQ2NLsnwmOaz
SLLRx30/0e7nnYEz48T9X2auVbCGG+G3e/rHu8U1+dl/R+Of703hDTTaZwYuLSCFmGBgMFEdn4WM
qTiGV3Qv3w4wNfQaXEk9vKCLI1RzgtFYQoqpD/bSLvTNxaCXJ3Uft79H5LKZgg9fIgxCidmCRki6
iJb5s0ipzzd3ZDrZZzOe0KOc+7CpvCyfOddOl9ewq54vpQjHmUVh723Kp0+DLMfC6cfZl7yB7PNB
uEzCyuBvdi4SyG5PbkY/XEF95JJa3EpltO3lqDFmqwZr72Tnzrfu+1nDX67qFRgpJ8V4MAFo8aiw
2H8T1eHQJXXcljA+cWzs/85RU4eEc91noyQI0AAyp4rBNfqtEHHdx6QFqPhKMxoyhbC2bTmTmCRH
KeSFHsTZuVeWxquQxOT2trfHg4pik6Xew6mBOIkqxz5qy3sOtEc3F5kDkH26NwpArD+Dti92lT00
DtPXwHjaA8A3Nje7nEdCfESWkQS1EwCQswUDGJOmHmX6yyHvtgRY1p0gvFlvOm70RwZD3leQg4A9
g/Ps3pH9sg5Ngt2e7U4mBLYL1SIQIoTe9VnU5HxMwwjTxWaf+fo8uyI8Mn/yXuLWt1sJ6ddoD0xL
A53pWzqFyBitCfpeSDAEN+7VsvyLJVKOBvmZhDkHHfSA3xN1mx2pex8AxukA2mM1z5D5S5TqqHkX
6GShZKmWpKoGBtFSSh4yhAWAv0KebRFB80oHFlT8tacvZN/dMZUwnJ1GxHFCiOLmbQktxZDiiwAZ
0b1Zf7qUwUXGD7kmwrUy3nu7FeDUUlH33ioLtqlqaxd0rDOENE7n+g6Ar1qkFumb43CcSknnfOpz
sabVE+fTjmDOIXPictis+Yv7Q33UN9n5kEfrpAu7iGkDqeoJkRROOJrMQxME0fUJNUmmDq3ozqQ0
gQwrJ9fE8+1zRiOFHJkFhHEdkTexZyvxVB4tXYcoEsjlEPI68qIgG2l2rYXzAFcvoyHugSL+gFfh
C7ZqUkDcwzLY38XhTnv+/xfpBHoiI7Z9tAdKjST61s2oVjOHVqVTsS6busFqmT1qf1gbTJIYDuY2
oGzUOiihkbgLTDnZZRuZ92hghNIhB6bBVoSoLWHZxA+qizcH7fN9pSxrTPKjRywGUFNdzGPTjU/c
A2YeZLDdOziUVpxDHQbLDCCTW1e+A6/Jl98IKeFEFRd2zG1vhTmVuK4bTRMEazwzg5yAhHRJnpPE
pkyGZowAuFcQRBl6XpSiJ0u9a142ejnvWA7M3bEKvIVMIj6DlFF0l8Bz9TvZiV5QerhR7AiBhLC/
A+bQSoiAGvHEYgLuxPOWMa43KbxbGYcGB7pMRkb9Z3KDAcRD3Q6A7VHYIPeooaKvVHw/4GaOve7A
6oGoEh6l8Q6frPzmSzYE7kIngrrS1tqjSUNWXagCF7e2BcO4H+p7egoMwirli4DD2ILr+MSvz5IE
kriromOJ7uZpfwR1cMeg46jpy42afUK8sPFxpnpT+pMnQdn8y+/zWPv/A6nr945un8es5EPHSgmk
CRJJT+FbRj83hmzktvORDSytO41zXTcD8aUC3dG7bTkFMWY/MEHQzmqt+gvnsgHFifcVs+/SqmSp
22mPpPTSBawVZr/UWXJD2ctD8tHAkIblU22YdW8+6kk2GbqUY334jE6XvznRiRGONj/D3USw+bDg
/j1Nk5HJwXnLbRHv17TaeyrBTAaXf3eZlZDJ82nlrdnKW0KGbB2DiFH9kqNArGcT3YANf3GxTQQf
4eTyRvlZlUZg9pSzAaSKupdG+ndUlsImJGnPYqyNZevoz5JHF7xEX+9do0ddxhgy4tKeIT9myVMD
wPh4aMsVrLJ+Izwu4gr2KSkezCUV6mIQ777LH7k9mtgyJm7+xsHKwWohJyHrt34D+Y8QfIIzkD3+
kO4aOLiPigczfAvZ4kI+yimu7SSfa3KnMpgRS5PnoMIx4otiemCal4SEbQZlfVqV3Y3noZ7mWLnK
S2cJZrRY443YeOa/EtimVyQvwvvJ5ppvseepCrB4v52BO5pLOZrfqA9Lvav/KMAtzUJyGpJMSnLg
cME1yRrfZpptg+7UBTnz1wbzR1Ymgc7VbQ5+9CFo+af3Bwm0ZS4DLXfAbtZwZ+HWmZjkwCuQBlwC
Ztgarp/1ebA1mIsT9qT2SmMZaEhpytg6kUtd4CDbo7iVySLh86SYHk95g1NDVu5CwR9YxqbAqlci
/AGoJSals0amWExtTIDzNtgrR+zxr26FSFKeMEo2EjO4gY6jYCtb7eM11N8aHbdQcI3meuOpLj6b
af/rAsXl8G6hF4RU7yIq+HplKxHRjJUMfVZyPD5MvEO0APLRe3x+bse2ftwmCBVb8xy+HJG3qccl
+nsZCOvZTR3jJ8fBcXMkaek7OPXCcD4Qq8n+EsVueyydRDlwypRkXa3xfbyJ0CKK7YTUTHVgo4l9
gh8t+ilLICWg9Ye0Zm30qaR3/seH4rvghQSLMpPRDpR7tCXwqD4DKKiuLa8UxioelFjk4OBX8AvV
FjtSraMYg7AxVlFIlKSibwpvoa8EV0rk/IYB61ruidM0JFpd2/vx3o0OyO+X9O9Droz1xe/TifRm
B++dh767B2EAWENV6jA8XfqzkO8X/QjNuYXZYsWxbWYTLTAiuyzBOmrQd4JMNXwsiKJZpaFPnUMm
xrnQ6LSOjAYf+f3PEy+U0uVoPisB7wFjM8ztpPh+zfGQ8gYSyPMoQUphrBUKl2cekun0yUrzLyd6
WkHa08hXi1UbT2BcSmjZFehNDdKGWMTQIyeSLVV2IQce3KGn6YBxZi6v6bDtLHs5V52g/1zpslRK
+deQ6V+T+eT0KBx6rjr9zKES2oAv6Gc08KpWv93Z9u6DLXURINA1fbGfHI+OuGWD7PuHrpr0kMhF
8mkRmiR4EWd7S1Nupmlv9eR9xftwB0VT3VrOKMxYk7L9oeaBSEhxiCY0DbBlJ52CV8XK52wo3PPK
+v8NmRa2jlPBMZ5KF+4RFt0PEltvcLJR6O5735SyDdYPY8VjVJlJC5jFx+vb4uj/pdtCavxuaZKI
fPHzZUYFe3xbJOvwR9zmLqmOAWNdmJ2ZwjbkZxIxhpYEEnrFgsmgIkW0iK8lf/x/Y0Va5LtuM1rq
0L/R85XOOatn226ivEFAS74Vks3dQnAfsdQdPf8zfy2URK/+lZoJizbU3VgLzolIcfRkE+xuFMKv
HoO4654GTg9hVrlrZqgflV0nfHVFFiSZmK2QYLCFgA96tPHxfEYq4gcmSo77AOyPcI9bO4WsxG5Z
Nh6DdOuUTh1hz9bn8Ak7xAthSQQgfxoADv/fLVxdcNUJC6LGRzTbWAMCjAtFwYQRmYKtRTX9yTmo
xL31GL8UCSoKn9ANzQ+Zo4IzZdFde06TeGht8Ke8+N/op9pKsAUPas2OjL+Nc/s/MLNNkP8L125v
ZFryASgLpgorE5ltuWIH436JjkXyOq61OQc1qdtf9LrGqcF3xIpz3S0T0zmZ2VxlXOaI/FrWE07Q
JCXW7d4M5NhwokB2vZvOW9IgexVC6kcCN3CjYcPsQQO/k+ER+Qeq2TqRg5CqLgXG6SLL7eesb217
WLqLbMcAnzZQnCFODp5LDVrAekOq7XAmg8NPNT9+c1aAhfaBSUuP2DfEG3jDfhHnTfXJPJqQcALy
+1WpJG+60gk8Y8aW8vTflWH6puK2iwFByGBOedUEirmeeGWz8n3djQcUGz9G5db8I97Qt3toqluz
BQQtK/nYHa1ypw/ztfCaTfjeBk+m55JzQgYEQyRpH06pvtuNLjbb8BcQXVZd3ZHRsWhCkRMyrA9z
fw2vAmnklcz3FjsQUhMSSuO8vwglGeGBRLYmy4MLYm58pgbGX8ajk3yM0eV+/mLRkgHKiG6+4Gde
xq2K7Pk7oTmqYO4+2l3orLIxnRlOeAmbJJyJfZdIhZWfhgm0Nr45gRP+/ryu5lWsVJifsqlUQOVS
FPcd80y6y6/EGLA/NvIPJgTxcAWG62WiloTPjzj/UrgdLNptVxFZxWqz0gmtUa4jVYMAVPQAIvSr
EcsrMV1G3ixmlH4y4Ovo/Z4Gxb9KHidfwu+PlNGnztecZE8r4+DNl6BiMxB1oSBQh2VbAmbmFClX
25+K+1Cf/ys5JE9+7udYtJNBkO14WZjvv4iWdoA1TOUf3dzoxg+yqMtkW0QYTX9nknz/O7dUay4M
3Mp1mwHS6bFNj9XjA2Oy4LB4UJpU8FKMx+IoDu10MJUIHZZIevD09R0GyNAr8OW4iaNiV6Hmcl8n
5dd9P/+sm+z7DFgyCtHsSk0yMVqIFiClQq3HaGxgpltiVw301oPv2tp9lINvM0R/yV5XBfBFD6jl
ol+Bi/nB7DNJGKt0I74RsAYdOTx4xEYIoM0HWWTB9AJvXp9XHYoRFKtS9rcP/vHp+czfIvoveYSc
Xfzp7WP0357wXTRjA5ZGWgpqabRTbWXB3HXGE43Kx2lcEwAswl2rCDbHK7UH3mT4Jyv4utvKHwn7
AHAu9FXEsQaWfN4FXJOP5lZ8cnudCoUNszuPt0S6HEgDM3EMeyLOKPtylG9qZAuQ9lGO6zmugmG2
AkzMgyLWty4+XJ03EqJehjLerkxUUDJiHLzvT0Mc56TjI21Xw9tOUnM4gCA+kSYYhw1cAqBmQ0ow
i5Nh8zzOk1WIgcsBdgRnelVsVyTxBXbsyyJg5gyIIq6q5pbEjltxkLYdDEkMlEr5oAqZ1/u/Buma
ngDMLZ/v1OamXkXt4VcZo3oPhM5pzSausAHQ6nnQM2gN5doG3nUwOkhEoKaGACXAF5Qq7yQwi6MF
k8rUpWr5A7iMbpS8MdMVeeXTMU+rxP8PclKp8TWWayk43vJ4WmziipjtXUiT/aHq8AM/Ix0oMirV
UHH68AFfnDiZCdy/TgucNrX4mVqYqijHlO2qKQn3xPExNdz79AZPTH7deflWr677csf4BhRYEK2h
1Xs42VWA/EvtRid9iWbvkSNzFph7DI6NtEM58PR9zy3FHogSCchSSk7vbmum7fADg2DklMjGEJph
sThpgbQSWbSqJPeaCzvduS0THG00LFsXBnJAE4pGasXJrYo3Escpr5CEf+vOY0qcD44MnL6lXSJ9
JRm+dVqmgmhTEySTtYZJyWdxClxb2f8JwZSvm/Mibtl1/zpn18pfLO6PWXSrS+UyTv6YqmozLSO5
MtSYNRK2mGGjIU5SZgMUBIJQBMsS6/57DxQkLMF003lWY5ZqbOe6rJL263vu+ViydqUF75iQ/zaI
ujU4x4XFTV0go8ChOth+VvPSO/zpkMXVC0UsMJnd+eBoJAAXt60Uy6SN0ME9CIC7iw+DIHrRL7N2
74ELKEQo0SSFp8Bt9uB+hu/ai3PzIYAlM9uo7jY8IFhBOBJjhueg4fzpqYQSl8zmLMWFJY+L4i4p
jURvjtivJhX8IhgVp8ze0VrRyVSXtppNgHCFyGh2HjBUJDbj0PufcAIrEMGXckGiF3Neb0ygAOdM
6Gt4gCIcDMUNecp4rH2bz7GfXxPUJJP6qCky8kPphv94Uk23lmgvN4OFkNiIURVZ0TdNCDqdhuM3
2GzAEuRDP3MWNwAXEk9JQ/vzmduEz5X+TYdJI3KJfd3oVgtzw8w0XK2U9UPsCRkPJ+V1UUaUvTjR
0+/ZmQmU551yn4G8lT8AiBnWvKl9x/bXIObT6xf/FI98eFEFWYrmSPWsKDWHIO6qCjSioJ4R0aho
GenWGbyLYM/H8CR8zMLGrgcd1Hyl5SQNUVroNaHjYUb4zhE6RfTM6+2nCozMk0Jhh7RYQrAEmQwQ
6fqmnthNUf5aTtMhPwXsQQRp8KZJKGy/C+7pL0Im2CVTs2M0aqVehHjhiMiMHdfk17dtN8iFgslv
L/abtZ18QBlTO3mr6DLe4+fHV5C6fJ6O6yHKW3ga9DX+Jb3kwbE2jg3hSYUL3b2ecrZnYNrxsEgf
zEmo4t0ZNEOwL6ouLv6aXWxgGCO2xwiHDLqZSfJ2LZ7+Qz9R11xVbkPX5wvDpBYJKyFNq0zy9NTk
POXZ9TTpN+h3qfaR9U+OGiA8Ihwj5nEgj1G9DLyfoSPqnq6u5+MFPV2LKTAe3uPFH9Iijbyd6usP
I2iYeVdkS7ee190jPNLrl3I814nOLjcbFL+A4Dwh09uPmYK9B6bnZzWnX2mN0WSK3sG0uI4rDJhS
0MiV7Hw6lGfeT4vPmSY85SRpQnUOUSoQD9jEUF7O0r2ah4pMx4R5voTMmv/qO7ED7eeSNDRgQJ8g
/e5k7NM6NxlZFSEu2JOVma6tyf4626afJDTx8jzQnXlvc+qGJa9YUSwrP+idZeZxCzMRVFFT5/mQ
4UxmpcQ+S6pti/OlRCxGAxgv8FnRTcQxjyEnPmH7AUEtZ4i+JO/Sb1sfBIyDLi/OyoovfodPz/G+
s4svLqaXv7XyuMPh6WUeUMwPRVCmcz4E9NywZsX23sqGTgcVITVN4z/0gdYLPdSI9e2v1jMu0R/B
1EVq+aDNHtMXpfm05WtoCtkQE45ndM93yz4DU6XZ0Xb5A2oWR/NN8VIi/yr6QWnJ8e8K239YNgdi
hSyl00EXCHarVy2UEaDaRTSNCcPHeQ2MtZDDb6D4SdADqGWjO+XWnWcmI7fSDPGrq0Bogk2VvcoJ
xXKPEnFNVVF+YyGUSMmialasCyCZNs5mdbLkkJZZgkHWo8gT7B/2UkEfC8CZw7r5elHMw3kcBTZV
Q3nxad1f2X+AutFCeY/A1Ckus6d4qVVVtcQuEuGIRrYjpBzcs3RkRdM2vtqyGxmh673IvSlPOwff
DM1zNw6xTB3mPqa3wk0ycSiVGvzuOmE1CzmMoKfkhkUzWUqVz6mV/LIyAx2LHEulCx1wZ6gRfTMc
2Dy8XYY3sibRPJnZi5dwmrV9WjlT6NHKmUm4bz2aZpeEMLGXA8bjm2wZLHMfyglwZ31C0x9sNviA
G8vQb/SeSDUCYFQsFfu/yrDCyFKHnuBblPIy5iQ3XCUSLRl+Rjvgqn26ksE1QXUi8UHfqRVD3iYM
NXXDowdUHTZ73sX07hAfeszRzL/sUyLrLHOpimFxIv18EznOszlkR2FcxTgqfooWS3Kj0LGvtb1e
+aNQbnq83BCYRd1VquM4TeOEcuif5hxeI2d9aJHuvG0MAdPCd0cIDMgrlma46kRH9u2YHYVT78JN
DFTZYxHHwkNBZ/EHir1SLldFSQ+IFJVnCiKOI/Lbs3m9sD2/uYA0vNSJbh3ouiXKGMd3reyr0LEs
kzhi6cTIMVvHLmqbUcB8QRytj5+thw+SyFKWkGcwI/YBS6jxejzSrYDGa3MxEZ9BaDZVjFOlDjh9
Di1UiyUexGteyM6tZj6wnQ8xyGOVPBzPKnpQEmtegpLeSPm/TGJOm53fJrPRg/+q0ShLQDXXtvQ/
AZwKTYKxDQickXsPmPLcygRYUZ39xAHZoTStjSTtueBAjm2/3N8vSP/CluAY2wwLv/eqlYDH8HfN
ouiycXM2msowQj+9CtcFrO2v3uZezblr9ALH/ZJnr1nL3f5g/m6rzc6hmIyTZ862rnlKFnm8iNDQ
6+afGSe+8A+eCIfL2r+E4TftX0o5d0RGnp5atV2jCTnVhZrJbcOwpu2hrnbYIDJbdyfIoWRBGkk3
3TEue4YksFLyW7p4zswDgWxKbG2Tn8TCwUiqVdbCYPyVZwMdSDp7xON1HE/32elDCiTAY3+mfs5q
rGsHHvGnGDUdr/sLccsDZHyY2eHMIIBTR+fnVKngSr5Z+05unf6f3pJvFxEOzZwyXTGokfoAQ6FE
xlNQe3hCs0YXeePtEFOsNqSqG8hg2KYqChuS5jm5f8L7yW7omNh4Y9/TegfJmFsVDj854TItmnFJ
tl1X0Xwh8zdeM+/JhUHIX/lI9xu7u92CKQrGzjkXzQCYa7/rAiznQDu8iLK5jNl7/bPdz33JISiT
Y/HjrlU8BMHqHGN12KiZ5ZZr7/LFQ7fKniWY7f53YreHvmNqIsGbSLSafQ3MDdvqgMIf5uHrACTp
xDdLalN4LxGcXoVo8p9qKNMzZU6zfxF09dPyTFzkFFjJJLtIVLWr6S/exq/5izPzUVXt2eVlOHWn
FHJ8ay3hN/cw5mSMpC2rH2Rbo7uNybLibGvbRL9GXLLaEcAZcG8x6q+7bShgrTn+prtEZjw7Iyve
u0szqSOgf1R6tqg3/DtECuxFuHCPQqwZsaBaiZyWrzA96yZNXV0iVGLX8Olx2gu5PM7LCbukkV7z
+3gxrntRoorzhiqF2IS9rL12v0D6dLZ8bgjdrwlVUwm6Lc4bPWzIz3v96BiT/Ab4KNqtbIVJxmCP
wdhFT+0v3WYhAKp6uj0dlqFnKaN66v60P3UChRBmd17NVccwpIMHnEql3mxC9BF705Rlz0TgMM1F
SsqAfUbHSTGDgLOYcb0rVIgiWR3bV/VtVAuLpQOq72Esho1AZ72sCaOiWmCextG6iWL16O2xfxjh
QkiNU1nnyWYtrHb3KZi7/DT8D/rd47Ft0irzdpNjil9cstlFgxwGz1GCrWCnDU6WvM/2ObFSTIr/
e0DtzeFMrJEEbnszdTarfLYmLY+f1atp7vp78CWtLFHCAsJJi8EBXMr2332w27pOQSQ3D1t2crUo
k9qJ0zLPq/02ROXHBm/PvgB8Gh55B+xqZRSCO8WZz4eJFFAAb0/VWL8kZpx75t2WLg0cvQwQeKmS
Y+Q7+TgRDwNGu621URWspLkFcwE/L0sjkC3IXONhUB4Vxe4+oMtvyPRl/N+QeaN0/eL1avy9WRO8
S0G9L4aIPGjX0JqLYLOJBVwa+mDZjDrdVAgpCLpiNyis1kuYet7MrTvE4jDcsB8UTy6xuRW6CJID
j4q+ZqqXmCxMzurhQO6MdomkmWDHdSUhIT4q575G21ROTX+I7AdPPyAzjZA1DIc6TiGME/a+9qYR
wTAQ5JSmDHn4VN4vxQQTqly6jSy0lHokU4tEtRjralGY4syMRWKlagP34YhOdKkcBPv9EyxXUAZh
FeJbVSHzW4zu2UHiwd+q0gzAGsh+Ynf43yvSri+wKNQgTLShhxN41yp6cFw6bEIsvVdrbci8UFbI
Em3QZHFD7OdXmG5fvwgnbp0bv1HJmZxt7XMUdeYFo7Hu9NoPNhxz9zIguQVIQccIRx3998ABV5sk
Jy23QI2iPEq2pLduOsnNKEN66Qi+GEH9XracbG/1dyhx7+NcmFT9XKXZzbHblqQ3O8bsdztDuRPz
oSpM2mH+F4smSBmwA2AXsPlHuUAs2d2IWC4JtwidtoF/lYs4qSuwvu3yyY3yF3O0iHJS/S36dUBT
91R6YI1e/Od/Qo/6QBdQFmrHADZp0wJsl7o62ejMsyiun2c7t0BbOrVqSIRO0IUG6eTwhS+UkfGj
7FkUN6xPNp7KM3W6VyzB0G7JtA/pDGlijJnrYJc3PDKxpvQUIlMaxb/qmBxl7cfdwXB7k5ARHAmB
op4P13bXWlN8xKhCfugdi4ZDGPOJm3Xv3xyv7Xt5wJcW2UVZ8/oo+mwszVgrCkw944W/M8SIKu72
0QuFeapvqKAu/e9q4XCXDNp+eyUl1C4VF5qZjH08DJAn/LW0JXE3i8XHV7UFqBWzBoMeVDNUNyF8
H4qL1ZVI1qCREGsII6w5/UUasfOzMxI/IccPD/17mIMlzZbYcBKIpxpY2xmY1+mGTD/WzAUrnFl/
HaSJ65R6vMlC8XKAphPre3+uqf/Ftm8zjof4Ws56E35Tefoakj3xMUc0VwDZDdDsOh1Ve1dG27aj
lhaR5J96iFAaKP4ypI2z79NoVtOg/JcTIgl8EsRB7NH8XaWvFCf8DV1vC5GFj3GHkbPiao7JQMks
RfwAjQtD+J5Wrk/+7GXpqUytgJAtwkwtGjB8xTABUhFqeauuHr4ot8v3L4k7NaoH6XRPL+TM8upI
JaTKfv30E45a9UBqrV5H9chat5qlu+CdB+DcBYWCL5PG6BvnQKXNXPz2IiBQ0TfuomYK5MYGodZR
nbVTIi1SgI8LuAOb0X+vLZGLmmZXan3IGihHeJyFHSsW2SYBIDOSQOXElbIwDX1rIaVpq7XDcjdJ
ZRA8kmyCWGYiSfBR+kZuG+hl85onQGJmytTctwpJaMKjyk9wWPyRxajwkkKGjglBgeuWOpxZAZIk
3RAJ+MPRQKkyJ9QWc5RAYI6dSHu8ebGWniIV8dGBVr07HUVzlAfPirwYBBSOZO/ig5z7Z7Xka3JC
l/A6cP3+aDy2SsbpF4zYwgldJNjFAvJ7gWtortSsvl9JVOMaPiYyj1uM3YOQu3AMXnX89NtIKtnC
xj+qMRXOZqbcWTl+6u4WFobzAJ1zpGcHZxVjAI5d26EaCdpC1YcIxy/mDFT78Qe0OM60S8Y2ZH5r
jtE1EzVT54vSgq/EuXJOXn7RmKL9fMOPVbEmkF3nal2JSrgz6XXW1eE97ZkPljxpihdg9nP03rP1
0CAfIG/w75R6ayRwqDiQ6T2vtRonLSH1r3KRcch59he3CWYIp4jLM1Cl7zGi6XNn7rU55UBqiAKI
5dKx1cesJKp9EMk4O3suttZC/FKJBdfzH9qzCFvU+Ds8LwrvsppcqQveQpmd0mKRyPt7tuQGkuyp
N+DmY1LS6mP+44L0p4Tj4j1u9ACFkB8Hjf4koRbEXiTkqUprHdDnjop5eW8y2dIEVCw27RsYWodm
4N928sukO47p9KLXgpEZUeTR3fsAz/C/Wy3iwPnSSlE/nsRWnG6mdpY/uitmIa4k+bmeGzvmXWgY
EV4bbImvM433aRG6nviD2IaaRfLLHVMLc7QOq+F6UkvFjF071Bz5j4Lu/s34fp8/p6Nckv77DEIT
N8ChMsQbVZ69R++BbBLcBAz9dG5tR/3I58jq/LJKRT26izmFNvo44q20jmqS7VeEdD/ey6brMofE
ftNfFZL5TUi8pHIWFWqBmQoQfrkvIFD5tIuAD2UxtS9nKTquwXLoDwyXRY0d2Pn0mCnX7e3g/14B
P2NvYyyi3Hoxb7ln3xgajlubXZ78wsU3T+F1ltwzQUC0ax/fCphrmD2KJwn7Z4VEYxO78ho2BOM+
k/h/HoUPhFtgS+k0uNr3Tuyv9TNmhYLyZg9ij2c8FO9EL1VAmE3Ezig4mdcSEC8k4kJgA1F5zi95
vPWNoLgNFitceVFGC+E4gEZRqf1CpO4ULswCATqdFLy3i+7JYahWOWbIiHIjWVuKKG3Jcy8G2Bt9
+ScT2U68lOl56VIZ6p8flTolH8oPrdDFVcKi6HLVIPlS0QDjqSvBbTCIxLevuxHTeu3m27fXZ99i
lCs+TvpOHYZSKlM2Jb9K3rbHMF5oKymXshGK43m7NLZV8dkvp57E6GRA+sxqr58qfbfkgKTkrS1I
YUS45gKjBxM0GcWkYrvY2hMXEXCR3W1BKpBu8O0Dt3BfkRq9A72d7h1qqhB3gC7toRfveQR7qtAO
fi1kmSet94Cwtyj1IQ2G6tm7iJxQVg9pG+wbvkX+0iBM6+Fl0sTrlKu8Sj0nxkOhipfHEktGP1sB
YSpdTRh8Vs1in4TOnAkUID9/vLn2/aYb4EO7KjF4VoogSOWkCXZHQTyvK+Bxn4b29gFnM1OtBzvS
DAUqUC5iJ0dXjqNM+yZCBGo2P5aJzOrQc2jrnx94nfxQA04DrDAjTM0oJcaxBB69ePYoa8EBUAJS
DwBLhFTmixSKlBgGrGGzpPIohr4Do7ctHwpOxa0xxfmqdqGmPfB24PnKiJ/HujYI3HvJtPG8w2Nn
YOyZT0Sun5pBpAHYzbLeH+ZJEjpwIgzQdaQzbEWn9AyWJoX9sugXjfmgr7oaCSlQjdCmUXaaErtx
y7bQ2E2FoPhSHQuH9i4UwWE/tNvufPAZb9Ag2ke95ffT9XHQSPZf3Ll/VC0LNpsZ7acTz3ipEaI4
qH1TV7bm8UOjKzCFdMgDRmBpack9D8TiS3qW3fgBeZil1jGjMJbHdA5kLzL5QYru5/5M4VHn0MQA
wG2np55oPWOqz8qTQm0q1ESWjxkL9Eo0Y3+GUbw/YZVX0p/jOBD9ThbfKn0rHwIEByDrvkjcTSDH
6b4STXgqoSvca9luoebEDmFSg2BN8we2own0uhZn7KOhNL2/+VXskqosLWHrQQUuMLZgaE226u3o
5Q4Gwn3kktQedGFdJ1cOAUbYhkY/vqWPufmyaeG0b4Cog+j7P+yGndjmTapxI3Ihobz6lTSeclPk
vrIVJfp0jkkHOVLUfZjIEBX8FyN3Cp82Y4+ubeToX8TSzTgA6IbwVyCKNhgdddXAQwGqvzA8MeMP
3OtStSvFMABKV3BuD94dges6PufJMTVhrpNbQ6vGOsxslUicfiprSeZgRsGu/JcgHxEM+5hdBFxF
Y+SRRW2vfHNfbdl5xGHAQXC4adZRLSXOsGkJMCWdbFF3ltr8sAxEQcJYsCv+Ta5WkMSRSmgVfBgi
xAUB+UPtdsTJiecNMVnCGbo72mXk4yfiZDcW6Kk1eWaMnOYZfMBoqxuczT6jQnanTDkbhq/qLaqW
V9RthBf772kxNp+nUoaNfSdGMAGdDFLE7YM68ghoR8WR4ur95/BrfM7TwHBNp/En2QvLkk4pT8mK
FpC6l5nBgcX11ckbYd6Otc/eXg0ILYLojdtWfZ4oGMcKqS8vchc5PRdFP2+dpaAwLdFcnPBTCk+o
XG/vjogLjUffo9Y8aTSj0eiQa8WNlrUrj9N1wCCCTfoKJauHZN9pvnyF+UqYmEDbbFjqenXXx1z2
+MMq4uLsLQ55WenbTe52A5MQwX3kpAFAx9N+HvbjSx7h43WQJffRkSMpvBscsNFwZA+KDMKU8sWY
H5plk4q7eq8s4k4ry8UfE3AlJc66GH5iX8SZvuEV6PZg2kC/NmiQG6WxXHl5ZO1fgr/cEHbWbjO9
hg7ZVfq2I6a3BRKv3bUFxbjxxU9lthSNwSaEIv7B6jb4tpOmAOpmFTBxSKfSv8rSrRG43lF0p2F4
eqdvEnaT4fajkWwoSD3KJm9T2qQ0AzFXK6CtFvkrJX4093KF0+GgWQaElXcRbVQz8vb/jtIp0Jtd
zBRS3MU0wZ2uAwh0ZCHxxK7eG0Kw5jMbLAEeEWs367ZLGLvkvjv8rIyUWPJoCKKmAmBlCxsDzUVm
2XzcW/VXiES3gLd7u0DyaEz1NZYO0Ojd7aMKuXYff0LcyrJ5g7wlQkIyNNNxRfcGqSlIAB3eLvAl
vzgQzEFMsoeKZDERyPgSzixd3FadUdN4ZP7LtFpHOhdSSbBdxMbaWKD2mIV+u6BQg7SruL7TvU61
fOsIsuZ8OBNlGlZtduYeUYEpDtWaGnpwgShal1oai959zIRtwHiQtm8R8a2kHWusmn7vaxgkD6+l
GexuGkPWR2OPYvorMKDS00+/9qoxeNSMUdkrNe92/ML1gf6jWRe1rj+OIGMC3KI104VZCUAekYr8
OWk6dgc4F91UTiJKLOOdyPzHYF8ACmEL7mCA1C73Chnbqo6rwX1CTLtvH8+7doUyJkn4O4Z9CIGq
sxWkkiVL72As4BZeJzUgPvUN454WQmCuel26VzsBiYdSyDk4AVOLuYgxkeZ7oBl8CR5/aDVHtisw
juXLHwn9c9jpxygaeuvQgmrl5KkhroMepuOKA/KHUgtAIcuOJ0QOMvscQTODp3xbUWW2gE6lPf+c
Cmpsg8daZ56zDPL9cgiUP87IqYE3uRdp+AtrgBFXfLiH1+XAR7s3YRTlNU2RdFsSkbsFIA9rXlQe
qxzx1mc4ujkMBfd3HYEEdObgmLsteI8iIlvGjLfkwnW+fk1jBk6heofVP1h4VZeCtc3m3PnkGBAO
i4p7qLTbD7175q3cINwY8dpaSf95mwkivoG4BF2b1zDDDpdazBDpjeiYOClaMh8cw0geXZCkE+RP
nU5v8ejL2y9oNei7SoUocMXBmyZoKkfmAd1aG4f1fKEtRJgtD7UBgu7IXlwLC/T5C8Wkuen+k2nM
GsWN+zVgirbgM8haIw0xCdXRI8/xbr86JjQQToWRDuh5DJfgXn95QIaT7/7dwU4ZfGfwzq1XAKED
nJ/XUEY9pxzkEGZuRgxHNibWW+RrAB0gtUEKje/7BsMEmBiN6cgZvu+MsErAGR9ViALxnTSI6/EI
A3Jjll4Y3Twx3Of8typ4hPPsr6okpPCM1Ezli8RT0L9BhZBtMPSQbN+yUIMfrd5rk2ikgjHwuJGu
XB+Uzsd04ghOeD3QDN1CEdm6iWBgcCMWk0TFSR7egOzXxp6r4ZYplWXsmsYJ0nvn5I19Lx4+uaaA
/7I6MTtgEp57vovwpgXBjGoNnzDeELkVVdTzie7wm629ym/uZ6zj4r2S4iBmB8lSQOx0uQSfd2P8
+oVEZbYkZ6OeWv4rkxSqtigE2Djkt4h7cUZR4R3YMSwZJ7am+1UqZTjQZOIWMVGwHt38aRL/88Sg
kauYaPuggAGkpce84UVJ+oAqVXrxaGg4RKBARuAhj3PTmM5kP9wGgJfTMXItA/RChQuD4xzFyNDM
BJI+rBFl1uz8U5LfEq1O+N03M86MBwSkYGvUkDhKDRul1eGNCHM+emXL4EwLB1dLUoB55/SKrJYE
IVrONuekksIPV15jfAN9c01MMGTO3qoH2iBvWnGG404XxVSUzcp+xghonzajUfGu0VZANYJw2p6F
2fEfGlZBrnxT4qVN7Ln+V6tD7wrPqOQCjvtX3B/qZpOt8SPxf5TPWQ+mleFRs60Pqs18hiAJT0cM
jHLXkRKNMxfmWgW02MpuMdo5+QndM4IlbikJD0TdKGEsVdP4lyB2dEo4xq9WED/+q3l/lztitJv7
LmfdtIzeWOlp525VFBYu8kNokvvyxRTxb5Bb5VGj5GJIWpbvSTpVf/sNuCEncU8L/uJsVVIKciQR
mO4VXAL45UEACVc9EBiwRMUU+TI/WkhACrThpv3wXLb0TsT+bwfcdxIeR5GrQI1rlFR8sYZkH89d
BqILpgvwIoEuI9Y+oa4eCQCS8TFIn8DFvTSqqRhsRS/R/csxJtGnMjKWqVQR0BxKUMAEZxMkYROR
v5lpdbUn1cFSpYHDfIbcvUt5vBb4K1HssFatski0fzthgVguoXwkDOupQXOffXGBxphq0X5svP7x
1S8e87KthfsTv/gRKGxmOZY7DnBkc8Q3A3lgVKdGdk1BRh/5aCEUTQrxbSULXRy/poK9JUB6oi74
4yzu4PbZNFVpf/F9GUDoyguHLVGP2gEsfv2nbGgTvdqy+7Ul4Wuoi07J9Cg4TVmvKd7Rtu28E1kd
7u5hzHF1UlCCGM79QkrDHUrVI3rW0+MvTdm+jqX23WnqDOA3zZcJ3jISQXgawvr7rCDf0QPgzgHF
Y1pFWar4FuR28sQ45zXxXOt//gzUO0kZC8VNrg7kM8AzZLZS1mrrPEW/FoSSt3nYPW+DHKfoLFTu
FJFfK9b/WYjqWAnNpywQGY92fVbpw6RcaZ9Fy/DoPczeXGgGukMLVf1KMimsrw5FvtHhfu4A7yIk
vJfoS2wXgqO7fRpI/lEFfmOLT685CcgtNQpaX8ib9DbgCQRJ56S4a4Jc3dWlL53vg2ERItZM1CNC
jkkBLnY3ZeZMFzDvA0KHi9WjRjtz7U4kidhgL0FKu17Y00l7xo/Br10lghmJ/o63+tFlJyoZXMKe
hWz2IT0zMC7nzS+d2zVB5ZWAia8mZib6brvewnsa6zZH8RVsOrdzVORrU1Hz3flnvYtJ/lHwRNyV
WNleN08Wf4UULcZJ5E8wtKqFg+EM91qLR2s3snvH3Q3Em2/sw5pPu5rpV4LKokf1m4Ic2o8sVHlu
NuW2p72x6X5o7MCRSy1LxWrn6OT+d7gtClX/19rzRr7gNeTQBYe3smoWKW7Sz/ab8byfjnXcGW8k
C3Dr0bTownjwWcyyLjwWfe69aIn+SbSiFsQ3PpFhIQWe7N9jvPBmsjGcZxJhvCooXqoE3P3u3jvv
dAN3dHPzi64AmXOlbfqk/pBksnXLgKloKTw+vL+7vqbiI6zvwz+/ub+u8YxlypNWzjnkpUW5xVOR
fg3e+B4AeIbSnxqXcOdJig3qYSQeo+Vch+JPL91Sg68JcYVTyyJcgm/iMxdG6KpEIW3Nz/9pG3td
4hSWjkKxSjIG0XHm1zmWqQjeaDq/oXHMdl/ME+f4nOEHP3WZArHiXJGzKUs6TDMoXEqwN4L8UzgH
0O7s1rIWNI73YU4DDsXcTdxPIYhHD9Nwma3brFOO68Pqg5PbR9Qbn5iCRAxejsciQU+ZFRHhxs5p
ia4EMMWz7R2ntEbSq2kcepPxD7/WFj4aED7G/6jg2HM7A0oznySD2CrVIYz8A1uEilWdXpN53/m3
oHNo5j9oLTLO1ruAWBROVXqzc7LblnySAy3JlLu6AvBa43G0WqHhpsivgvk3unJJdE6NlJrPuMtn
7z1oRYcod7CZb++r8v6JTUo/J/Z+INNY+E5JFrCdBLJiYfTzEWk3QX/pmDRSn06MWmFWJzCVPvDj
S8H9z1W4Bki+pK1eNcnHTvb7V9LrKiqhv1oGBQPagNQRIoA4597XGrr5/3haFc2U4QsLws163XPu
MPb+4vFnXPldVgoASjWwejgBFRq0ZFCRzpIYkGYgOPBQ9rwzY6gGwuIlinTrCZaKX5LqBd1MknET
UDhnsds2pktiRiphsMWZJzN9Z2Wjk0Mu9GOTG6SbnfLAluFptv9SjGC+KGcLp0bDTeXCi6wvN6Tl
3elVy3//Wk3MJElBZGPycZ3M1Qsh5dEFqcsdUl5GNtETkwncybluLZCbMpTJt9guNh7eS0pbJHUz
d60ygRAu6RYO3KA01lC2ht0hqB6RC7zVXN3gH/2koVVCbJ8YSf3XWQIBtKZjIiVqwLCZ+/MFol4T
tkqi2zmQ+wtKy+YjNmkwwn1Pfi+jA4B17g7h95FVcPYTXMKLz4qocPGlRgNZHrX/h6R2aqTiisti
4us1ylz6CBWoSyvoaNQzTvV0oFYJxzzl+/+L5YKZTo3OEsVXykx+eqPnplLqJy2Iwo7aFfcAou2z
wTPeCq7iCXcwLDIKgC2iLP5TtfJVuPzOftVrAm/d0muK0JU+9fvwvzrIVBMf6JiQZplql0eBgHqs
CWMxnCYEx+Nlxw/9Ife2KbBXSsXqkmUqN/fcvCuS/SBf7C4yK0qIkJy8fihNzimWVqSDu1y1X/Xa
xLXkIxGtTqfMQ28eMkccY/AD95fL8QmF7ae7zqZCQ1s5cBQ6yyOC91ohuZSaoUxJ4i09jw+CR8Rq
gjMJfHKCoUSExipF9v9RzhjUZOlJCGdseV/OJaYl8696gITOBX1/bfm/tH8erMzo9c2QL9IpJWS8
lsbdf5mVyoMQa0p3vKAxNKdaH9leOtdHGFkU65X3AklWNE9JuhBW2rSpO00hY8dy4vYSauKi5qzD
F0duyXCzAeFJZcLxW27peCb+YATw4rigr8CZ9uQN6orOKusS1tweFeze8KGgej+cjLdnDpuMc5X6
1oU+A6Ft2O2PkxSdeMl4ZxL+89gP+cx6xvnYbdJ1xwKLcUYFeyYSKPZ1i1ZWHwUbIHdJAKOgpU8G
k3GBv+UBqpWEtK0GmJJqTKlfIkK9x9CIVJkyWJ7kAssspwkOThV7dz0cmTQ8uSOjD9kHi6rbP8NO
saCgFjgk6z1Vhg5nOZ/uBay/247fnSPnyHEb8VHQScehW3H33it9LPIJ/4MWGFJmiLemvgJmCLvK
s+A7P5bpWOoP6xaaIDNk1ieukgPbImFw4tSoW4/ej7AyWBtFLtzf5EubO5GtBtu1pbKmu3PWEJAT
xA2M85SUJ1cQk3KeRZVvTd524V42uZQGCSseGt/gjWzcfrEth8NcxSM3ryIZcBFIMEgzvN+U197+
LPZgeqmq/JxGCYoBWw/ZY62aRl0D18Anu5QTfNsKbj9PRI9CjxHTd/J5EaSCW6kHNkw05OvW6uvb
6leKQV5wPqx5z5jhph4xI/Z3PcYy5p5jK8FiR+1Yjh6XeB2X40t6Kc0uMMsYlsqzILQYZ1OnlGWa
fhfGQmbM10iFBsRPI7na6YVWJwLiVk5Zh3l0VUZ3ojT9rOaLnERg3h5rWQff9+ZO1zrivB/2Bniw
XxuXCc3o6iki85qBcD44ePRL2kBdm73ON6kr2mfmVOYffeRVUTW8MtcVum7wEduN7WKvHd/Y7rEm
ZG9SPjKa1rcRRLIafwQvvVYxjjgSkFQN2NGb3eO+Va8HCHiqrBhEw1hVekgTcRXP+2bpQlu67Csm
rEQJ4SRAHoBPOhIkhU6Tg+Vcip3j6gzpmRCs7a3yqGE1dikODrDjMQvjUaI4D3V81YVMnaOdi8pJ
TL7wknh+WTOM2Tf5p/8yElpaPaOyn20xI39JicvLUIPN7UvApocFrAeX+QslemLWXFmvWjyWKk81
9S51fzIggvhk7a6425jelyZQLaJM/ENXim+rpJbCU3sew19J5C8flwchcAys9IdY7pej3AZ7YwWX
8fOft+M0OwOlWh/1O/pzAuUfIvAPq2zQjBxnnR/7oqoqRUSE4tLWFgzPrIJwg7lYIyr/4UzvIBvZ
SqCdt762p0yImjLNOBGkNvIyDWSp3txK5JYti5Tnpdv8EeqeUbTzQVnjpQwmol14WIS3cpx1gYE/
hSOrX8EPi47EGQtM6jAB/EJ6tqLJSk67PRG4r2VrmYPwnjENFyCU3eFCCcrFbA66+Gm7R1jPP0m4
E255xjwGgtKiwlz2cYcgQOtSgQWNLP13TySGMhVJ58FrhX8NQZJybXSPHqlLTv1NosG/6j9sh1AH
INygtnZHDkaUtVU9P5z9kn8NYyqxmLeKF3popZkuZSISgTFXC5JE9rk8YpOtzvRwUxqok/e5Sz5n
KFAzRO7ZIivrpEtm7iEP26Yg1UcTWX9RBIG32E9sLNSiXVsZmXWk3dl3ITkbq3WSIjNJc0mEjeAF
Gqsh/VfIbAcQkGxc41ZmRbqWOHR4QWUOQLrn2zcCcWP3Zx3N2WSP0HWRCh3TM4r/KC+bAl2Rqzwi
TL4BAoVyWh/mY3oPRkJX0u30C1aQo+/n4jNQ8pHepvOym0LAVz3yN6K+W1yDE1roAYa/Q8LOTU8R
4kbsUfv2xs5yG7Fy0yqeXBEfHmL3saDBZoAf9N3MBziRvnZwCJRICYwjSm+JR8FSlcjQwetpEgbk
YsZ/GqG7ki7icDehBTwtk/4pO3CFemQ2M6X4XZVxV0B2GidAGsQd7Q4XQLqyHrp0cvfQukIxIAWH
hnRbokb/hDomU//adJS5ZPkhIt70EeJa4sSs7CyGEXuQoOseCdadHMSmNqLlnx7B4GzjXTYRPLpv
khKQ8dkQo02e/0p1p8WNv9zckmLDkDBn+Ip9V5Rf17q352iyzbHPCJSj2/P1lytihv8uTJAeo5YP
E0DKwiFZ7BaH5MQBPAeO05FTNUi1HltKQcg5w9YBtTIpp6v9ciQF1YRYo33biNndkl+ledsLbfWE
6o+QxGZf0csQY2MkRn8+W5JqjGHUHllxBELk3cyZuSINuzIV2eQy+ZeJqsH5wNuvum4LU+PX7hgY
/Ze2SKBXLFNci1yQW+8aG2yRDWp1DL6c5CyQL4k/7zyfx/JhthZ5BLLYd0T06KbC8jjjH1sBalZq
NpQQGuPnfEh2VJXoLHQh0jR0xRZylWNIhrhl/KPbIeMgcjDXSNTt8iaMRzB70d1E8HARzLNm5J96
nZWQTtQ+nosddPnFylhi3LjZaND+Qz/cUdNh4xiehXxv73vyHz79iuHeIZ/batutwR6z6FZ8jDNO
sUmQo5TlTmqBbTgvDfvo0DsqI5AfMouu2i1Q62GyaqdcqRyhD0nX6YnMqJfMQOkTrTp5W1Bc6FDw
i8Kn5tq2yMp9glfcoJO6FE/2+0hQENMTjdgs51fglDXmgn+vmfJv9kjHbc/MfCvHfkhvC9FfvNK0
zcZtl3YHShoGtzbnRtYSpcksXy3605hnaz4+kly94zO6s5JkAZ6bTSQMQLZ9CMsn/B8+Voc4Tq77
IIWRxSuqJ3h+R1cCTPCACN+fOyJUf4bUQYIukq3UeyeNCufAGC+7AnlPXWRPDbVhrCAisZSc9EUU
ULavMTupKzkpBB7RiucPJPOHrlUR5fN2WF+Kjs2vLy/OCAG1kT8e8mrUU8E6+gp4wp587uVyXSpw
O6BI4kkXm2tWT6ZGLX9Pbm5qi1fK7AAbmwlsBhSGDnuMq3epdMRJ31MSaNxbWgzn/0ZxsqR9NtDo
i7hftD4UtsdIqKQUeZqIYNgWYVwQigip4zkoZWvISdh7NbV6tnx062Rb97H+wdKmzfAFHaD6b1zf
qqs3bKAje22m+yKs7Lwq9Z+sH7rURntqaFbVCfFcrs+7fUVrTsY0Q74NBUTAQXqPlC1z4DcZzALK
oYEmd5foU8HO+72+oDIvf9fW/hsp9diAfBn4xiV/1/oM6MxSyTvT7PyBoZ+ECPClKx5vT3yPqKEP
XdWBlZfsRpuhwRtgAGQ5sWi3Wvi7P3xFyzXPTEENvK4QXijzo1vZHtc1L5baVAR7Fu+ROWg5zEEr
wzp+O7XncghltWsqbmysCeCOAKGlwkgck9K3HtkSdfixjBdfKB3sgsjYXFdhxCtvIyW0jM6kI7+9
7O2pELLXq2cHKys0JZ60tgsUHz5iL9L5VrYzi9wfwKarHLP8ECBcARXJJaTNIcaG16WTyAjK7jS9
R2ha8rdfX/r+erjIH2tCP0eE4iT4x5r3uQpmwv1VBUSYDcnK8kcQ8NfMI/ZhLnuAxHKqfE8TO0Op
z5pVQx1y6hK7ULqHrvER3lioo2xASAnZLpLxb/QWvr9GSaebdoZgI/MUbkjS0xSrYQ95qcRdMZSU
zxGy/mtvfsXMEb71FZwELwP9ynS8qO20uuFgt3CVerGLDt56WXSZjDMns20P55ndbajBz0Oi1Q2b
cLSCeiuT2I67rykLuPYDE3srN17u9C3Pl6a5YjNH6YKZF6nGSiaMt/Z6VSu9zyR/k8JzNCjb4Egu
M5X44ROyjZTNGgudEeyYJzpx007RXAazK3YjhfWNO7Oj6jrVChwuyN2gb4ckT9C+GUHWslof+Ynj
axrK8Ibq6o1ZUq8TemTku5+RIhG6bn25x4T3zkt1WXqP3kGkIqTjiZmT9rCuWWM7matLsTaFfCE6
vZWdXskCCFdqAG4Cw73P4IJTHhnTIiOBq9M9pufOWein4kylIXFl8s169ZDJ5QlXltOhkzoyq6Z5
fXXP9JuruJx6+nyz9VqTzHMnJ3ow1cYSpm85qKfP//zKNHJT9Z3eJIEzFg6pR5PeZbkbc94v/oaC
wl4xH1aDo5Tfus0NxDL70NK9TScKR6jwEBI1XDZsytYR839qu17EekZytZzbIf/WE/K7KrZKcPj2
rxFl1GYXY78UQG0tcXYBMyYniC4Rslfz81Fkan93/y86OD/YXlHuqV7RomgxiS0XAbrmBnHU3CuI
EP4UpVTBOlcC3yAFdZI8ev+ieiiNNFwr5YCFbtBXLEpV9WpK4pH8aMgSIhK7Zw97rkXJIssYYyLx
Aee4KsmahgRXgEG31aib+T2PPjZRPo5dr1C/swHF2jmuZNkIo3c9MDk23oAMKdHa2HvtXPwfa5x8
08VJqeVzgWHTSf5F64d3TDPLtK86fvJfQ7fI9crKIZOtw2xvr+JLal3ZBoMpLChRvSdLT4P7f4QQ
w3ksNRrOu3MzHAVsb9yjCp3KKBuqCEjl0VyCWS8Edny4gM1SGY3ZB2moNkWiL81kYxcW2/QVydXx
7Ae56l1os27DwBkNvzEceObBe8ThjJqAIgGAV03F3VzH4pFBR3Be9Ii2D0D6VVokuo9Xd1fFiBMJ
Bi+vXipoJDOkdzJ7Rudr3s+OxczuKk4gGW2VwTzGNWUN/bRSj0UqMZ7FraEcfhCK1FLBd9PHqaJ8
sIFdBtiCimJ9Tp2BZCejhGPzVkb2DYMOOF18/UXVRIVP8NavUxV5wBl2D8WWAetDnjt0uQx3T0r0
81KvxQvSNad7p6XqzbMcpHwqCoe0cqJL0HSskXyyh1rcc9aGb7AgZLZhHTg17nNvvLz9Vq+EkrqT
8UMgRV3zFCtBB8t526mhAoD+WD10r9H3LhTsK2V3yGfyI3xn9Z0p1jtxy4XTJoZLoJn2BiGwk2K3
442I/cKajIXV21HbMWP5/uTq8bDn7pUmtp4aWg+Qz2yEnhti+K9QbR8WqN094pUXbg5TBFi+IXSc
zW5wU7mBVLxtdfDPe5rQrNyyamNC8QQSt8UzpgdS0xHr9W4le0dDPDZsxvbFtNmaI10gDMPNe1P6
UxCyv6EQo/oed6Orb8Y8sAEx5NhM+ko3HlIDSG3S+0Vk7jrp9MUrUsnv3w8JdwWICA5lLlS2yJb6
679KYJNaU51qiF1izPQBJjRe+0lyFt3q7lm2hXJy4MmhlZi3NL7Bm2BIJi7Ekba52SRIJvz1xoc6
m+zpt/xUYsIW7zTyOdNRS+KP+TlOdpAgHY41U9RQJn0K0rEOO1uyO4rYoO5WDSBd8LHhPl5F4GjZ
x2QMzKk5Jm1z8WFc9nomXqmOZvohYpINeNjq5YIJ41aa+lkwgjLcvWfK3dZY1jePJN8pMsJtMpaK
Hj017pcAGEQzfnbOuVLs1hfefy4Zpn0blwEkc7tkWkk8+9Mn6i5iatlXYFVV0TLSpSyElxAQY2FN
qhjGj8+U7qb8a/hK7VbtY6CDX+g0BIhSPI/KX9tOXZT7iM7YkjC2N+61PTLLXzQ7xYOB76GgvSDE
95qznLWj2ZnqlPgx0bQRd2950ORpQIxXTn57zfSvJpZWP3wfEdpNzbpkU6nSSNqhPX5djfONwELK
uedUXg5rk0FC8n9BJWvy5lZKcicsuz5ERstL4wJF8YhbXtnG9S4aX7q2p0s9H0/bGvIK6QnnNau3
TNRvHsSolLtlJfJ5kaLp3eFm/NINr2hem9BolnW63//MZrywkgF8hTnqmUFKcs1L6/Q+/jffVG5U
5cOeBBJrEEiF1p3FUNCLlBDyQK81Kh496zF+/rn3wt3Nzl1vOKeOQN3n7lZsAGvw50sMRnGjD5mY
9TTXJBLfoBXwXOmVV4YTamrl4yIdGsjWsdrQ9kZ5Mb2GGNL6gqEQJTGxkGRLwfFPCvZlJy0N+Iz2
GfzAln74ItZjNwdtwj8JdLqOyrWHfPEQ5IaHZ9mE3SjltLIrPqsMdQ/fbbFea4Er8nzlnCHfYVfO
CjjC9lK/hTOJR2O/P+eSJeQ+lOaBu68CIcYWjpVMBSpF6Z9i9LkuOLJqEyasWo6zQmgVDeZxUCKQ
SNBd91Q3BZJfEB2Muswa/sVllNn0rbj2QSdB/q689+zJhDZsaTTC8Ox5gVfIaDuQWkmzg+Bxpu0h
NTrQaM9GUONGcjTTZL2a7o9slRpDIjZcF7sfVuBj73M8rTiM8V91nKCrw7xAlJI7rfVOLYFDJe9e
sZlWQuen+PAOtnAejShbSdTMyEWufQUr8dbkcsOW1lnjFROVM0/OIuXBclTuiY1JOLt0H91+1Lb8
0GQhmnbg/x6lg2kXOe/WcNycWQVBWSufH96lcM/qii9krCqGHir9rUw1f+V085oA4S7f6w49wJgd
ZItsuZxROVEd/Dm1Q8Me1518M+mEvcnYKqVWgcqdu5Szg+Uh61v5wc8RLOixcJQg4xtS640aZtfy
r3u31oN51LlGwBcFsXDIYR7a+9eY7NHHRaUQ8vCxfl4LPZmZ0IWzJ+thEYHyqU1cOJ5yLuVHg9BB
7TBdml5rwJsGY9X8WVLMCsc5dfF6D8qcyh80JKdwrfRaTPOfP0e5wufUgA1Q5E81w5kKorTa+z1G
S2upLY4yd5u5wNdvk85CwcKhpiyJOBlRHb7PzTS3EHwZO42CpMzUC1uZfnrQm6lxHJrtKPWqk6vC
h5b1tWRhBAHRJevfmaAUJYAHiWse7lLDynWTngSNaChxJINxpElU2f/OfhIiy/citdpn3/Fgh5sa
9Ns5mxiormhExbjIYId3BKMtu9qWVheTI64BCi0rYUUwYJy4SpSSJlPxl/oER26A+7KeYxBAjznF
jD5mRIWanhI8rNOimgAxpbx4TJbBn719DglSFsGWcw++Yn9/hNVloqXyBCnbvEXejFydvhxNc8Np
bQh6ucfr7H5M77g8R0UWo38UhS3khVLcKS/seOnIyS/OqQJkX4KLMySqUCPmxgfDWOdvcChwn4So
FdFpKzABi/yxZMkhen0oIYmcSUueLktScwfl8FdKihStSoPtU7wjsuhxXTqzaKZsBgcwsGRf0iTd
aRF7qklyBBVNJ6hJw5DnzNUlVAM/fJzai7mPBenRk1C5lEA+m3uKGNz6QY/EDaK1lB6LX/qC0Vsb
1CBi52iwZbdGH345rk9CoVhd6RnRHdQkcd2t5RBP4tZpnmPdfXymULQSZh6GLY3t5W1zv52Q8okx
jA8hkkV3JxzKiKVhoKS6mULz6qh1UdZNv3OphEzLMUTQXYczdoxCa5mKB+u9lceUCsPOs86rAYGb
EtdWSmV5nU5kqJbVPlPWF+TuMqw81ZYfI85C3SyUs/padc3csUPdl2WA83fJQH81j0o+4eN0D1Ls
xm0ZYVUPfJbqEixIQf/GMVbDU0FUDgRIeT4PiaW0V/tG+dNUmPxoR0V4U9nYRNzkkplQ9848mWJk
oEw9Q9xy4ctsqSkuqoXQBddPRUTKXJ9JbPG1SA/TaBmT6l251yZzqJ9kI8RhH9D0hWOiEhgQAspT
Y03cxWasE8vwMMr1v4IAOYbaSyJDadQEF00kLJwgaiBvaOj2Q6z3x8YyaECg/UmfAr5lwfMiGuli
CnXAWO0hngsahyS4422SylsQMEz1bjCVaNX7Xs11xvZTlKWz4f25UI+cfZMs5GmrZlyw0m82bZ/y
H4hn+hui65VS/e/XxqP/EkL7RiUhEOYQ75iIOHIgAkJCeta03c9QYQ0bE6CcG7yQEllQKtGgjSva
DYR0cWW4469er75m8qXXRu9Ia4GEiXkkyj3kNj03u2a7fK9vv0zuJ9ifJVT6eKncKPUSddla+Mg4
aOavUDc2eYgBiggJ256ixQ6F6MkysJ5oCOLAb3j1F4FsGst83uWVX3/7RzWXcayYcO4wPmPO0C4v
GxMhqL58GbBReQceuAnzmW/h8nIw6jwMnXzCJAhr/rgJgHGCp9pTorLcqaXlxmtqD8mVd30sjBpE
ItYi7Sqw5tPkGudZhK0bDV0eU7zBQ7rJd83HEnc07y2Qrxf/5Jo52pHM3OKDvgzOadOOrIK/c8L/
k2kQ0QqL5XXxkKx9gwlnhw0QrcIuKrqqvBgXPVdqimpbrutVCc3ymOpuEMzhpXSYJBZ3ybS6VLV8
IvJNRMgf2nCpYwUn2wf6iPV95WiMNNy5Zt4ENbgIvDOtVNjLw0uoylNDbksQkWkFntwgl8arPGTV
9fecIAcZjIgiTzNaqxfCVo/ln9OzosSFzfDh65Ut/9O2kyowOXMPBYmdXCjy2qo+Y1CBVYq8BrDa
xTTRcSw0In+NjlE1OCZut8RgX/S3BQNfeSiFSlP7U37Dmha+dIYKnVWIBQvpj52HS4Yy+UtY4PM7
SscpTmKPy5xp7595T8IOtMavzW5eGHGaAMbH622DTevPHuu6fTnEtdks5e73b18cnBaGnXXlQBGW
N6wRPZBLp0lH7Sd8YNRzYwyoa5NIZUens2LcRejPPUFprxFj0C9tQdqnHL54eCi7znBGF60LpAYx
Ymy9KoVanMsuqdBecGaAZ+jTpeimenUfda0sZjbnSL0F2GYMOpRAiTb+iN/bqvVgrcNd4oSgEwWw
DvJ48vyWy/oiKvansA7lQJWaV8FYkJRbK24OJWHBVEDHfLbdN5vrFIfv4SUXELJC0wme4yCFT6vt
O7IK3CCW9KMNE8CjNMlTrN0/XqH5D2T15ZuI2PrDWNDqX6dj7/U0bMLQq8/w8jrzsqT79r37lCFF
y/k5xlmncYTD2yvOGVg8zY3ry55BajCdtRH9hrg9Qx/n3wQbTW5of+qKX5Xl78Nlg0NBA+ZnYpeE
a8Ix9NprkXAbUan0E7GJo9tNJSYuDw6vZXYBd+CxtMGVLEsE7mouK5i29j7mJpopUpPEYsDjpT0+
ENzSH2zxFgQqXxrq+ifHQ25TiMhBNbfeXh3+U/BNq2kxTFYJa3ywR39TVp1KGX3NDJ0IbAJlXcvz
cWkN/A8QvydfpY3h4ViG0sDdhX3k82Wm8gSUE1ZCGMpFtfPprD7FCN7ggONVOgQJPRuycVwbqIaK
9SVS40CbL2prvzVCtlrkceGb7P8j/Lr9DmFFiaXJEXKmaTtdVtTyQaIKD/oGxtc34ifUB5Djwqqm
d6/YlLv+Mh4e3YzqPI4GhxoxrP/1s7BH98KJG+9AZvt4tNnEe38sBLDmhg/fz+ky4iESBxbCt4RE
NlSOkfF/Evuo/uHecdBbVmHKtDfhoYHPcoXGLt+VUwvvAGNkm7scCRol5S8PSkybGHm23ptPyKav
3bg5brEqu++cSaiFiEz7npFKEzsnMVad18aEyuj42EYRmd+CRZOcaLiVs/E9yGQeRfNL9GKx0pqj
tLqXdV/vkpm/sruU2wDMvtWAcPO1d1j/jVDoNpmngK7yjWsaCXXD65hCGV65mVZ+IF/H7FCaLKE7
a52s8DKnBKtMDehp86nlLebHEtQd50cJXSfmRfoL7NM0gnNLG2aZU/v490iAzS6RXTdACTmSuzXD
8ywnOOL35RPMxaMiaaxBuSWTPr0tqRcAgkrD2YPxlZL15Xl5qjtmMdQQdbQX788ldaPgxJ1eWdZp
i2Df1XIgcn5ScjNBgGbAWEnAhZHrIyJ7C6vS7rN1Y+3bG1H2+kiEgyiACLPICw60L9zLY4T/2DAv
cBYcUXvBRvMQieqpN0RHQlAp+NFTtdD78QRxe+iU8L/AbssgHqUVg1P/EPKol7LDDRph8/V/HYKm
5US2ELfpvpGKsl112DcRdAt85NLhMDE7FBG2B8uZh67+Wm5VsHZeBC0w2hhe2CcNySPGv6Ggjgrt
pwViASl/TlhjmW1VGgCk+sEwCNqCFnc4X+7iM6uOgGETv4RQL18hDZbqeC3e0TIiM8pVHG6wAemt
OH7pUSuODsS4fx0mvvG7yI/k/Gg5wwoaNfWxFFYcqE19E1mt3xLDsH9SmkOeJblDrbqVFgp7DOUk
b5YQcTwZtw55oMzDl8sbEqTNXCHizLkQF5Tq/Da5DJuV1q+0lcq4Z1sKK9imISUl0UB/GuPNV4Ip
ZbNHvV2PewhsopQqLEcGN9FlRXy/wireICUowqTUaz1BIWPSQp1yOv7b0rWYbXGy/27RaQ3n6qOV
GLDmSnbsEL3XjGYhoOY318O5ae+2Vchx3FP62c5KuGHBSbgxjbcTBSng8mIQkILYOI5a3X8pB5gR
9AEq8xcS0cbpa00RwrgQqW5Hvrp1QNuhWV89Z1yQIHakC7OnER64/RYal6kCvXYJJEmwECs3fhU6
d8SWjGmFdgwkeVNfNdZM7PrxpPvklVuEDFLOv3UpyGxCePxxC8f41qT00o2+Xb33EKrunun76MXO
LYYeikpXurZtYqq8m6mS05ewG2N6BVXqOhVMFpnK5p1cMeArFjpxcnOSZLV5lBSji0cY7cxVgKoR
V9K8+4aPf2oEus3SGP83K1pRS4toeJNhn/i5X5PsA8IlyucHM3pbXvPI7kkF1ttaiY0xGvr9A9EZ
4w/+3w/RpXrvAFzt7QCIroi0dEPrJKjMUtL6yWYth/ahntoOvmC0XfBq6A4Yg2wRThCo47y03MYO
5cIQo0L3cUm0KPnaPLfCbVkC04hxv5M+jW2SEEwKPlBLQYPpdrIkak4gRr4t+Wd2liqfUUTN6kgb
J1zJuPAr1Pt77/dhDmy73/i17HSay0n5FZuHYVsqcBpglBF77j7A9bebBjft0Fh+yzPGOMSxvbbS
bxu2/Yc4x3H/g/UErUKqIn5N0+cu7fYDmY3IqrW7psGLRB9QAcmkFwUX9BDjzhuGdOFYinWAoH9/
fHunEI9ZuvqDc6FGPoJiI1tWxCJbqj0lrSpYUoO9djwM3iCg+QTSb70Is6W07EQpizd0cYMcxntL
UPMuTzNzY6lJRDPU/G6UizN5o47K1X6JmuCZftzWdOGLPCa/hfMeiiFkgI/7vZE71s88dU0MeEWm
Gt0XGxWVIwEb7+tj6qJMHbQAWGDPqk1mk1N9Cnz8nu8CudGfa0RwgHL/URIt+9h+zQIku7PMjo19
xoapTor4W20Jsj28QdBRZ6TJjxWRo4Xa8/4b+qw3nhZCR6BXBTM1i72zWFLS2MHnbZqtdXbY67xN
Cmzbq1MJbbnW8bZVLtUu0aCs0rqzdJDtHtPpnT3nXAPnKvCICSGIwoWl8AjkbVlWaSsG0NJ6atBX
Y9DmcOUxy2b0v4G5H7DXxStJiFxjH+BoKEbJuLeKuvZn1oJSYDttiKFhxF+Ss6CZp5ZS58CVofje
/nY5ONDSdJ/pPu83rq+iDwR+5wqjRefHV/Dgiyr7j4LKj6C71ja3Qg48UUnVm7DKJMkZEwcr89s0
GQLVbS6guIqEFJ9jN7PqOZ77/59tXQAtnVjTWjblH8cTnzsXzI1OYkiaVX5yAQDjchHNyVWCfCiO
KJKhE/rVjgK6znKDnmVYBaoktln5SUFQJ/0GfUUi35IDGdNj4hRR+lroS6JsmMJntD3HR4gpf1hl
Z4Ywlxe9UrF2CdjRZKLrFxOwhqRa6fmjZZsJ4kCeUA9+g++87Hl5sX0L217Zfc7pUQ5JR/8NuL9U
GEsEQzb2i4LRh91ML1C9uaskvH6WSGpBnD5JZWfT7ZD/gMDIlp4ZpmhG/pbGKLudKNDw0iiUGcik
ib8g4k91TjNJOD5EoLXWMQ1dlNUuQueQk+vX5hZsm0Yd2nzC6ZsGoGqHzQYRY4It2oWMELYdpqTZ
/KZyOZalq0ypQj8MgwF3mjFcsdUjMvYF6XlLD+BiekOIu8IQlcnm2EKkpi1zJ2lT2lOX8WJYIbye
/gF+1abJAFcqHNZSxVHt9DGVsb8J9btgP777igw2+0qTPqu4b+jaKgtRagu6iF9RFe2iB//ViLKy
Wm0MMdc3XGlqeH+0nI+GHIkWFDDxL8Fp/MhBNuuA8hYUr8f6uysCAfl6KKH2w7E8Bd7svK+uYlm5
1KS/HPiqCXVwcqBUTYKZYU9dqL7ovIjxRLzIz0Pft72yE/j2N5OCtpqyUfFuDiz5nOB+nDHydy0v
UB8xF2S8S3XgcKPvOQYxxDryoNTyWWXnCLs0lNalPfBwmBq0QNF1+SI4XDX4wrJYv+WbLDzcxNaG
5HD++7/h3NlSySSbYzDU7NZQN9EqPO6RUrm9fHlpcR65yPc/eJQ4A0k7s8+znXke2Mdc4Nk5VGwZ
nzTy9zb+rdXMGSyDCUJRGQlQ+QHt2NjaWRTJZ/X308CYMmpCK16U2eRN5zDi/lwe8Z587r0el4YK
i2BdsoOwWajBeApoh5DUgEfudoGExqpJ9cV/bYjQ8K/swHhGvKG/XikJizXffacEP/vTsX1lCC0D
vwI9s2V/pBCL4zKr2Tobn/UebAD1zNJJ0os4r2l81Y5hqn5lrjW1JhDaQIQKb7abt6jw64WplLR+
fVzrzZJ9vQ289A9CKYMtyI1NndbsTwtChVrMUMxfFh8GDM5+8K+AkR73lCF9RZ+gvlOSIfFmWxdZ
f7AKTaEqPKcu+nqoHxi94lvqQVx0c41k6nEQ+Sbhx/21LGtgQu5PTAHoYfirdXNKVzHJZJliJsn+
E9Me8K9hhmuhcaqp+HoLvkwTi9/XEFiH+6DBAjIzJM6ByO4wmMCST+zpvox0bmYXJZbpH/5Rr5HW
cSRSV8olHupHDN+O2mdY9ztbCNc6tP9t6kdNGbo7XRS/HswPfHXcEWtrp6qjXNhEkh9tSlGCWi2l
VqXV6WW0s2Q8TU5K64qNsgJPGQr1hDFFyzDftItyUDGQ3xdcVvUCaRWj8udXvYDq+nfnLfyNe7sm
QweGUyo8AcVdnKwj07opUn1n7DAv9bQuFRAHzEiAadc3BjlJpflP8heyLIXTkiqEUEmKTC9dAg6C
0rXEvspzBWpGMQZlB5ME2cNJ6T04Mr6boFARsG+1R73RiFHfo2iElY89k/k0s8Vz5e6k4Kf5SvsC
VimJ4IbEaI5En6w7BObi4rTXS6of98iyE+Tm6Jhc86V3OZO4vWTCk4fXopDRsXNJY3oGY0b7QiUI
l1Ta/TSvkfnHYqx4bZLIvnLgcQ67tgvGqYlDohtmTpptVsgEUlAZAPYZ/RZ8QpoAyQ6gPexwfPAZ
FDpPoGvRGNsJYRbMeDvgPYvnUrhbbqtK8TnS45wqL/eUd0I4idWh4hmaOvK3pI3JOAlxIbLC+4lI
1DSv9jq23FzvsSuXjapVVdL/EXd6Drxh8qD5YZg6LZBUIJjrERw8XruDN7q2NOQYibKXxejgPor2
vg2wPengbjY/t15OMul9Wo/jd/3DfaiLWucWjwLdwm3hiX+5aFD8oVCLWJ6AgwbqFR26RnfpJxsP
KWNTOtRjhuwDIdNNBn6gMReroha7qSRrDkdDsneSg+SyfzTz/9s8kh8NLM1NS6j9Rm7PepF5+xlf
23SH30Qvbha9QlelFAM4s0InVlt64iuKwcOpSPmyC2nVTKUZaI3udPXZEeYBAOqeH/sBrCey17yb
pwsoAH17n+gZdWmcdwVzCjtBvyQCOF7eUbyH9I1by8iQV8vtP7acQf7GoXeBQAIVk+zbjN/0HN6r
XXwJq54t4EVK10ulXfR79THuk0br5B47NYcY9xT44McT2u1Cj1QsOvxC9ivQ/GdZaqdkwOzSUTUM
h7p/XPmtGChI5tmF4+COaX8kN2DYsN8oys2HWGfKNU8DoiJymBm+PzAK0OvyWicDv9Vqg7Lryro6
DEvaMEXFtXiG0IJF/rqJjfYh7J6tW5cmOa94qi+a64eeR78lcgRmKuqIK2ikEFMA79if+BECWaYv
fxLEpUVJqtDX15kbnuYC+hLodvL3mf4n2zorFONQ7qAzQzAF+K+xedu/WPiqkvg8xvitAvZuJqvW
lrvmKx+DORziCz+kKgxsRfqsnyy1pTWysQKDcNPWP5fREy4lHieKWD76SvXx8AQmwVlNCgaAFPnN
AJEYN8cPQI9pF1oSotBotrU7Fh19v563Bdf3nlsItrePsHgxruWZghhn7HcNO1qQoCUOSk/LckNK
HJiq6mDmxlCRskzN5y2nfqqynUdsi4aJm/tRUvNG7hIvQPJjYWgLag7A48VZoSHUNMBFIxH1QvlI
E0d0zt0g0ZpWUeEDsHjvle2BepjFpEtBPlhlhQo9yCEyk2xp1GHltjmJa/1X0rL1WU/nJrccOBbT
ixniT/LRBdlSsr55RiNYYtmi7NL2lSe+Coo0UzVqWhIc9UzdmIca3k60yTWg8pijkTO/0JxvnEfO
4zceVaH/iMtSbv5B7yVhxlIy3RqE3ZHX0rwXzRP4583uN/99oyrnmROCcufLjI0muf1qKtlM+iKS
WuXsZ1RZkyKzPzjj2vmb4OesIxmK7y2kQA6P3fv6cMbhrS+nYqhDhJ7bOIIvzvBUQskxLxf169/+
2t5VPy+rrUS4KEluWHMtk1QDy6CRCxAbcsOxaRI90B8pTrJ2pXHoHLXkmmligHQzygSrIYiGQEJn
6+gowqfK+BnRkxUZKBgFPTFhc68Op2po75BZYkhcg6e+bDhOWsYqYuMpha1IBYh1K4XRSLpZFgO7
9h3yvlfURrRycSJei6tA2Saw2546LcuV4HZ6IHnt88F011XmLKMjrBuzQtVv6k40ObtGipLWC3t/
fGYRFdK2nhMDuGRF5z6oeOaf/Pdj5h9sdLdE6QX+NKrmC5Cw6ZcBn3evmJXEbhsT5DNUG5/EzvL5
/LJBEz63Hfpmuy/Kur7BYMpDSR5sVrR1plDuwNZdUmtQHE5+IXjns4hN057eVPcha76BxeE2n3kX
oVOGZTBqS+8BmSaOP5AwFAC15PVGnnpJKRZovGWMvpfRt+6s+NX0hYMD/clZ5b0X2rsKf0MQHdE7
ljs8dFHwYsnkh5G7z81c1GIx0VHHoWhY563WAlEyupnsb9mYDMtKDUZn20Q7anyPhoDRa3M8W95s
yGakmxBvD/RPIJEaj4YrJ/9bk/AvyCedWjcrN/lNUOSbnItybWF+4lVkYKMBRoTpmd0fKTv46XIj
eJGjFoXhJ34AKYZk3QgmzEK4YIyLYGTUAnSAO16Fb1CXKjPDpN7KVVVxrpkxfm9VBxaF5fxeMebc
JHFUO7sxqFE2eqn3+J29NHB26FGNSYxsmjB/vsQKF9IUACtQEgULRVJ2HTvub4JN/xCO54gKGVPy
3gzEK36PbSGM6mFXvhkR4AsgD4erDI7aTZwj9gpce7WilnSyQBsnvEOWBR5NOpz1KDHvta3JWni6
lx6VX/CE1oCgc3QjEVEWo8FGi6f5VGmR7ZoeUImGEM5AUfYyiskxCAqzX27J57JQWAYpdIHmAq5L
i0h/a8Enn9b1xtPnALIZ5r82dX6w6DWmIrByJP3RUOgxxD6DPMEb7ZuK6V6dfSpxhhqb4eRn1vJQ
2ER5OxjqskvqgUDcla2vqTNzS0vFfvXW/oX6qOJpoairAk3neF54cVCckqgHLbaWMwzs1hH72ZG+
noTOGXvYfV9WxRz9eIeaCtzuj7o2ldsifYGJ8KZCdMXsHxT8Ub8B6KAORVetBxccLKAFjK//D0me
BtDAYpudeztTqzAkIntXSH33pQNTlL5x5LqvrrxwKemHoWYqJ7kxoAmOF1PE5nk5G4lTkpMjrs4D
vCAQX1VMjmDXkYQ+JVjsetgxk2Ai+CMk322/OMVEe+Fhci6+OOZNM0UOqiFK8w1lDvK/MYhUfyYq
WWJaM3MJVvYMJ3FrfzKMR4dzajoDpbisc8jCJPnz9fqi/NuPdIMHiziWa5e34/6N+gauc2z7t1PG
6ZkwVEpzsU0Z5tFzAWsQPlVwntnHvWSoVix8PyMzdPDrdPWIgKX6nhCotwZJC5+8IsFnaaolvaTJ
UFz/aX1mAEr9A93JL3E0x3q456CJ1jHlu5PuhbL4f+yPkD+xusyhjumW1tBuBRu1Vu02+8BvUJZH
BqFGZDoLFRaKa9eom5Z109QCIXMN6eyqYGiCBVsvcTkV8mlr3foba68SZWKMiQKFw+MlFu3rpqfZ
5422jeqgkUPJHDdmqPfPsHM2DfBskAypS92UC6PaR73yem2mjXxKfEDtmF4VkAkx0FSKZ9vrUcS/
Vp+SyelFGWkyRAMxsBgiRXm64acgpknwnrt75gZqrgE+VkYjXxSLBveEQYDzDUXgxlITt3OP2qaM
XAnSth1CDiokbQEwR+GdhLeWId0iyQbhAqKVUSYl1jBT0k3e4mJSUX5IkriV5TVs2kmNsxjqJUSC
qJ8SODAqBeXBJ+nnCu2YnF32ATrd7rndHrl596N9TMQzCdUV5Ov4ytTMin/LTltqhFFNA8j+cGgQ
ZwzYr3Dz0VW4X+xRO7pOugdZGK34v80kB6h1Cdc0aWzP5lX02bY9IP/BL/jX6D6wRUaGoihwR3ly
E3SGd0ZzQ6vXAngZGs1CLOLnoXnZZkkl0AsRn7mGpyIa6NkU04hFRm5BOiU/otgBmD+yQvy+visf
jw2YgKUbZ6IVXx7aqkfZisv3YQC64oMQOlFwwP6NsNG8C2LY5q4bDq0T02aClv2jehqkR+yLCqXu
sYF4Dmjg0zXkDrknvob41fWQhC5XEOm5ecpS9H4YiBG58TBOUuv6cF0dR04g0JsroC2E1qpJ7mUx
yoQWu2xemVccR/QNO8+z9l0DqQbca7pw4pzvJSiARUUoeAUXUOG935xgJeFTNv/rU/jKTeq8N2la
S+FpaJg97qAaUFE8YUx4o8QDHQV3GvrtHqJ3obCW0/UVHElTX8IAhDQRptCW+tiuKvVBFda+rkp0
M2NPnTVBHih/Odoml8hLJWTZ5xN6gJIppfiA0/H8A6z7IXWsrdwc5KDAjfDOulcbmE6zSFn3zy/y
UvdnZ2YwA+ifJNa5Vj9IwRuiau3Ca7ikWRG6iKmzNOmeWGD0Yhyj4QX9wXV2mWmadxCGskrpoGnE
3Mx0hU93IMQ3/6A9kPRZMkE6L4MuWOw9R110NfFZMDGhQK9oARokJcTSfhi/pi/LG6gF/hV5nwuU
FC4AKUwUL0gLWCvFVsjCJOM/7agsHghWUYlgvQFGqum2vAEGUlduaPif1TQ1/mWz315tp1hkfXlc
mNTSbrSAEzLRkWKop2ITaIobIG9ZzXFDm8KEDh6WqOxClCBCpK0jP8N/tKjnl99/yuBGes8VW/Ws
nsN+IT6FhNNljAKYeK5+fDjerdNlzFanW1JlyIyhwk+D2WQ8+mYwjLH52NMJrWV3rQl0PXx4ZRKO
HY2t6oTVh32/Zpkf7qNsgs5TJmYrfK01Yi6euRR7UVKAYY1uNw1WFV8Qnq4W1CRDyKrJyZXNoT/w
577OyOCVgjMcpsySyYJQ+aU8LE0LHvxUs8hlfAvhg90y+R9uKMZJrXcb71wI7dij08xLBdos0aFM
n6f+NTPKyUEqer7p+MhJqZgYUz7rPJgrM1Ax7mbc4n97rnnGPQh2WBk+znqYJ4uDxQOv6ShRGDT5
yfJKQ9S9hLzYVjMipafVeY2jsG1hedxIgZkoJ3TuROo83Ml+1dvMcMiQi9qf5GP1XIYGLzGS9Fis
HnH5U81A3n/jJSAifYCFR2iAAecq/6f2c/PwGAyYnHuzoDQt5Qf2RByVLBiYPZiAsMCtICyYalrx
tlukvzRiolfKqbKsxMY+lDlI8o7sC1GU7jlnEN3nYav/wj/St/i0IbgvsDkM4CvVZP+VmlSlHUvC
uUrb74lfj1ICwBJeoLu9hv1Q3El/X/3WmPfE5R4aJxTsdM7aCMnIvjNjsJVKvp2wc0J6EpoRdByS
qehp8vjPrNyzXAE9zOR8RG9EO8CGtm8D4Sw5S9aCnSX3L/HF1QfBPAv62kcNW3W8o5f0mTRq8Jk1
fVQKKYut0oLXCH+Plr4b9z9xAmq8ipEmDkIh68EgQwVE/6ykFGLSqRt0KQoPwALKqOmEOZufp9hl
ac3YUi6K6NcehLfOUaCvdGFUkx1xax7nZsn/A2aXS2sFQadYPBZlatFVSU0ZUW6KDgNPvizBSPUj
+0RYYEu4IEHIM6Naj8a6ZOSNEPfepROdYtQ7XZwh0aqmWBKnuqARSW7qeVz0eeOxYwXZbbIaUD35
HwSN98y6W3G0+cpsh/25+XNKfDUKR6ioIL8Oxk2818YrqR2BRqErYX3wN2woEBEpXmTNpduUlVBi
+ptsjfOMZiu38oDde4TlOTANTEGIv7k2J/dNDEHdxdBaZ+dHoGsdtJ1j3VlTGiUbsuJRMZGMUFgS
f857hDQYF7erxPJcyfUKFR2E4JyjeHfTrjQhz9OdB5u1Kl7LThrSE5pzcoF5Ovp+unrmseVX/cAA
tK1IDWUIk3vYNCbXkoNdC22LoacNNGYHjEBurQohNPl9Wiltr6qYYXLPbwaqsZyE4yVoF/H4YeWq
scAXyGUGfCvfdV8e10z1aVIzW6RTQuyFPQnjpo3EB2YxkLzkfLN4WlinPgfCABUvZQw39zd6mVAN
31N94sN1T/9Qumr41+puvt1dxCb/JwdUDziRIev3nHQtxnx3NzeJY5wvOasRm2mOTk8nWSHXTmWh
mT7iAXXFuK3S74jXraIVKtTh7eupLDdNMA+ChPsAKxtf//MkZm2/2BkWLdECrODvGWIfmWKadbuj
68Fd6m/lWtDUPmQtdRS3FiYN12CmIy4fTDorYSX5pG2lBUAUOeRbfXPg62K6hS1TNr83mUvgd1mR
mooh1ZGE0njd+jgW1whcvIMKD8hNryxeiDaYm0EmjVEIKVneQLfXw76DWkwd/T4DNInMOilP0t2p
vFDlCb4HqjkHa+5nT/QL5hyhlILiREAFKj4WX2BcyZlwOFMXlvYWcFrYGHmHKsOAcHxwIUeSxX6a
hYCI4VPmn2Z8VhvEwlMwgKWSMz1Fs4m6jpmlHQHZ8ZtHgeKet4uAl2Xbosn97tnkFor6OwAtzIcV
Oq+AkVhesJLKhvvYWDGqH15KJEiJZ+7DcgrD6QfOdKyM5GXD//IQ78D1TwLIgEbUI31nmXnKlaof
CsCIxp7xeX4lLrccfLnSnz795Z2FUnRzGusZqDYzp+oDc0qW4Q3CiDbrEUEKx6lcA0EYO+3wa2Lp
1o1qHRRg5DLXfrDT+mTjujNV4o5F9HB4AnlTH5zw57j0u6tA178bpU4nd6HjBXgChrAAj6+PtUeQ
/vHG5OCTI3s8hSnyhgVTvmTx8eqgNJYiOZGkD/Enowl8DMJfjkEfQ53u9Mm52zsygnX+yXV2SWrH
3PVknvJH39n7m35g/TjntaPhqYB6jpoeIKmCgBj48KU2F+7LANGsbCM8DzuACZcX5dKxwLY7fjoR
KRK9uExfqDqI0EpHQSu2qC3FcutSIosBttXGsXnf+9+nl+D/6SL5uTsuFX+wXOkzATuSEpX5aW9n
1BQ4NlQMaYb+KchFn/4Y0y5n1im0TQ5ajc9u3KxN4AJck6zjOdYZKcvxCc9Fb7EYqqNbhIoAOtu/
3EdBtVmWYbJlQD/JfVAlJlFk17Fxo5sOz6CXWocIlinRY07WNVKuRyBPz7HOnZDnBPYDex93Gh0y
3cexQ32fpksFR2hYuanWZenpHlM93U/i0aktMlz4GK4g4lGvRDnvvfrspA0xx9jk8qKPFMSDhhS5
DuWxBR1vKxO+hJz6buSYs9OeogxXZl0ZmNbcqkIVxNmHOerwMc5QCQf7PRD3CJBED/Jy2onmTj85
vBhD+jL4gdR+BJxH6+vnUCsvPPGcS5L81wxbK1UWl4hJUvExsvL14OlHJgbI+6+JuPaYrGd//Lil
NWWs38X6bi4oxLgvtG9JYq6xGVAfzBcxVJ1Urk7fNWVK443N2koC+Dg1bO80v/NTFTkg7d5efkez
tZF7UJinqcqs/5zLWm+4cvlPBU4PWRUwZlRPLzWIbyXjC2S9gEDehG2EFAzyy78nP5ohNZkOBHZo
XWnEFZiWqSZ9g32OWtdbkuVwRcQg3D0Di/dk6FSCubgXWayiRlaefQu9lUZs7EFkYqCvqUiw+t6q
mf/Bu0+JtGQqPyBF+vcMxYxFPfiO509Nal3MaTnzJS8ekV7myYn8O2VXnRuTLjIR7D0kxmSOI5iX
Fo/6b429GzqYzOwkWbDVjljXExL5paSoAenCv7/Od0Qdp0Xkt/3KoO+uwy9hecq7mtsjUq9NNtin
wf2ce+CCaP+guBUOdnvJxZ6CKYnZJucW4NhLV47bzm2Eva+jCSh0ZpZkEe/w9Z6pyOI2WqJqzoGH
YYbUHLXm/kNyzTIZ+QCVPl7EPqbND++j9P05ozp4QLi6JWPFNhJUdfAFoSPFxV+j/+uJ46vBpUNk
iTBUO+102oFrYbMXGHaPynusdK/WSqcpPwEmO3yIomALOp7MRthz3pyGO6mVms7xaVh5SVb6Y8OB
FJj+0qwxGTFxFuhIJGnylp63bpcmZ098stlXCVCXmZju1KXrJtQeY4yWzhGZC+KFjnWhJdN09HaN
GhL7p7Lyljt8KyWAWCBChWDEFLOR3tTwRLfRfiO/r8sQ/100JDIpCdSB5KSR4/2qr1BcLpEvGdkf
kkNgunZ9qCTuMnbgIZ+L/fOdtKbd7r8zlQ0e6g4rHXt6I8TwSQJ1AY8j4sWoTnP75Vgynj2s7Raa
Fkivb6DHgf3D7xsu4DT+kvtIm1a6SAv8+LoRRl3OXtmXnVSxUOo93a8ZqGCK0Hzs8Ih8q7OYDreb
7ZmRV9YrmQgbh/vCNyFcGqsmECjHSCplJnSPrWxrv4yuS+W4lzyk1o0gvoltu/TCiksg7NNjMQdp
OjMfpcy6Y6bybGSwqDHaNbNofJFHAhtGxpmsL4wcpBCjA9UHUHfoZxrgdQN6j5XbkmwziSHtwe4D
c2wbnBxu2rBWwawURYKQjgN1uaknTdaurQykqOB1ze/nZwJIVk9d/zfsY944aRaC54L67xYgwf19
YVgiozIc+jA31r9MT/fcpu8NENmvKC6nL/bjYravehOwovrLLfRuChcfWn2ulTXmDpHwM+ODoalN
2BN9FPP9ls+fd8tjiHxhuxE4uxXKNCm3sZMtOMj6WnXs4v8JvFYNDfFLaFPHgcurFcYym59WY5r4
9wyz5liupKXEz9TTk7Wz/aombuA8+qAD40yYl6itJ80bIm2/8nRMtefDqLVByXT14Lxpm8H4K7gK
oJ239Vy39KLs9XdF0ILDt9YefIPYJuVwxFyCBkFPlaEuX/nU3X7DQ8aWVVvVqWlS056sS+BHlQ1r
kJ8OK7vbYplRFC/WRxEMKZUxE9+pcLJsCuaHwU98ANlRSFwf7Xfi6sr3SQLRTyrrJgBPoIOWE2MP
eNIBaLawQrQ4saKwstVfMZTVA5Ov7ItslC4ITT04SiAIEGZz4H2HAcDp7BT3hBxC1f3d39lSANQs
5TyNWVv71EKfNWOphIuNfom7fSJeOQZnApfTQ86OEFrFsN+Zh3Cv1vxNYitN3XK5vbzPNOW/0MP0
CssQOpUmNjAbYBG6+CCkO+q//rUS2IMy3qKGWqJHpRfR6TxFnLpjcntwRE3ahBGQe4k+/eRXQqGM
zNeZ+bUkv15iuIWOGBQS83E0qNNhx1xuBAb1VqhBDURu/LV88o3INV33uaWDWoQ4FrY3sHEFW/Nd
LGawq5TvwC+3QQaYwqPcrLZeGr4WBPKEgVarmSmS8/0xsirUOJnTNUxKIaagFCcTqmb0IQkO4gdb
OuCit3MuToMBUia3AT/ZuYH7VHRTBeSfKy6xpwdrZc5DUD3v29uoukZ6e7UXjzT50h9Tu/mN6PNH
6Fs3cVfVerEJVtrm8ZlXqwbBFR03UmQdyQK9MakQzOgTQ0MRdy6cJFAtrvtpdxYSfS9W93EaaWr4
jizoGbLwYDOVn7EMBc0pjDYEKoC1eDHd0s/JeOTknB35YSpb/F6zLpG1pZHdLKyXAi3TcPyTYCXI
tYJgYsk6mrI6wOGU+Ze413vuwjakHsjPS3mEcOCJdeiLI9uMSPQ85KK+1kFcLvrkM9yG7Z9Xk4A0
4v3/5fustEquD1Q6PnDAYvqT53A6Mb1Ugn+3/WGGmLFX5cOXAgMnOq082XkxmyONgSEHGoOb/IHB
VY88KPBISLqO3mQKAl7CdpqIpyffIUBOVQVUusFx9idcL123OhIS+jrpyNVQO1hXSf47B4xVSC4g
4k1Yta7X36E/dlEd7WQyfaKPDu/eEBag9gYNi98GNTIGOiBFsovouoLFmz8XYSV4/7HWZk281Nva
QkprbaKM6KTL7Bs2RVjMggRcBWuBeEvOXo1bYPfpB90ULkFBqw3Wz6yYRWIJYUb8fyGmZcuWXJc2
v59VvxNGsOA8bhRfMf4qYyb8TWfYIR9ZkOGFKMZZhwtbXZ4wITKTEw7+hZ+VMghgMtAdR95D+4l2
kO4rg8Nfv89xNMp9QTVEReG/uEE9lWJ0rVRO+xKKiERRFAEdsKxfiRVGbJMSZWS98VxdM7C4102p
uE/Z2tvH0fSaUUUM0QfFHI0404ATIf9nHMcYnrq67w9gbpg8SxXUnQKZ5f4/wlGAiJF3YnKgdqlk
eLgjNncg9cbZd+6GeB1PGjnUPt3jmkXPN2XAl6t8Wrw4+TE9rF5i1qF4oWQMnhFPFI8tYQuCzduB
Fwz2VVIHn7tTJcZfCe0810ipgw38JDH5DyrtNrWnUHKhKhMlimFEG8p5yNOaDfK/VpSL+ZYR3tUP
7i1T4jWufHQL4z51wVBiGa+okzLJYbT5jGji3TpDdt/spuMsFwKForNGC2nk0nggmcIpT8LS63NX
SkssVq9L8cW3lsS/9cir8JelpEFpH1BWYY3j+Kan7sGICBJuBjsqX/xaOzBWBVaeYZ0ISabYAvVT
qOJdR4Uv86c3AcjWspnCxFopS3Yggsbv+ipctIkAHmoU6Tgp00JyhXNmu+E7vrAeSpm2kdURZNej
hR9yWbryZBnpQmkUP+8JqGRu0E9lnsHs4sgr7cHJ30rMtcVz/66I+6iuN1bi4zBwyqMK8U4j6YXU
CMUFGrs4pxXIHJ56MObSxpfFkNPfMQ9Ng/tyxZK0Jp46YzsxW5nRjkxvoCb4kuB7PAk6szYNgh7R
H0FR+tgOzTkssjV65FvG3AnPtMjxY40N+dVBVYiPUhDpelVVv2f3JxDgZzBgeM1hv31Tm/+TYhS+
0rq5mPKvf/mJATLw3ynMN4bgQiKdXmBq6/un4ZF7HHdu6h9zcX7VDYWMPuBYDLBcNnIuYbDc9Rph
/Gf/6/p5zgnnMyi+lYA46XEs0szggbVDttzTIQsn9zI0bYxz4psvzu2dMx8t5L+Kc7LQrE6GnCaw
agwgWDY/xwCqaH/L9GmMFqxt9EQ7l3TGAcygYnL02xsZJCwaa1Ql30YRv+ZJus2uPYSUfsfz47kY
6JNd6U4VJ71wTBjZNnCV+q/1SpvmWERhCkf/eO0vlQtuwmu58jvVziFJkpTmgV6B8RFc0e2msx4J
o6dajlBVLI1AI/WbbpAvMCGh1Ef2CkvfycaE06ExNP9jT0aCJMYOgdn7QpuPXeTE0A7fE/6V2bjk
3UHLxhGwQZqounq+Kjtkwn4Lqul+fuPpNcQUR5vhgeebAzAsvgtTh2d5E6m3CgjggaIL8suaEwFw
UKGRo/abFjBwqoTNJee30UMzTSwMuZ4bvKJWCGSvJxINkqH9ve3qollzislTw0QGRMMIM62EXThO
Iy6QpfOz8R8q5A1Lzv/rqhTHkV5xl5J/IgrKgZMuYlD7DvxA7SKKLRx0A30XfkrsPwg6HcxmHyGu
ne6f+bEkU65EKxBoGvhDSJsIiy+QCO3oBqKbw1J34losRCQ9MKCGoiapA/V+VaPGUGtJknMgljDR
3bsvVE6s6II99l4/0LmHoeIllKqs0XMXn9WDGc6oifSvNU5nQHiccimz9ldJ1zRYFMnpoev+huf6
a/G3/h1K0p/ugnl+OqwDAXznG9QnD0yiT8CPhqPmoq4sAIIi9Y3880OHI8GXVc75vo4f3FV5ZiJS
z/YO+rqSwNAQQUl5xm9i6CdTVUm2pg5VNy78VufP4gt6pMx4w67Z5Oi9B5qwG4+HJUhJZzdm06GL
nqMsz+m8yXKhk8cIh3JsB+RvMNxVjS0dEACMNMscLVcRnztVJ5aYZDXzVaj4mPUgRfSUMlayX5Rg
wWroUdAt5I65TYy6GzN6bSAg9mOpGxpJE9piYDEIEImRuAQET2suKTDjn10/kX7r8Bw9yUlbLYG7
M485MFnW1ZKQ8b/1fGiBch6m8E0x8/Jt/P532snBw7TpbQ1wSR86nCDefDWk38v2g1CmZAqsYDys
y0lbsJYxvZYTzOBGB8I7uOhPzWhvV7V0PsSWoiMljxqziqurIVAnmKWOuNypAOh4H9OPS2WWhMEh
JaVkSGagK0kg6T2v78eAoWeRmul395rHKmSfnU33c3BkaD8X0xueKRrhKRfyiiQ43eZVlS7VQFt8
skVzLkvUqUmiLXdbOdlQovRxg+DEhHlziMjtOUBWWWttbx+uxPF44I4Ti7PIuAAfNdf5v6PsBK4V
q/GWl27pIlMF3KyLIIfoYqcgd/Hv54qnTgBNy144Wi81thlMdPJ2Tgz+ZWxlx32VcWyFGt1T2F93
zF1QHYpZXD3oQfZc5uxWrWmoEyRXUMAzrGnNs3/lzuREK90s7DAnfPKe82yoO3nh+aFt/rWyaslE
NM3BuwhZlIp0x1zSUnkv8W2Mw0eMfvUSBrpH1Fmu0UNO80taIEh/+qtNlFYYOjmrqjkpghgV6qoo
ZaSWhfIOdPybKHYMBIql3/PzuJzoZxP/DpNVflTJkABPy4OxiEOBf7Q3FK0dDcQWtTGonh+pV+I7
60AkXV8cMhI8JXTaHhPYb0ym+Fpihxd5WLjP3awTCVnGKOP7Myeion1/nR3my8oO8z/wJnCQ8fLh
IMRo8sGKtft2FthFTk7o1kP1GAPq+W5b7yNAvvbgaBmzhdQkWFpE9wq/Nept2co55tT2TW9zOdAn
NZ6yjth3ez6i4oi0G1yC9qEAFMTfeOgrwM9binsBwrO1rEHD6xgXthL4I6n1bFZRknHH41z+4KOm
9w8YiXMN650k9Usc1ePPpIbhUVax+56mwdViPUl9k1du3s+QZIgHi/s8cKNwdJ+pfmjtsYqTg4Rt
V+P92ftMJXkxRv3xb8uJOfMGvxO4K3osA1WPF1h6a6AchfmW7GJNYxqsM1dYiETCkQk0vwarZ/KF
vjeQgD7RfD2ukkSnglPHCiuc27/OkvtSIq+3h7+izIe3cV4EzNlXKDymciW7k4iGL9HWg4Ig3N7X
dzJO7AfnWdWv8W9i6EyrdxyDfOJmzS5BsPvGhzZpfhLNnch4W6upB+lJkkw9i5tCmUAAi5gNyY0E
FugXyuM34XGdbr9kLpPlMANcCyq9473llJ/73d5W2XodktEzOn5lmDIap2RpxSnrGPDUWpDbbAu3
jEnnS4ONdzE0AN+sPGksf9QoswT0bPfZ+XHs1BC2jHkWzCPU7i3LdMOlrb9IUpt9DnO/ETEMGeOr
RD6jmN5vN8Gr6/WjuapGMNY43l9CUlZkZ0eKRlu9l+NiCLzOJFHXUOthIQzTcbDNg7PLX+OegaR3
zkTIj39K189GhB5IM2qnQE5mPvnKPK+Fk/bMgPhE/4xP7WsKr8qaO4Wdc8qKrQ0P2N4tyBV0bbBY
/TesNnYkhJaVoV0VRr4zCCLuYu+v9HvOVcV3IG05y2AWQmcwQv+nZbtEDtz3IZOIq/8xni5epzsZ
DQBQ3w74b7XlZQhe0S4BbqDQ5f5Evq1sJItPNJBL8T4NSS/N81ODyEd6m9yNKPlBgjgenafduB9z
J/DzoR2BGo9yUkxLFIiPgt55hlrs0Bc+2kXnd2VhKXVRlLEhkrmXEuz7M0vq5JwR5EsqTbLC3FKW
NAK1PHn9gVn6w1NyqNRUUC5gYBnTB8ChwDoWVi2h5EdvYKhTfKBuZ+IDL04Ev6wd8nN0WfDzbmZo
Aq2BkqLrIavtF4ohpZYU9gIyRknIwvzzwnU/RbtkNKPWNSRiWFSTlBLphenoXlYMxMjQv+WSJvlY
u5lJwZJCktDw9lt9ONxwbquJTCapIRffV4uInVVxeMWe+nsIXmcV14nq4qCp7gSNF++AMygKLd1x
beRXnGAT6kLveuOfctcs6eTQEqc0K6bZERSZzC3ZeuLY8yAm9p56GWNgWW4VZM6iSyxtWknqQyn5
TMGAwJWDftxOb2FdG8xOGAVNGOFn7CcOrFhE8yjTDnSWBXIimznk7Ml5CaV+QXL74ZHq2bJSBQpT
FKbTAguzQCv3n80S7Udb5Hznuk2jEpsxuJtI9AJMpxuh23hVFUlBZMEEf27+KBDK76qEA3LH/DwI
QT+VCy4rvRMvdVpnVW9RtstHAiCQhSSB2jsSAk2KiE0kq+KFIn3S80sdrdShTxYDpCi8+/yu8n1L
yJnu9NO8ajaVDXs2GklPfAtOnu2I9574VxbYqTWMQs5JNHE1G6ymvCAjevjwvc3UIGsRmfu+QlE9
n4Stk37HuYPhVaJ9xLkmkHkEZMMgDTBs9LNaqHeafC/KSbqiuM0F+U9Jo+zk949qlTkIMvGprK4d
8/vyNUxfE75j1z56/918Q+7hC7H/hTbmuBrS45vWoCKGsKgpJvd54CmPTq10plPpxVPAOwS26GFn
GsiZT7ab8H3EGmu8VLdtyKJfUNug1WUrGV4OBSLnU8zLvX06dHVYFFCZS7qUMNuYl3niWVURLvEA
fNkVyYUAYrWp2NmY1ocFahwWBxann/IrsCnk8pQMq7kvRkmmCxHjw9ba2BvFG4AUr/22C9GVSoIZ
M/6UuhQImmobGBEJOKI3zxgAml8761CpoN5cNFl4ENbLvFlfOQYBM/4WeaMOuGQNrzidHB2Pv5tQ
/WRKr/XYvaPVhfFNe6QG4xS5cVmPnEEzY2EWAhyX9wQzz3FPzy+/k9gYM4VspA6rZUEoTdvtixzM
TF1FgoobTTE9Jc47GT8UJwJSyaWla61w8yzyMbtBVrVRKvM7fL61khGdbQ5Vo2gWHzxNPQIV+oPN
gLR3MJAyc+FmJy3w6ZP0P+7naAfORb+bU7fzDE3pSlWydOlty0Yb+3gJ9VXz2oKBv+BP3xUP+4Tl
UDNIOOt6aaIVYebGsD+U5vRZXIMcbQJMyoPP9UVOPK4EcArhLiO7cUkYy8dkmxhnC9G8KPCKMDyY
lw2PqHGqYbOqmgiAAn9PIL3LZz4zqZoDI+Mupe+Zig+V2Rs7d3QbyOBtbehdNgU6bmhROXw9HGbs
K5EypoZ4zRGDF2fSsjeN3teraOrsijPgvAoQjaX9nOOxpDQK9XGokosQirXIux5QypdhJKCPMNAj
TQJtphTjY6fu0y//kXnau212bDGipfqReuks2UZ/5rFD+dr2HT6+pCyzh32edAjAABfdVSSQw1tV
o9kQ25Wo5IGjFbp/RhkKMmXkenV7tsbyNvaNfg+y2KFlf90DfH6eTybde2Lg5OXLS7aM0ShxZ2Rm
6IIUQM/29wEcBkSMweVjZdJETfA39s8rWC00qBIxglRRcrzNs1Ur2MkXS4IhoKRfW5kFoiL41Ifx
E8PGxRMEBGAfx26HMFm17CZZGYprLI9W1TU6sdqLfgK2F4IzLfuFF/92sHY7BqhCD91Evujs+T99
BOYHN5RqNRhq9prKCMBvzwRMZF5EDsFgs1hRGzVy3+t4zsEoZa24nOc8GoWB7vfmxaIhFLN4lOdc
gdGepF5pazVlYEVzPiFXvHgsTbDMRp54l0PeTMb3zN5XAmy1pq7N0FzwUDWDbbd/myHpfgtV99kp
q/PPfqausWss3x2wiCsy3pJw7UQg8ye8TjgcmXR2Y1k0nSNGY15AhYgQ4brIE+EqWwQkW6DNpluP
upQXWZ3laXEIQOoF1MSzFN1R3/OrIU656c6zSOmiBVyf3wXG0OzkH0BGMRcEhrAMqJ3uApneO5iB
c5c3XnUXumI93Hk54F6w+DVzYk1KrmUgNMFVO+0SEBxQn4ZV5S8OXSGMcKcDFbo1JwsQhwtoGSEZ
xSG+rHQcMYbpvOsbKM9BNeHbILJ7g0L09PMM8ZtGhylMtQlD/UkBKRU+j9g2izpoy2DXzjQ5HFZ6
OhgqFOa9vyD07KdjxESPP8k9R4yYoRVfgL+BUBw/1NJS41YA33NthCyHGUiWijyT+vqzRlU/ck/k
VfLQqsHH4EjQEIJkPt03/7ip8kyu/K3PNuSprHm9fP7lm9MPDEKbY4Xjs2Et4wbN3KFb8qrGgZaB
SsPrQPylejtGtadJ1jTw8tWjcOez1fAf80CrstMqpzG8/WeTrQZEFzGqtUifD0rXNucp3b/4ctBL
Pjt6fX+l//QbOJqCbxakZpL3IQy11BxnHL7sVj+ffQh/n+Me0zpoMfx9TXXI463LQC8VcQ8eilJC
DE8pY9qNbA/v76hKfmzPJVVFg7iv4C0xeFYvKsOu1uOHPhT9EMxaSVIwbShZDFtccFRTOrjiFiI/
YA52FsjvgdlNH/qzh9zNwvQcyRdc9x57IuaYFHhXolkMKTiZkm8Oi2YGkkCSUbtw+wTTj79qH9aU
aS9XKo1c4FDjfc2bGvE1meQARHlzNO2cD6P6dJpO0Z0USD43oNHJPZjdU9XDbcZDzIRB3dToyQRL
YZjUWiNPsPzt41i6+gyRr1dcoq0au/s5KnyrLF7GqYJTxqBlQsP9CwbzzVQbdkguYtHrI5bKCoDo
EaLkZ3rfufUpmR+1bSYsJ3yblPTwZjl6FlGEzOnGVu2btVRWuCPo3b0aPDw1kMSn/jPKgL82PcVq
sbk8Wz4yzd2f2FdvYaopf6nVxsN2/IEZDO1wYSvqsrut7PvJxZVnDBd6f/qqBpHE7+UH9P/vGrHu
/NyM2CfBAbl0UbzPE/q8B6wezD6tLvfUpJoV0Rc7BWwc6EG9xmNW63KBjw7y9oLgI5ByiXWEtqE0
bEBnqvEltJphXok3i6EJWtoFxknhA2e993X0wLzHCYVTbaLDMwENj6R8pdDIX35pb1ORQoS8QOXM
9KqQIwUY2xiK3i4J0RcA3c4+1USel4Z1FAyEqIwwPvzHhOsGsa8M0HXRfChOcFvdfYJaQvrF6LGe
WVcjBQiETRCb+FAOg+41NttBND1tyucgflfScb+cEHp81MYOepXlINudxYGTRf0g8ow4zcufFmh+
fP018c4As+zvDqKDyPytwSxJsPPvaVumQ4A0EBMcb0LwBBY0aF4E4WW3wVDpJ6uzkhpKSOl0yc9p
mfHZVm7Y/LIszUKtGzrTw4KdOrgkWD5Aep6ltlknpqQ/20LLJJIuV4LBgEIIW/wuGvLJz9iZClJj
8Yl8COEQstEMSozkRalTOct7qy9V9v+qPEwa57R0hoRJZObgnArllY4MhDGtZB6ENiDkFWwuP6Oe
hzC9FnkNgT3SlaSNNjd1SaePJ9vTFkmMnZ/OeuUIW4LItBFpadJ6DL9VOQH/527EDfynLNrmMiyY
RCvZzdmq2u5MmdAjl3WRi3LqOGqqZ8OVQJScbM+3CkOQA7x+yl33QEebVzos0Ur92A0eidGnExUp
T42nQVAzTf+HD1Z2J/6zlL196N0NEFldgl11PJmkGaeuIH+XT3US9xav40/w12lOkY0aJmKxsvcK
aKnA5tks9RB0FfkCcMtMKZEa2IF0IDBTEMgThW3hFgu6aiyFQ1coWfwpBmte4BOvdzeb7b6g8/eP
iBLGMm/reYLc9aVq6AbK3tEiCiQxc6dTDlPvY4ULSonQbRTytfdKfDf+apYoTRsLFdfvVlz/DNP1
i8Q82h33eA+BaIYjkaKoBxHgemyxzMN+RzO3VoqdCToB9IbMriQviJ5KTqIR7oX2qi91rim+wV0H
2xPq07N05w8QIX32bgrPyBLQFElVIpTy4q9YlfwGCjTeSzPKnNajbWQzU0oT+TSda8WPOh2Nz3kv
lfkmJ0ll9Kn/xe7+/z2jKtOAM0899tKJGatNmVqP4xrTppLODoDuBYHeqsYuIpI1m0RDSXTpHIId
At7OW263YWldlYdLf8K1cqEI7zIxwpcuyJhI4zG8yFbZCbAPkxhFCf/VWQtkIOoEPBYO34ST2S5l
/zdkes+ybY1LLr3NC+Ppuxzf60R1aY4BScoCzk5dR6uYMj3EIEXwdv3uj3QT2EHrWLZEzrcsnIax
oDT9bySQUAkinyyaScCGVnimnqEsRPsIWaH5s8aQLR+1bMdjGabxR9deE66x261FXsGGT/BEdyvg
vgH4cEO/GZ4O2g5zLusd1m0yt8Ns5w5kVK0Rd0cPGD9h5TsqzrM4+8yxPG3IB7Ti/+7kDSeeteyW
x63Dszekq5oJJyYTARJkH9E/3bfpsC3RLAHmrz5T/K966rX1EoeQItHlfswuAbmGssbq3ZubQTLf
DAslHk714+bNLXVQGxCrjmkLuk8tlpomRCfzGXa92SmXR8DX1aKqJHPU57/UM7ZRb9QaXrSkBszy
GwSn8SlmkZMvBRGStGZXbNVLwoy9Ls9ZkOhPV9Wi8uicPy4HRaoQ54T/7QS2nLvuTFOavCsKA5Un
r3JyJc15gxpDg3Oqv4uCN9gLt4eKQ/R5xnUoTKPTJOG30UBiMNz8uNpCaA0AT0tJtktD8x5rw8hT
486/9sxtOqMiX0vUm5NT4cEiDXGFXifMC7vkqqRT9ERnKpu3k7WnHJk3qxiUk6MIUt6dYbqFF2S/
jXtxkMWkZ9gESudXRZxoVUryXQkvHfarEsdjuR+YpQFWiH3f6M4SNiqGf69ABrBGNBMmhBEGCjsS
q1rM0RptjehnRBTdB6ZIRko/qFBxqwm8gRoUBWcaXDjWaor921EUsSVPzCEanstaaq+GJdRCai4m
peqCtz61ifOkZPA79qiCMKMgUiraUPon0wV1oc22SperJZ/mS9F8kU/791u94UTAxaQfd+ALYU3Y
Jel2QZDAJnRs+pPPikmT12xapGiVIAOj4t4AeIEGEfL3I3UBMKRdk8krOjjTULZSLRECSU/ilihS
MrWZbI+QUxhu1U6hQjeDH9NlXQ9c3IUqO5Jl25AokNe/nyCy4LeMTTVuH/aMtLWJIxlIoeNWzJrW
4j8T27sLsmTiNS49M6AsMxHbnfOlkun6Fa7UXy6aLzkIyBoYyS/Xtlmyjk+43UmJyDgCwp+3eVt2
IWGzZCWNA4xwy9JUUGSQ9Oz9D4yd5Ihv+KMxV9ldjdk4ntlUDf3cV9dlHT+yuwn65KbCIWx5ZGCy
LU2I0ImFL7Z9NU5aD21YRQaH1RQtgNAhghowE7OVYqnpOj+7c2RgIOlET8cLt75/BX4ZOZavxaZg
2anzGk2vhqM476M3++N3exq20qnGgWl/Y6aL3JobQ5AcrKltbr7K/T4zs72h0PsbSUCi3oE6z/EE
EZzz931khul9grkkQR47VVNVuDF8RY4I6yV+B7nHraT9AaPU/26m598SVdxNRtSLzXZggaXSpZK6
MLoAl6vRCQ9/dJp6zMjlqbuG60y9jCrJzU1yIAielezLGN1jQu2drF2t3jjDG0JPP7AYNU34ExhC
eIGx9nhERoee/qsRJRoJP6vZ3aAXU7+Kq5XLajfKIx3S8yjUc19mcJIgl757l5RwnSbVL+L/xoJ/
GBqcAI8A0kHRexDziODi74756x0r7mCKeavR82RFfgY1d2r66hBB0Dw4tNNLOaOpLhBpMh5S6PDX
WX4kshAiu7J+LHG5pgVXODIMgQxJV5UZq6xgJzQFwarDrAyaUTscb9W0KHL8ySbX4hmW35LwFxaM
/52G/6A3bWl9t1c4G0UtJPvGNGJitF6qz43KzAd76sYJUTme2Gh/sp+2ebxgrZBotfbhXnevZBgj
fN2PVSWRmSZUZJCulTrhjntUL1vrJZfGokKPwhI1NRYD5DXkvVtwCLy4vI0/el4+29o18puS3ScT
wVjXeGR1ncgJRGFwlccS2KTHZN6h+psA3uw7lXB7bvg6snUbR1gOcv0/ZHN8adTSoZ13nuse7MiX
sSfsRn2gEFpVClvQXSUaix/QX+WE6ERwbeFScZ1QJVxUVAVLGMieVQ+hyZ3Vvwtf+G41JtPAHh2W
45BMlkcrkQSmkmoi9iSpULo+WvAztzX3L/oX0G4QOXgobiXTyph5U4S5J5lxwl99flyLrF/ffoZ8
mOIB0zCEyMiKRyp0/fwDcqjduB2eeEJw5H6VwY1QxOdQiJU9aGSYM/fWa+ppLu++Gy+aB+ULeuc6
3SeO9vLRzULDoB0QdGQSxmFPC+HVrMdQacTopXlM3a77jldB49EKa4Hm9TU1yp17b51mnSYv0sVg
3Vzzg1ANlAGigj6hzaOD5GPliOJAXuuZmwnTnUoNzu7pjZGyVzcZTXH8spv+Y0VQ8xpEA6FYybdS
mtPS6ykHWR3UdipZ8JjHDYPFCsr22tqKdbsK1smRbJQ4y8Wxq8KnXvTaCDbgKwZX+wDjmY7VOU6m
J++KRAmSyItyGfa627/CbXpalpHijZvCt5RXb9p6ygFDz6OqB8YwfZe5esro6iXcYUJDx16cKuuZ
MnJ2+zUp2fyfDr6r9gV3MgrPS/tOezUsz8G9qoMgmDDqo8at2nLXepJ2kxLwddMd0ingn8rKQhwL
Tu3kjBOQj4KWcqR7XHcb/8N2jPaU38xwvphRkSE5k6XJpiyVN5VnJJr3T5zWtchp7D7AcU4BwDpD
Gt5P39a7zbSvrUgpgGRXMeRqN+Kpv9QYrVH0AXnUyciVRTR6jp8MhMklx53+wKX+HKW1mfDPqx5T
Lb2lfBhX4Ca9FyIiqlDP2cS6jbtD6/T3RLwZRllhlLjAKVig3rHlGxc8wU0EPpFK+kHG6D0Npv+/
XFlKecbracGurzCzNKzbpJBar5J4jTKAD/x85ePt/ybWFDQPM6JaD7v80pTkpStbidzIo6dlj2Ce
HvwoNGSUnTHLaqdw5rSKQRHELomhGdo+QHrbnGmnKC2R9Uc3ygpf3DMPSttXrQZ93tZBrbJYXPfy
uY2LXTrLxrgVQD393QRgwNtbTZ+I5dN9VsSSL/79f1365CwPZcNs+abPK7Msq9ZHKTcAJ1UWsXp+
ZgJD/81JfuQ/lqULlK3+CHraDq3yEHjsf/Bq5sD1o2isFknpUxUH6g5Imz2u3CvMhK0bcEJVyIjp
X3JEernO9lFaqOd33KHmOFL0tZLoWPUWfvbGDrl3nDyK0dChJz1DtrlZ6zbwnHEvk+8Bkmau66cc
glTVgfECswxgBRjn/3Gp4ZpCwG5z19AFEnfZgbgKQP1inLWjhtzWvfXhXwkmwyILbHbHN25WNuAX
1fLelaViQ1Pw1lTlqxVWdYUmWqMtYMTa7mH4Nbq+/kBu8z1Jvc5BJx4hu7C+ihsnnF/RsMOfB7uB
QIm6yc+Y026qSZdm8bGuRpYqycB54rQ8cfmRNgIVPjWvWDxrpRCLBZ8QUMHQet2I2nvZoL5IJGcd
Znou/CNGXR2vE6D6/63gy6Fk6E2W7CKcPAURxNt1rhYrWU2/OGYq25g0IdUsUnDMXL8+IBuspVDD
KxVvzV8i5n8BnV1yCaYd9CPLpDuucZAXL5FkuaXPCmdZtsySp6d7KQXiJhsFpKy7MYDXuYWvSah6
W5iWTzLR88s341hCRpgqHAncqf7nEV8OQ5VE+8Yvyx3OEwtZDPtmod8xdDWZW+ZFSYwfv5EUtTIO
C+9w/lad09Wh0stcARoAUtlv7WLnKVNuy+1sP6KlTNYvR4qR/NaGZpMbq+xOyH9agsGEpTfn2crQ
efPJwZ422Y/7JUecc6XopNuTNRuqE1LxdiU7mNrWFjiBSAeJEpN5uoOO4pUERS2u8+VGH7dHA7QQ
PtKmtcqOfMUfCxEizWG5fP0h2meXBd8RHjWobpuva/0jCqwSHPKoCnyajgsxBpwYgt3U7+Z5HH7k
zXvccYZQq+C3gF4fsacrOdPUJb6p9tLTyYwB0l+S/nqunXm3rLggYwwxEIEfUzsFlIumas4Fupyg
Uja6+7xiJJyhQ/T3C7+wvZt+GUCrHHAp8WxgkrqlKpIgbZclnG8RhST+0X7Px57Lin0/j2jaKr97
U3YvtxBMMmSHrRUeXDFk6UB9GIUe1DTe0jj/gi1UU5dlQAhrkwEr0B2EMxoZiPYC7e9U0PsaA0j1
PSrvaP6+ETwzQVZ2oMXGusCDsQJZJ8NVoeKz5kv5+L4DdDL90HDXJEtxfMe8jmdWQvR7iKOJdFph
ez1SaHsNXrvT7bu/mbpRmFUwYzX69OYU+VYtEH0UFQ7TsSAdhyYGmU/ggfXlstob60GpcmddIZgR
aJx7+97qpds292elx51eSY0VWuCD1DbDqQ8kY7eVuIS72TXm1GAYNj0WqmCd6jsCi08TYF1ffGp3
6/K5o+orRkfJWw3uujc+Xe4wYmYwegNZjmZru0Nh+Cf6uzTF4QB4hmkkv55fahyMwRS+N6aZBqNY
ll6od9VbgfSTc537ati3aTheBCNLciO9A4rK8z3mcxIzD029zghE+G0xy/Tm93k/FvjKkjzlB2uK
1o1TU6sOO8GmHuxNBwVs1ivNFcTIckGQKIAcocfxakY92fhSZlXhd5PrBZe3ee0G6TaPP3n7rSms
ILgzsF7drxEVRniTNfllT2zF7WwzySn7rdIploO4DW8r8Iu9sygptfLGRuc8l2XoBA0dDYEEiFHP
ocUWtXpE7AG8e+m20FM89vWIsONP2fQx++ikP3FiyAUUup1zMdYPGC4nLogxr9+js1BDIKI+hjlC
0NgLmQSYzzav0DIYnuHzHTpNxq64V0ECn9GJTDSzs/Pku5QxYk0ev2r4o2ZYQpg9WKHuJy+0hwyQ
z0XXBmrS6ciqTTbHTL2d6QW0ZrfmQ/EjOflffoDKI0t7DlHpsB67DU6Qgs167ku/iUYx+Cr9s5ZE
/n4z8VMOCBHZdkB/2YHG8nRxOz5Fnh9+H8ki0F9vBdsChx70ao76YsPiC5ViXwcw5srrk13eo6/+
CltHj56YijT10y/vfEmBFquZ5nmn7e55t1+LuwaeLzEbZ/52hrIReZFB1EZp0AB+9akxSOPJOhUi
CKQJyxLbIte0jXTx/Jd+BfHx4t0Katmkd3RO87EjI6E7ZPKe/6yhe9abu/WPLGEFXLmILbFbASFS
Z14SoAkepPAXaYfz/Saced5Z5KVvvCGnh+crnwd70d5/mhY07rT0lNTIZR/GG+Bmb8yRF7K29pyf
oUyOtH/Bdnx1FBhWJheXQpB1xezV0VZmrhdSX4EHkuKIA0nutzfJQbxdl3+p90umgSs5uiAI6XJI
dw8lHYaozBXcVT5HklNLe6ZoQCeTWDMND8VOp+Q3yJfT4yzxTEGbxsdPEQtTJJGE/NcXs7OPUCFM
r0i7C4qelF2heciio0dg2MbLyu+7VIPYUTFl5wzn3LjLliqCi5LDJOJ64GHAjWZTRzJNg8Qa+7Nv
CexYyZl5O+LNzhJODNuf1nqpbSQoOi/2g6pM8RzAgB6YowX9z3siKmPiI8iQ/MPQLjogmmV9zwN8
4qJBbx5Q77jElKLDmkr2A+gSTIig5F8AteyZXyhZ1NqCNDsSIKwvVaxslXfvTu9qp0UoQPJW38Oz
Dl/f53Rg8X+Jis9h2exfJq5ur4+89zFd/y+pFdN8TjoxOQIhVjV4DsJdaKxs9+hkThebETnFbee8
MuEQBNXgr+gTIX9uokvou6PJurkhstfKctkLwljB7zhd3EO2g2mTi/W+ubZNjlctQsSKGo7412kM
DRJSVYu/AmfQKYtzEc9ygG9xepfkuHXa0fR6Pc9a5MkIv0Dhw1TaH6Zk8G1hzZNPiIAazrmiLRU5
En3q+Z9rkFcW+8A94+3vvTKohZyRd7wVTy9zrwYVJt6YYQRt756/P3b2J2/V4dabhVZmmeSoHXOh
POsUGoZlzYeP0TDRSbxIxkCVf9WouTYegjfFkXcw5F9S48vEBdfw9nchRofQfZaYwY4kQL9fGgbh
ctLt0O1fdpgHuJCiYfZqfUieey4z3oVsLej5/LNEqiQJRZEUSkJhipmdd53rrFSg675drHCCeuO8
1YFJpPnY/4RhF03JvXrCPEd0iYkbVDA/AYkWaLdKpkApr5/aZ+OUM3Zh2AMB7QzeX9V8RhHj+V6L
u/ZWxyW8bXVretRtUgKnaBjmk0XUwmETcmAYNKxGid52LUPnIKDXlTzoU4kqfAL4FT4k83Ktbdtv
CpHaORbCYjh90fymUX7QNQwHxjKDCQFuCkQEyfTX6SzYsDUNCp54FOcxsmHqBxPKf+Sh8Kzr/S03
bGI3wwA/cxrUz+Elr7gYtDA9lpGIsZGuaI93v8OzBhoBv2lbJHqMaA+AMYG3EXR2n4Y1+PCSU8gI
T0F1Un7MEd7457EZISSM0ii0ZHV6WM5+Smd/qwtCCj2zfpBdusvZxEt9dCfXy9lKe/f9npfMGb0t
V35vZVcsF8HzCC/SwT115SeKRBJGPneJfEgWtwVlqxdaT1KdRH97o1RiFKrbz/z95o4P94Ao9HNl
0GGw+hX/kYZ8oAMYa30xj2/kzfFa1nYpN8mtS8OaxHBt8sl7dJSuE0mX7fy3fwE0CHK2SejoM9ST
VErb1BWArDZmUxTsp43/76eSCEX5oinvHjIQT4WKnUuOiRnG9HL70hklv0tNs99OPrpWpmjnVzOq
TdQA/5ey+6uHmWfh+sFnhaHbQpmKouUdqHzEisXMTcLaLfReYaW84IDYOVMGBkbbrLH2syEwDHQy
iSqVTOWNi1X2dkddpsH13EoaCNC+axJRgYYNqvMlrlmJPALYb6gt3gbc1XF43UEo4oExk7+NbMgv
NqZuxRFtserub8k/k4HHWulWQ3mSiQnflb9XkFGEw/SCM+mcxCEsRl8QPSv/wUCaeh7Ms9sTqf4z
qAHtXm6K5eb4Vsy4mVl4HV7RF+vWzUuqMYxcA02X9ZerK8/8bF/nwxD2ErOffL5kU8IJT9tFKXVf
Yffnf3QtIqRCU8F091AoKokGLgt+7bT+eL+UbZh0OI+jiI6S/SPFRG1+3P+cfcyqGBnNxs24Blg5
Y47AhjV1o2SwATvhah4OoLU9zEJ1PpmSVIvPhJDkQisIu40C+C7sjsznk86NWx0zDThjJX9E9cge
Eh4ZmXLzm62uU6mSno237EcV9eGVtLOJC0QFi1EKGIuv43ai2jeGhU+OfsKbokyN84sbu/XGNm6X
WjBByIRCAdSrMo2p+p9NbOcTcz9uko0zVvSF56RduwVN5jaU0sL/bQ57CS6TTPdjrOAQTz/zpaIj
m0UfUfdO6Z2zXnl7zffKztz2VS9ij0EiTAXUNFmntLZ+cfbuT7gM0UKKXAhUfznaD3vTGSxBtoO9
c/oyB663ctOQzxZDlF05LtE9q8bQLxNYT0P3OKDbYUJUmmcKDmd6xWgeBZWvKo2iSYiHqqeqVmVu
2ajziODKI1HWfllIwIBSBO5ofkd66+k/UUDOGBZKWFIIXZcHYSrA9UUNlojK8/LoZzL2H8TGNMYe
gQUodXlr5dlWXlzCteFDrU+bdqE1hE/giVLShq6jdt7VABPCtZ/N3DN0MSVFIcNzSZxsCNP08Y7g
Sxc2sc7Qk8sLrMBFoD6BMmmC7MXz988q9ud23YPWGwuA2tdAXRCw9e+ctOOBbluJQlYRTwQShN8s
F5GyzlqPcrbnzJN1bbvQ+W25sGUQkWsC9KFPsCD5F3mZlhvVQyfS9ArReOz263PjRIYUn2UANjOY
eVd++UszOeLlZ0zfdRbnjb+wb/zzQtDnNRmQhNgbzhn7jQlfM9N4dxyQXetwjl4hvc4YHzP3TYXI
UNDNIEAbLtlz+ZgLIwQQetXXpPMOj2ERv0ZlyK56CJW5nPp2AK9fM+P7MaxYGShbR/40w0vzDTOd
Co/WrKq5/yWCWFM2BlxE5tXprMtd7V+0kZfjVucqDC3dCmKKllw6oDAiEVbwmpxYGuJ7gei243Bb
bjbvIlSSbkD7ll/uoxe1CRMMlwXDu1m7DAFa5VGyeYyzlIuy5z1cNaoqiMrPpQwZIZJ02FzWP2ue
HIH+EbfioyRJzDLfdJbQHiS0zNWwoLaYRjzatXVByDpXqRBQ1z6tmijl6zaeeEF6k+OwRUNgiFcO
slWbFPZULaByhDZieYaqY5P+B6O02X25AG3zCgQxjNNL/l3zR3Uhsgxa6lgMHrbrhfaAECf2dpDs
eOo22rmylOmkvUClFebhk0O+OgedNGCCZmptrAHkkA9hS5Io0NyNtapOMX3bp5d+APKkBdfW+l9U
IfDeGxVXuXOcLpxL9Rj+H3kYL87TSG6BA/D/A7WHewMRJloYmyWDkeD9U2R+ufvfJrE6mGph5fPN
zuAFcL6uO26JhPJQQwk1ce3PhVBXiO8F9gWZ4XUaXqsNTS7fCStMYsjbNQw0+W4CtM43zuO2Mz4H
KmxaH32XgIJatm/MhYbpJ/0DEMas3vepDXWctZ3kFpviGjB84aT7QzfEpuG7Y8RXxGWVOPWQn5NJ
lntVx6zHx0d+eIibAADwQAsQnpk9KsBd32D18lWM44TbFWHOLMSXi6bMYPcciPtZiptmBvWxIKHo
gnb5iRQVDASnLmOrVcCmrjW6bfvsvlrJtib7pLHbzCpCAm9TYDaG+9ijzKNih6OK1G7jcn673HTo
IAiw/5rgrnRkfKURh3M7vawxH2e8plt7OxT0fWXmZiHzu1U6KSO9787KNKgRIb+69YEWdi7OfVkq
Q2QjLd8YfzRt6Vfsx3hBJqky097yHWUyKUZEJp/+PBO2LQLfZIoNNkbebjmpFttBeTYp9VByPuvT
uCdTAPygNEWp8da3MCY54Wmvpg332pAaEgBHiOW2FtDyEP2GVxdMHawYWL3B7VA7wdfdirJcxQu6
vTCTywI6/4VX6XV/WtVuy3QvfIcn02nLw405hDRiYoU7gAHOvyjjZ7WSPyMDPtqCrD94SilbFluX
a2CfL7cyeDPbXxXJPR4C2wC024MQ6RQk3rkT0JVLwUdCQgvGzbidDZGQGa3XxSSnrZerqSF9ARSD
B1QN6AP/HwiAY1mLIpVN10Z7C2c3u0x0FSQbQzCtfVNPDLkamtHG9bUzZDRksSH/vsk3RYusJ+Gi
iX4Snkj11Ze6YaOCraj+Le2yzkbuO07hoyDbnBF2BjoQY8Xm02GMqmZnrnevS6ek8x9+u1kwezip
+8oig6YjIdX9MtmVS3pASdwoT3pkBKfVvVZroPv08StCYODZNkEwQ72wu18VDGzvXKGvuJKWd7/P
498jA1TcQAqwTctONpGwsoDYS7wHeD8Koj6bGuNGfcCkmFrbGyAPFW0UqdJfH5Sklxw8tshdSypz
GbnM4Kru9O5YMPXhl62qDQax54vxNTTTBuC9TXvTZEs3ewkXlZq2ccnwJLvHMXPYZVuDygUrhsin
/4I3dcMFvsKce7Ex7RzcL7OjoNcU5rz1vCMICWYsAW63GYA8Py8rIdv8dmsoVJ7oM5ueeLEwHmWH
Aw8OyRQ3b1uQCpSPuLYlSNGBgEIXLtBJZ3YAjXWQO6cm4BOoEilOpJcu/wYk8FEKpuyZeOqEFiv1
+dJP+wkhYYKQtNsprSY8C9VPA17GMYe2hdKihYA7RaxIPbSxsAZ04SJL0GifNsbefY/wEsXf/a9i
TAqjftAs7UivuuvASKF58S/rAoYstVME0UbnaqIIrD4YdyE6i24hN+DMCfIbF9CWV7NdZHJtFdMf
dpgaA0k2RQBRwn4l2P+bEGt+nyxVUlK1wOAN7TQyGp8RSO122RSfBo+77rL3ut1p0MM/EOBF7lOt
hFjIGzhHpIc48e3EgIhJNjSIqWRcAXRbcQLGixtWY9ZgBdksvS5DyUyPI+gjAAVgeNEVFryQouuh
6VkEL5yRGvDN9gj1sgXZqQ+iF1obuIqpJhGOI2jeXkETdGgIKOje0CLPD7EkC0q8+pxzxlmF5TSw
ogY3JhLSdcNKEzND9M/wqUnYYCwGE3iYRMnbfW91m1IckcEuML6WY23bVEmb3k3kMWNXJcnQTOXi
k+SAHs5LtRZIIXSPm+l0sK5Q6Ltocyr3PhV59/hP4qh82uP8a9cRv6V1mjPnHmPCLRTeJNwFSFMU
+A7MLrXTvjFQi0qeEkYOX69IMki46uJst7PRIFYKV9pywy4VEckyIFvKs/06WBLWcz2gfHh+89lV
EJrdZcAv0vrT7Nf3L0+qZYa7vhvYm3mQyy0qYFrQk+jxBbSRbpeuObBLEYgirv69fhcMcQEzKKVa
BTznjCD1mJYa6GGVcSPtaL3Lg+r+fkgDBWvHkTOrzKPl3PP7WtusYgLSvHc/3urVlhx16uQ1GBrH
Jvw0Iy0KStJ/6PDluSNRyAX8EnpdgHI4WrMH11PZE8y+5PvjaxKBSX7GpXssNMmYfT0SRqQcY/n/
lZZQZ4NLWjgTbWX0kUmPn1NQ8Q552OxTvnR5wgSc5hw+DwRjVtOBSTm3Sx9ByCL4IrHhBYtnslSV
YOPA3IZB5BnzWpWIkEdlIYR27oHBXdYIM84EoaOcKTpRk/rWuWw/VVCSr7Dw9ip1bdSaTSDY2CXT
yjUVMVMVMTEw3WImZN3hr7580uCR6YH9HmxYL/uFiIz8HY+19DnHwyjce6iCa+uIti393RTCGB4u
zOh4MqdL9rjA/gUU0P1jkfffEyxx3OVNtfUvdk6W7IzJhUoecFvkLYgsBdgP9563HEwn6MKqOhw4
Dc2cUM3KuJ40Toe3/gxN7LZWTrp2rky2C+A2HP1CgWaxiIykYJMI6I/iQZPzjeuFIcgEDmIzuR1O
SB7ThshFeuMTg2vZ8ihYOG0RxMoSKaF2r9arwKB91uLXa8vb2BCO6y+9Q9NzvOlJ70r9WWooepDT
0ORBw/yTeTWTmFF58tXNirFK4eey3Oiq3F2IESiIREIG5GxMnqzn3QfQSqo09eTLIFl3YfhoNyr+
prmzlAFbai+otsiVieJUp6AKboRfYre8XcWqadWtq4PqpdtvjePhBUfrAciEPmCVIFcwPbO8eCoz
Yo0A2hRdW+xdVhoeSoWfC9ApK1F/hlvCBPQ2mLycH8pAl4ZSi/A9SXNkYH9ppzC5w40CdfbjkUZ4
8kmXANRzZaerw0KYtK0Exl3l7iDI8slYrF05Gs+JY5qloY2gblrlZ8DN13I6kilXUVAOD8nhIeyM
eFKcc2ohvLK+BAW8Ahlu+COWNk+8j0B9dPe7QrNOX7nTusCZ90Ui4quK8sFQU+zh8xMOIEVw3SYw
Gpx53q4oxE5WZgLMM9PhgwylYYNS7KQ7caH3zaz9NcUjiNrecYw1dxlo1i9nLYEg5VPckZLmIvYQ
heYANGVlz402+EzbpOSyMEGT9sj5yeIXJSuYxtR/7NYSriBy7L7MkNcxuCkwQZ06T8b7f7Wh9+Ft
SgLviYxhE+W9fKMdxWLfVg/q2GBtnvqqs0xl9ua4JZsbkYcqzkFHI9c6yfVbFZ0MvYfwOiUym2XD
xJkQAE5vEiAcPVxcUkiG9WTtFJ+uC9MnPdzuMvUz/9Hex5jFX6sv0dpQTHszQa4y2Cvwxcyl1ppK
/q0PCyvyY0WUFs0eGPQj9ADyEqiJGkMznVu0tC+Wv1asgcFbf/mN8gwgtg0HaW1dpfuwfpghF7q8
TerQ+p3+TpFpj2tR88GT6uI7URqoFsShn8QZeD2206zsTiOexeJXF5azb0cG87ZcQt+M4O3TOlLE
oVpw97/njpa5+c+EMY6SPXtuAD0BtSYQ2IAgUyOEeTZJXvxxfu1+3D0RWcSCYj0HEa7bstx+MYjX
ZgD6OxWdRV72nssdYSDSCKqpoIZVQ3us+Pq+Lc1jde+kTopu9qKSRUvtm/rNz51oZytrFEbosuvt
ciKa2v60/v3+NDlc5syYSO3NFaNDJBGlPZmJXyvzyMCjvlxJk6l0NszjYfLpxZ197u5qzBIhJfp5
vjHj9dMUXIk6SzpaMwiQ/XVgxgO/KX/9+NdYWAXkIUeDd/UbHt6MhL1miVlHI6p5assGMge7vEcb
OY4WZeAkdUy9XmtJrAiN25wL+C7UCV2alF3QewrWs5ow8aD/tekpn3MQB5cc+4dHtTGPZVpGPqN9
/VBks2ynsUi8CBG3THr5qYnznK7OCCSbu6oat71BpjPoRgLwhFn/akB1s4c10lBLYFWhR+UFdBVu
X5TwSnKaNFNpQ7luv8UNSjHGbb98JrKIAErRGkIMkhwwWIwCteKRBpjF4HSBxiObwUsJynotqDq+
enmQLD/Eno/4+juW2H+xxPXXHqydag7IbNhDd3zTz8YPyiEdnrFBYRdiZxZGOwliYjQqoaQUMfsI
lWQFxoV6RNeGrKItLBDWH1DRcS/ZLd3PwDqA+yOIWkoKm2cu7decP4NNnW3eZGYyaMz+tw6uErve
pS5mq56AB3XKukmUuX2IAI6GRPKhsmxEVvozt6yMaxTMc8S5CSgUHaVhEofx/nua4gl5LJgmt6nE
nWYIxV0X3E1yj9kWdiha/ER7uqdPP8Y+6BEtiKt4+JJoTin5lQ2He4dGmJQABexdVonOA39zOwhg
TERLXiGeEI/XM/eNACBv0/DD4BbpAssQaqJrUkkMiB8pFJhOeSlWtiKzUx47ZIJJcsAsibiAAVNd
EKiCsK8LldWmlNVDl443MXOthTb/NwWcLeajjcEtbFyZO+uYZzRrXJuJDPMbS395wSEJyZM/zmvc
y8KstFk+OTqwhk5UibQMQK/icuQ5xPd+E99pLPKvq7dQo4jY/Niw0HN3ql5b0Jj1gHdxJU4rYEAn
gIkmb00doa9FPFhm2E++JOvY8nyk3+igtOGDtd1MEQkrSv4QKKkkg8toIyf9Wx8UcMNPqhCg2x6U
IemHRBXEfuZPZGZDotvgmj/nED6RSroIYtDYLbYOthhclf7JQQucue83wIHTyPUJAo66Nrq4Ti+P
FVzpanBEzc4ik8s2B+AgjT/3pgjamKIeJwCBNp0TR6CjwdjwXVFr2Oizi2G1Sq41vRSOqB7b/+L6
kHvJZZFfPC9zWYhUkgVwNjHCcKdhRxvAsU7FBkvqDUxWNCnw3ED9Hxi0czNEezASBJkA7DvTWqlT
okG8gD2JsMVsFATZKhtQDCXe3owhkcXqOmJTVGcTeh+gIY4efeytzVSK9iQfZQI0kq4uxX5tC6Ss
aYHmH3MjCxASIeiT0SYETOpYVC0Hux6nGmxOmNKwv/2+hxz3MUqzyG5cCGRCqFj0puL7UnpJ5kIr
JyWllT8zfde97HdV3bjaESvUtNGt3ccdJlm0iNikzPN56BRXJ5N6c/4sl3LxNx04WA1NT3lTVPIY
3I7Ic44sMhDSoUKyHtnsKgAe1Dhj6pdz0TauZ3fzJ3FQXJHZ162hw1BbvP+2OAgEwgK3rDGC1cQU
60cESiye2XCwXB3Y9MbeTrNGqCPRXQMpKvci0rF1q8cMNHzkW0g9VD3qEjT8VbC+yea4C/W89Kn+
7avlGwFw17agMSy5h3pTMjv/el9nxcDUbjxgItbAr6v/gtV/z6i9F87uYvHLQR3oeds9cuxyM3DR
C3A3ewxsjCe170LSxU3I+O5B2o1Q+y0T6G/WMBwXBBUqdK+uOVOoTGs5fZdlNnLRJBl0wRdtNRCM
h3SFgIwZ3Qnh/oLRMLMemsWkxxwIIJhGMvgnRpY4imQ0WPRmVYL+cEJTJI8uj9+Oh89tSBo6ZunF
2XGU5tFfD+Y96c7OjyEpFUeyxj+1SZORUw2J/K9wZ7f+o9LWJcq1tO97ZCMkiBwLtuWr0R/tHA0w
ENdpI9Xhyvz4YghAiOsIHPx89ylIbwUZJfbMJumRQ9eYsDYSH2x7sZRsBqkNGjaOsN7Rzhu1Wxpk
phu19/1THACr+n7ZW8z9gK6qFG6tsdJijlSrkfGzfZK1ZbJnhCg5alRNL5ZCilmKMLaG693HhyIK
iZkm4zksLA8NcD1WUAUYcBjZCWqik1pT53Zh0yhrsq+7UJHfN4XjgCRY6yjocqbN7cLf8UsBUdTy
AA1IxBOv4kwVT4fiN9oGX+334pb5gCBrPImQ8wfHcAX+Q3GL7kOpzdbh8rBgqZ4cFBF8XZsJybKC
0tn/u4eNLHhlCuyppDq+JgqE6RIgMLnymvdAzfzsmYgck2VmAruo+7MDg9RaG66m+dfiwim1ujJL
nLho0b9FpSvnb+tJg7C4wpce3o6MT/AUCfW6JzXWJP3LZeeB7hz38nVjcZFQvUpe4o/nFiyXWMoz
WHaaV4j2YKgAuXGwhBpDplhT37quqPQTvqA3Vz7ADhYbBXwRpfS44M2iHIElfHTJDOT/ehuApP0b
DlfPaGCkRpeT/nXdDd8YJjrXgVssmUD0OGNuq6iB3w6YOczRgMuqduLXvE1KY2xTA7KB8ZPoyw/W
AwdMDfIV0NGQbr6bS+e2PFndTxcljIgoslXzOi5vQJnwhaummtNS14DjsPlDX3ux1scquLrZDwl1
rF451GdmeuDIg27+czSwWfqIL9KFBnEdUCWHingz3GUz8OcQu8ofLO7Fw9OJtUX8COSkOzO+PVo/
l0mKWkzif/jlraE0YZIsuL4dABKZX9+7Eb+IJpaY3V7LC3gCvyOmkl9m4KemUw5jgEbXeTA+gZEz
JPCMEKOc3729qvuIWkLSyZxz6HIp282EC9RPQZv2tpkor6a0gbNBTtBrmi3jDhaiq7qwOKugHKUn
qK6P3DkAFeXVBIkjQfz9/L9Lo/OEb/Yhp2Z7vhZWXodVs4Qsg/XTqWZ7Nd8An9+qd4BEVwMxTJiM
f1BJtZNsxPJvnhI/2+F4t7C2PkKB8ujjwAWsj2NUthmFoyg43VoPHOp3Fg2l7wqRoELA3S5xURDS
ci/D2L/9FvM/7ELe/zaNNPtEZ2Bo5zgHctma2iWDdmx60Kare6VRyWpBZod4Y8bMiBmDF5NytG8Y
yNJRuDaR61Xe4jTwcxwdcjLoPP1cABv48BZ9inHXZAgCxskrCZnl1iXRqQBN2NlkJ5WkO/m6sa4V
hMjU9ycek5bE9JU1KajdAE7F50Z0x8NTseNwGgJvEXLlrAmCx+aBq4QWbErUjmywUSInswCZ/9kH
thOE3NmTB/fJ7GNYkHZzsong8gLoF781Yrp622zmMoo0LzRRJzDfviwyjSLB1RfYigkzRZEG+MZo
qAdlbN5OQtn87biIcR3ltyGR2dp5GdLP5/K5MD2QUU+ErxBI2zD9iRwpWSzV7YPK67FhHMH/qc1M
gVfmy8fE2RyxpvfHrN5zA4zyudqn+Y9RCaRQB5yjNq4XHFKGlm0GU4o5EpXxf2KvsVzR7/7K3o8Z
kzK4uBLiSptRzBjdxHNyoVx0vVCCCXn44k5oj9TgkVAtt6db9hJM7xuyllWijrSPrxugvXGzXSKZ
30oJjOBrLRv0IH36KCvVcPZwrbkn1jwKY1SOQQX4Rw/rdMGWs4vxX5rIejtZiBgKBFoqLwqF+eVP
Xwrt6kC+YSJ96klgk5TlG+4jk/AYvGNPMy0qHRg8kDtRiaaVVDazWiqL82S4bR/rZUmhOkrS4gIZ
w+TZSjV1SPdKvjwVR7AmAfs7nzw97eF3YnvnOg+Ys8SUepU2T7GArA6opAJQm7y7uF9L/VHObaqE
Ndbq83Ufee8t9exGPw2cHYwAN2ctUtRCkI6rrqOpVEM1w5LYBHHNnDEsLPnw7WCrU84N9b2k4WT6
0c3irH/2K0NMcJoXhq/yAvyQpjbkndPL/N+M8Vre7BINEq6+t11IJQJIEr/Gvc1+Sb4jL0jPkoaL
G+SETIPp1HtE1pEdh2vCV55uzwlhYZazvOf2Ms7RrslRRwzjV++IccEZXsXQE7RHGdmqMLi0a02x
kMBkV07QjCfHiiVd8l+BGHxRJmx2mCt4vJetG8UqvhcsOaI43T0NIOvISPhm7J9e8LKjvSVyRfw7
PEBhYDMDVyTttqzPaP/rlq5J3HwqohLlD8YMInrnvjDoyDWo2RItsmX/GRstYvJF+ubC34CgBW/G
EOzEppuPsQigxNIT5aHg6kl2CEGFBW0Sk3S2HejF+QxaDob4arFGqJIat35gbbDsej8EAdIyw6z5
nkQYEeBw4tOFj0JbyJj4AOv8stNeaXe1DzxD5J99XDKPxW/W7HHNCNNuirZWaRV6HSJ49NFCpnej
F4TkPWZqmeHMhBmpCBbj/7BqhY7E3rSKCCRuQRH58KdhmdhvZFibYi8kunu3VrPO3QEaDuL+bJs0
dALNfaG+/DfazDoFMuvBGKSwgBjE5493+F5n3w9r1rhTNhFNBVv0R9EiXb/a2MBgVzsSylOOG/pY
6q30i8289KsQeTyHumhgIHOzOpVQqzqq2XMe5ODWiT5CsRVNw6/vNfDUXa2z2UqEfOgjRGV8+cIw
0Mrsfopp+8J0J+Z3rhN5jNojzfGxsPVgLM7Gcqz7ujflnEoh+0Udk0aNRyL6kB2Dd5EWI+W+hjlM
xdnsfsvS3pSe5haHzZCX4OEufc6KDKziCiODsh5o/aeRGzdph/9VNf6HkK9mMprSFdYMIHEVKSZ9
rc3IrydIjwmDVgbVokQwlCHSLtp9C+jvSCu0Z/nmt1HaR6Xv1Nd3VKgvsbGWCwtcQMEHbnjnmcFW
jChgFYbWF/O0jMxMdjLph3InsrHojCQ9tm85w9cZHQOFn+NM809CqdZ0gtfFefxKSOpGT0jqQkaA
qXXab6BHdoRnI6+gxuGCm1nUNxgOSiRTyDgNlS/oAi0Nc4a00PUrwQHKXW7SKwMmPw1qNhAIPNKv
pC1TELTgRYuWshOzBcOlEiWmAQI3Hnl04vFOYcvf5HRpDgMvBz9u0nzJR1nzW4y3AyEvJw8AJSGW
feAfifc5EirgS9KMC7Dd4a/HfWo88ZsTKhdGa1SP0alxH7jHp1u3pE3dWO38NeNgQbprkm0PsSBx
sf2PCc2Grn8aMmwY+D4Z4+Rd9UqUEECgZnh9EstHAYakg1XPq6oJZytI8NavLZlSZamS42E6BV/6
cjwGz/BCShugHQwikY+LB/dn1t6vczgAiB/7DB5zc7Hj8xDiJsvGRrIXmwbedtugR9cTKZvC4e8H
pqNqFEp8w3+Yph81qtgElhpc4xZQ6Ko/CQidMoL7qiaExwj4w2uMDoAURpIPvPJaZQQaby+VerUo
sHVUi90dFYRk8ZALMz8KGHvmPq19QbEWz6Qoae3X82jRPQLmHOhPg21yCEVT8x0rUuOvUI9YNZYa
4yuoThAD7yRZ21IwZF4pjZIx3Jqzl40fB8++7KY58uOnLZq5IRdRBi+Yp+BjmICsUbZTLclGPa6o
pp/r/raSWRRwRK34x0m4GSRrl23GaamxyUfnL72y+yDmeRoIiTkUrjREkfdwqWnjhC+6tpCitOio
KKSd0rsBl71To+HsfBn/vq3BFqtnScZs9o49ihu4kvkgWM2aU7HlakgWzPBD1d2ZbIbPby9UAGMp
dF0Ujum0mYhP4RceUd1J0wJ7xhyMhWe9WooTGLgCLgYVMovRd+O7ecjb6HATjeeGwi4UFlQ1YyMO
pIMSTIfLzgWaNqEW90vEIk8FTiduNON5yYGsGD4iw1y1Tw/OutlSy+SKDsNNd0U9k3+GlFt3CqM+
ylvl9+JiHhMKplHZnRvQG84UhGszys1KYr9WgnBl2AgZUCprJZaVNfUbSKed4y4MvUrA2+Uz7zZT
xZM9rDYaEQNTQSx59NTHJcwRuOASKFeSPpTUfzsF16uUazLVIDWMHgYyjEYOybQ0pZ8y+omAQsgR
jPmZ2BdRxo8/nhdwbIQIWUaYyZShuUexvYu9CoMhin09zVGE46jbc3OcsCqzC4Qut+wjURiV6y6Y
XfakxDd6rBMJDYCPuAFc7YYqN19DzZnNLaMpbL6aqN91E7zwrlRyRxP45Ul0g5r9Jfv3ngxFlNC0
6cHOgk0EJenUtzjyO8p09xQliX++ZrlMsdOptZ8gPkkFwL5lX0vYZG9NKGSW/gC/6VZcpRLyvenh
gVkUhhK2mXplhnQzmKx0D0ijpxSmEStHCWwtjbrefjKanzzT1vGN0FM3XkQXkQ6Rw1wdhINt9AuI
R/boEMToiw5xIN2joqBBgW1wcprwxAGr3f2gnEtucsjd8Y9A3El/yhFf7DgHoe6NXmgOW/sgiIi7
Bfi+f1pwt7NZSEErg4H/mtcsdODpcW026Y7QBh75I1bGi19M+lT+vtMguDtGxlbBxGpiaB8tWtNg
FLIpBxh0OZffX9YGzk1Lb7lLNiNFxsWxAUbziZC1Wcxy/TXtXiEL/2bogxjNFGPc7MlGvs8Neeo4
o/aI2pYqDNOytZsHcOaz6rgOGe9Y7kc+zDNbzd3dZnhSXxOSDjfNT0N07IMv7tpNib4NnsVwEWP2
Y9eOZ2qwF17s+mykVS+yj7Y+WrqG0r5EsZfnTuEHGf17NlXIH+PpZXkXak1boNXGjcJn/HlBrorU
1w0D832GaSfC7dfhL2i/s4q3j9/vUkBGDoz2Q32Whfj/Emghbx5KH96aF8vaYpwhcKKBc2pKHU+Z
uX2ml1iQ2a1h95DHpuEGpN0y1dqEkKfMz0f2AhEyi7nfT730GinizlYgmTqOtUjRZP3IG/6UWXtP
Ohj2LA42/I83y8Ue/hn25/UM+Unbtuarqj1AGamoDXAycfEr3SNPUUsjMjgsfq98IHa6kxhv0a24
Px2AXSDh0IFOrTXe5/niJ84RVp1rG/89KQ+6wuZNLfvMi+G32WjjDhXkAMMuTxTuZfrak41nX5v5
Fe/ZLVLouh31xtOGkzTsGf89w1Bv6h/j2ObF8t3fiVqe4DLVBvKxSoA5u6qHmCbF1Dx/26uK/rrs
3BAyGOxMIdMj06Bg+jatDRQ+j5hB4ZJjSjEWthSUQgwLweo90DMQy/BsbhGf+EKJqDNfJHGGSfli
byeHDscL8SUEUYDFdpdi0WX7aOqyNAumx6OuZtMGM8dUB/dCqYioBFD3LIYrUBQf5LH2HUKJKj48
PkQUvHHpIxVq0aJjGitMYqp3L7c9/ZzpdZOBxBF6ViUY/NqwFg+UDjICcbu/XsaMDJF3v+9WNXR9
932Yhp11hAJjd1QSmkNH/vCFhpW1ZoLwLL96pWOtOL1VrlqtYblLrjTB+PKpH9lJWSGdwKYx5xxY
1eRom5Yir/m/rWKAl4LyVs+RfH03yDYs7Ey5NdSh728ROjrOosUrbX2SjvsDbbCSPTSnfjlrYyLf
zpZ9j2IrzvQlHdPKb7/AvK5JoGhH2T/P1s//74Q5bXdip+3reWcRRiZ471H4BoTFW6vj0HQUwdqN
WrNBgQVsOoucXZRbdIIT/m269JMPTzDE0pWcVRIhY0jS04WXkHiDYgVUjxrpJMdJJYVkID93F/R/
e/U5BX3TZgGmqoXuiNDCtr7xKnTBRZiH6f9++jYbrLcriQJn8gZBJVOrVVOd9jYApL6ycIJik3tl
xFTpWYmZAqEOgD58VR0XwPiZ358gBAB4IZjT+ecxx0wPWMx7Vxro4wERMMgYkyImCxAHiC8G807o
mnn9oZdGjme2Fje8DCJhCWISbTLltwuSay/N1ZF+eXqaYybHZ/UGanhbCixqVuB18MLddzlYlYXo
y5DEjPylYyXMEWYzCpkiLfupJ4ebsZIq+oTqPzC/7xXZpeIKIJSy9+u38Nvzy8xRE0wTvm1t1XgM
BgxT4FfXjAgELeVvoHsE9cJgRYk01jirxee20SPVS/I1Ghdd6QGLXDup5LYNpLkUExSEWrh+abYm
giI+/n6s4k68tOs87blEtCOap54qj/eItrV1zeYmdoCTNU8d5wr0RFMPFgau7hfjlXf1Ie4vi4F3
PoJHZo4V7Yz2WVhaVyNvbn2YPaD/5LybYQab55+ODaRNOuQquJvePuvGk5Pl6JN/I48zONRRn/+E
1DKoaJhtAhJUfDn3WKHks4mTiBhvu1JmWGfeDRP6PcggzhtGA9BwaoTpoFkFyIhpy4291oCGIJab
4Y3IDIn3CB5vaHhv7eNUzl7jvCzx8OfzPkxLlUV1erjqkSStvGf/jo3M7JiGS2hpv0usHaT5W5Z2
kfpzMX2fhclsdIuqJLyTxebl9YihbImPFEDfuQ6Jcb/5E/tN1bz8uqX3/ujRlLY+3lEzTEca4ZU5
9s1PU76WyOmdsluh+IHDKsZ97u77dclt6zmS2CGorqXqSsfLkMDXCOVeUQMJLTtVMxS3GHBVOH2F
cUAukvoFL1kmpTD/Pa721a8nHGLe4yKSdmi1oCk6eJaC859b1+rMieJwkI3dT1JMxBL0dw+Wyq3t
ALkY/7cb6+1NZjY68mAl7TgIJb3arosh0TIp7tQM7LaxPBtdxiOI6P22Y+GLF1WB8IdBbOvYExId
6pHUbfiub4d3gu52Dfd0H8V+8qwM34jxIoXpt4Q6NhGBUx61iGTI0pjNH876Ny6eWJoxhb2NObQ3
ZUAJQ46rATgyxVRtc9pXvB79ZWIScgtT/4SgzZRm1Oodf8YHV/sazqAdIEe3nwXBHYg22HHuR7ct
bxnpWO5FxbMdStqojuL5xMOTlC6dQjrwP8/d6/HgaCABegfSxM9ASt1xk9a9RYTpmborHc+FHF+7
BlZPVHo1vd/lTxeMtgTBMkVc92A5/dvn2Hupn9WJ4sot6RujHOLtsutr9kcFn9o4qVckDDTIg2Ug
OxZnjPGd2VLn0q65Ub0SQJaOSTSyqBDec3ggwkaaAocHNx+t3TvkLGz9HRVjUQOihfiDepCncHD3
DlNyVqN7VBLkAKgMLfjIaWiN/306dOqyC5NJRlXC/zKn6MRXd087KRO8soYSas8At8KRDuSacfQI
bG1pDmSjhexOgZEh5vMx6HpkkSJNZbOqtPwuovOLYp5fCoRgr0Su3bBK969ZxedR0NaLiqt2z9kf
6VZx+k1lGony5QIhnd85Jzlqh3yYUjuMtHdnbWb0C6Fye2Ibuzydjklr+nUAiSOzk+QgKHLJvZt7
uFS72HRHBmdvx8e2cTm0eGHAY/sMo6aTYQI/DGSqJYwBifixVLXuLMwv6fUZcvdqq5VSjrG1s3F1
PU6mBNq+w4fKYjUZox1bNblV6XMDapnZ4ijagOoBY15dHeF15IPPs6YQoK/b+uccf5GtlHrJV1Gp
td5eUAoGz/e7S7uCBC4x2dhZK/qUfHWJ8g/kuE8Jqfjw0TokJ045peoZEbcQZTPgyrLiJkJR6w4k
jNxkPDFAYd8/WnLWc+M9cmz4zDbhnN2VTMpChMaTCgQFDYPmd3tYoGU9DxfN3OEnXVD6DN3zH0Fy
coZrc3veouxFk2kDY4Ee4Q1WfK5vmBg+C85KQZ0YDzW3/O/JavZxeBM5TZdnO7LlaCesAfXuMGqU
IMv/6tiMx6HVg9h6sLVZ1T5wqJXgWJexWTtU6dbhsnhAv89SNxw6b/HvGW6xj4d0BAixqwNvrnkf
vC8RvbMEeftWuB65RP+kX2Hl3tE0+aIW5XRljH2eM8kt2vm9cJXnF+iXMgcpsvE8RAyaeGlqlxSM
Ts7X7PdlV5FQ9Kncwzs8FGT0BfIXihpgJoLQfZysTiGmE3Dfgd8NiLOiTUEaNps0QAu9iBESv2AS
5Sy2OVHFpDz+48tZDqAY513AiNraIGxZZ4epWvJrRRUGwHrqcqMwl4V+F4AIsT5mW3LfSg2cm+9+
hpqYQ2rD8m/5vxormC6qAIXX1YzYgr2rkQjm4aOPhUCuq3FPCvrWF86Ndz2+E78Fshw5Igw6WRTU
AShCdB5RBjr4fY2jX20omum0HIaMzoXH6U93MdaLHVmgzVahWn/M7a5ZOxf90lTi0+cF1ME4ppjD
56At1vpfvQDWXAfE1iUpKYcTrKhxCdbhB07PGm24jhyQKeOII7TRKnzFbM9Z0LDGGPIDnQDhFiGn
BtM5TpEEDwmou1hLyWB5bp8zPIrg0Od02Eru/dO1CaUbe0QMx6IQzEBx9FnzLswwCs84VjqngQdy
La2Od85ryp74kYRak3WB79md/3PNTIX1kqAGpHdLzsaN4V3XW2uUX72flcIQe49Q4ueMhoCXi69y
7VNwcUiROOX9Tr3bgQqeFDBd1z8OAzdw5c45gaUqm0hxDgLCZBAg9vlIWpY5CWKyEYlUcSSMIAXq
s8LkBYt7jb59sZDwbtuxYH6rKXOaEvswE4kN8JhcY+1umWe7v3/RtImqPzlXqL72KU6bZy67hE+m
0VB/mzstY7uuOYAYoy+EFd+maM6mY12TK7QhXlNdLHLwH9RM7rbPawgxKqWKKd/5cTWzCsk7hWYH
+9ZQFEGrszl+xryC6o7xzafHWEJpczj+gSmhUGnljPqi7NYMXeL+pelR778FWfneX73tNWKjIst2
FsDRgPVF/AT/fNJxL69k9m6Vixfwplrm2/ot1Jcu3qdWj2j7AF4qo9yZvCQ07RItakp5lTumYMjZ
NWg/QX/unVVF0yAjWYP/OLWyL23pkE4MZSWIXgHpZ7TOTswXwJDCXjbXSiiVDMeRpOj7HV/MgZl4
5BNiA7MOCVE4oLLz6UUZGcmMWLm/R/sXokJgURzic8y+UAqky1XUeeJ5oEdYupoOFmhkbtw3CToB
ojP5f+nV5Nvp1ZNM6KsaBL9BlGTip8Axm9OvpBcsG7nhM7VC6R3twiu2mFZ5FaPUZfmZwGRi/lN7
XzM20CY7MwOmvokFYsY3s/xM/GxDwpMTFFXobAbXo3TNLYzsbn1UMli4G6zNvKYgslaTXd2L6cK7
mUh7hg4HvKJ0WdqJgjxTdBsHIWrEgbVrLo80+1/BDxbWpo74DtAGEl5afVOKiywY7+aSmgmLTpVM
FgaFP7fhrRGUrXBgk+U4vKmcSSuGebjQ7tTuJ38jTc7YvtCSYBwcOdux9iVp3I000dwtFWOd0nD8
Eipxi5TQ8GpSfIiPmR9WmxCb8Pux18Z8FsN3nag7nF9PU63d0bkTJY+Emy4jAr4hBFe91mNay/my
jmzbTuoY1j9WdEStETi1UjUf25rn70jNE76vH5kT79NZXtjdq3Gm+8ZmGg9iI7XXidl3auxMhizG
LtFm3VBRbTI7M1yCGhySB3ZxU9weNcbEB5LztK0Qz5m64s4ypqge1kHRcxyE5DGTlNENedsRTDP+
iaWwK8y5gmVYV5GVsYlv+dKnbi7RfXindY9BoTfC8AI9LJl+xdmur8LHf1Y9IP+eegsKrnOUNEUH
OFLgTzAYGsGIMCyWvI0yiYO1OfG+qi4nSZcjKcCry8dRWn5JJDUhq5WGswu5Td9cO5NfjNsZ9uE5
Y5V8ZTCR5dKwJWc0GfX5Kgif9+6ndFiC50hVr2hDAwcljT+P41AxoWED47otOL6P7njk4/jaFhD2
rRIN8WhB6wnt8Kz9d2jeH9tIu0D1iWgL3cxARr6i6myB1j3LJEctHfJI6S0m08lqXbiUqMYQ+N8/
Esxjdh37R/I1MSj4QRXoseKkqR54lgtpBYJYahZgkcu7RteYt3sW+Os8pk4Lpn73+o80UUxaofhe
e489SNbELfyxzhalACWNrFiIZQMhVLbQS22xX1jQQcG4sOEd76VSiBoad0P0k5RcnvDZejnpS3+O
Uztq5jL27KxS4x8SGmiv+I3Ah5UZ/SNDqNtPgUE95WdKWW5Y9d0POeKPmRe//DwQDcxDGYS3Eb+Q
JOov9mQY7gioU1C/Jz/qz6zJzN/qiA9ejDldMUNyYKEfY4NiQ3vbVZWk+anQRoiv2Mw+e2SPuDl2
u3gm6vACd8lPrXD6Juj6ozTWItUrs5Lis2PwoSBIJQncyJR4t5J0pvAJpdaf00ECISXubZUlALUI
dKQbN91kx5p1kp2Dv4/AYuwPXi6SnOmwyQcE0ppPM2uqsS3yShVqrI0gkd9GabKfhnj4MydBKSsd
P7hf8wP9PgNTSRxtdL5QI1+fLjqA7gknmAM8wUnsfFAnz4rmUlLkpn4ikC7vxU3rnbSt0WaUWcRl
L/yY7DxIl0p4Vyftk87wGfuw5E+7XTRTpOVhUktvUS7Mx/0PrbeVgBr+U9Bi60//agz91+dCfrn6
drDQ9aS0hwU6KqWDaAAZFbh6kfacUF1x2gprqDOws3PAYWFwjTPoPv7b0yTf2ig2lJfuKku972ad
OEAWs7nsocR4NgUjF9JcICA4JYjijnASuGIQKSN082YBRHZyCrfzuVUhXbu2iYzOocIPeOwvPCXl
Y79Lmo8ieb614IuUqK3xlkPmiOFz+PI14v+9Hcfd6X4PPnq6VXYguDQv4+Y3NDpPmvvqzJTHEWwi
eC2LmZC1myLfSzTytUnvTku2DBcXbR+ikeQCWPOGhjx4n8pbrQl0UZcSjmBuJ2ipbydhcHuVNrQ1
WBjAdcZI1+WRGTdqllfDin3rsh33LfYfvtUiXU33wxs468SZ0woIS/YcgNEZGXj+rrcul5WL4ecY
58vQ+1Ch8qm/7RVwrZj5lZbYImsnJSEG3247x0KXabK3ax2q4QOJZjciiru7HnT7/ED4rLFuqvp+
Jo0ypy3yUaP8+RhEF6VnOoauydmS4Y0FM5WsLtsLdSoYJYCrdtwLqDgtNQlYI3QCqgbhC4ywIpJ2
KOdtfEhKjuZa66elzeXZA5X5mYhOSH4zOdKTa3b0crayen05uZ+ba1yLIqqX+vIpnBtT5abpBFwv
7u3ObXmcQ70b757+wveAlbR5wJIxgE2sBTWnmZjNB7TfKijiLbApnK6Vr2htPJk9sQzEtqHO/hzU
slvP0cWgV53W6tC8NbqOOTX6wufp17HT2I49A1+7aXX+atEuqy7xUmBYryn+SjS2HlpoBbpYG3a9
arVLpDejNp2P6RrWaDBuw/H/MEAG11D/zu+Ie65nEQ5+BtRa5k4h7o34VuYAur58xKGx5BJV1ecO
t9I0xqd0UKhpl+aBHnDSZjUo16tiWkZ2U+W/8qypv7WUd6Tn3CxXMN2x09NtnKEgStH8BIbWM/f0
cFZyJyzYib43LcZqPYVmzaVSMxnq3T7OPz+zXrbFxzdojMgB6wMnoWEAW7aWRRAfnPpHZLb4sdKq
yd6amyPkZoM+SmhWEeVjmGb4k0MqLqy0/gRsk52N6zz5G9agk+XzN42NWNJcRx2BLExEnn5LDVWS
OznOeSeea6T9K+amvCylSsIhVLH/VBuBlXibTLtbKPP9oip4gN5WizId2EjtYfvKahX0R5Sla2ln
TMQki+DR989vNWFbmDkAxyuuvonPSUmTrOzynPzojFjFNNx/0wCPsXGbTzdIWT22XIMpKdns9zib
opg/RrloJXBAXqVFFuyU4RwrfFUkFJDkXk9Ak+U8vi1ner4qkQ9shGVIAHT6TLCn3T68tWhOIiCk
5UrSNcZ3xuyPlNb20U0cqfa6IUjZ35z92rS5/Un4yLb3i24XEwc8ukLJf4Am0td7LZUsa1BDZIp4
rd0pUSOHKooGblDokBQXvYdPkMC0BXk2LwleQexQByUDF8Z6EiMKrL1CquZwNU3Vx4QsXnbNqEUh
MwKFOFH2uaPpSjknbrMfWARKX4IU7C1xPowXDYzh4klStrDCSK+0Wd8/mX9OxoUj8ociJjFza8qD
NjExW4NwT8Yjd3MRZqwsBQA26/ubCsEe8LKRR2e0ezHW7jd0+ODjN0kD+QA6Kk9knh0t2H6sRrPD
hoig+BEviVd15ZZefKAhVZTK28YpW6Gw+aLeV38J3NKFRRKwwekAEQLZRxh0cWLVZSFHB2frhKxH
QvhgcyvVisnRPVz3GR+trIyAVKbpbNpJfzYt4LUKskLlnFjaCwk0aIQhpfUQjGYSIge6jxtB63YD
Pn/upYCdpIEeOQmIe6dUhQMASQotSVl73VjMoUUPwGjMYipKpGyvKBgSYQdj3/w9bjezPkbIKi2M
W+/oe7cjzgxpWEh38TVDOB0GafFaZeLxa000ZoCUys+Eu9G+aGWpFyIg7Y3kLNQkYYBfgNAoDtHa
Y0X5Njb20X9H5dhZPP1zu/hRi6Dkm4S++Jh5W3lMKts5d9eNaw138RU6qUF0I7OEFz8zvcRatgyJ
SNh61LBR1qX5A63JzUeVVqFWb/kTiTcW9wO4Iai0ZwHEdPK4tCr7zO3kvCm4sGqk+4kmXD1elbO9
I2wFgtZFkF95kvXg0AeGM8l6AjgYvP4r/FjdbKqJiWks50qUT5E0ftBg91sFyYBpkV9mDwsY4Hmz
qGDS2X1gWdDYu9ksSQKaGcTAiRkwcIFlviWwHiDHGV7Lp1UXSQv/yIqtuf5x37AKcfmiYC8DseBP
Bo8loZnVRMeX2wzlJRkRhNyEOw1ouJS2L4IbzGuY8ZZIGeihLrFTQarjWGkROk1zO+xATVI+LXQ6
X2dmAlRH3f003aYuFb75+gGWqKrMBSjUC7hbXZ2a2JkgSkkGRQyO2OQ6n8KUnhqHjpxgWMjpFHXj
GA4DHlFUfy4pCTu1/tomZvW0WVY1LRDMCaJCS3jDZjF8AMtB2d0PvruurXZlG5nzQUPo5EFCJqvC
g5vjAVrXv/dptYCMO7rSG+72JKBhrVV1qvZZGrdofWemoHyQTPMi8G6F33KJYT4G85Y+4jWlK/yA
rkvov9oDkVfCjfTaOzXVgE6B8iPHTKdxiThN5pbvZFykImP1NhrNJXiNeG3sqJSUCDbswy9p7MXa
vABoA4X/qbMTtMbDxirstUy3JUMgT6OSv1WRkzvo7j9PmShvmLPJRhgrRjMKq74Uk3dtG+t2Qe+s
UtB7HCXCZHw0NOzLezakoFR5jRuQNzJe1lnwzwZZCQcIQUgcWWIzBC5skQ7kLP9PqhUcSpMD2f/O
LDqXeKynOqOtz98BZnRAj9uUBz1edSPbyNT8zO0oKH2tykPHGYBaXBQoR+nnNTgfuE7ima9eUfDL
91/ZBvAdXEbt8hO6caAhLBkdg5G+SUBJ6v69CtOSI8rereOkTY0qUveJiNep0SHgyBKePlyzl+s+
RqM6kyJ9o5ZEI62UVdhQp5c7z/RAUXxpR7pNMjegebkRpzgxXNvZ7+n/T6sQRO3M2groxyx2EAZc
uMM8XsusVq0dpK1XVZqEtcBw1p6MCV7fGshnbBOcS734bYzAWuQlt85puczDkjjAA+9HMsKVLW6T
5ehzi850mM5Tt2re3LmsZUktHMS75V+RdiotGvVC020+stiURJBc4CgymaJ796+68hvxIRaNE2GU
ZSaCsJeZoExKF3RhE4htkT3hDVpWivq/GKVqJtR5iuksAUF8dxo0OSIuSQz2uzMKl7dj/oMev5HE
irMOqhGU+UtDd8qUPE30ZSqCVP++eI2aZ2OZfkmVKSxgFETElVsM4Z8bcvSWpeKEsyeCW5x52oHT
cDtf3xxC5p8E+c4XGlQaCxrTYTqm7PFoEWE/CVbaSN3beDZ82gLBKw45os5jb6yDTuAyScC2HGj+
PFE+Lq+S4nvMD18T3UW5AHUJVMZPGJnE0GbgXF+OKjUt5uQ05RykqwEOiZC39lYS7wC+gXClF6ln
u0Twmj4tdSPCzd/NdxFPj8zQl7Gct600M7HfoWE844ms7cIS/wgOhWrJuDFJIyRs+ukm6GcoJdtR
Djuyu15Tp6w0qC1UlP1nKZjsRxBb8C69QEKpDLvnkktbcr4EHJ1QmDISo0rKbO4Y02XErzjTp0zB
80ocS9B+tVN2PQRW52Eew1INWCw/iO3mzHxRg8BxUKjD5OBZDV5ggrEAzDW+/eve2kNdwWl+CV1d
qvKSuLPjxeMV0QxW2oasU9eCapm4YnFu8FxhEDfKNI4MuIGHY4s0zpmUgZrn36DRhRAasuoiXIaf
WHguqwIxtsWF+Pm2eGCnJthPPig+Y6Y5bT4YUM08j4nsMz72F+4vtNDJefhvnQZy7qfm8WkJf/gj
/Rv2VRlOGxHmvwvVZvqAU2e6knUQBhLbCS7E/3PaQUpNqj+CQkm5EGmp1J4T94METZ0NKa/9H0gd
Uyx8PJzCE+jI4SRhKQmG7YsYs23SEqzrxos6sJ2KaWLr8s1TemoLa4f7aXfHL3zEPr0YODg3mFP7
cw4h8kV1f5ip9j36bwsbGkqCvwhYcZGuBErbT6w70flL+hFRPjnj0+v8ZtqmNaIYJuvLwWqLBv0w
ZHk48hNl50hY5PeqIl4FExi0O3sx9FtBdGSkzzmDmo6cQAVKuyLBG0p0jLR14rMyiH5RgbdbhBSi
nYivoVgyYIAFIgtVOXIkyQP4/e8+qxXfpDgKTbL1Cux7teFYc+H8gKbFn7keMGtcTqnZ2C8vQefM
eRWK+GoG9llRtx6V7X2EUjVuHCUUoSCZlHTrcvmfsf3ZJ5ZLsEynDHtLkx0S/hoGwONRpq8JummR
rnOd4/X2DOVgJ8iMponV/URwuw6TZbDmfUJhxYSTrKwq5V4F+skk41dJhaLal7dsHdYq/4CYa+yt
Qg20R4QL79kS4i+/V9V/ui3Z1+7IUvsHnutQS8Y1g5gYMiucrNssPYr+y4yBmVz4W/+i0A1afAvY
5rhu5ue2m3PZ8ybSPnndf2j/UTaWce5rd59dcb3vfoKixyd8q2a3BbFJ2U4LaYQxbeG8CAjL4A0s
Op0hxWNgovw+WLVOQA42da61yS8unG7zIKxI9stzqXbCZFH07IJ0FJWoWqIZLgq4wegOFpph8yk2
+cit+ClDK2jSxsrpqnwIyyna8nhBwtXzVzOVS4RUf5D0jkGUCW+x1qiWJmtX3VUV0CsLVX/jmBGX
moUqjyUVSNPzLXTRUCU75rsySkjr/4jOOD2lt6Z2gFvlqbMnjXkbwhjE5il/QHE0OSBNeMf/rkHI
uMIVbgSxiaM7k12nt2Kl31dTRMDnrn77EIAr7eZ54FO+LY6Wg3QWLcCfBBFa4OkPwA3OFNPm/ou5
ihMy70srdIE0+85XCScLTqoywUTohbPieVQo4jCH3+SoE45oJnei0+rlx/DkOHrTMDqwLJeCeq+z
2jGbPpqZS0urU1WZEvSX8CiFTi20bfiXrhU6yZMda5zytD6DKHkZ0JHWWgWIGzJYWshOhp21WUIB
ectx9ujYLCsAgXkOR6/Cj3rLi2QICsFdFmv8zyG0JtHSuYNrnLwKhyLZK0LmEUBENeXB1Jy/SMqp
Jr99EUV8+o6kKwD+/lx/y+g6zm5zPRHAkDOKtCv8f/O86XN8Q4x8Zs+g9snaq2zJXSzIxCiiHa2y
e36Y+I6P1TcCu3Hh5TQ8bIhYL6pRVCBbYeQcw/S3IdTB//tK3BjTYSsP/BYw63nZVt06gLYB8G44
opyqC7lqaynT2CVAW735OqDq46WbxDU9FjFnGKqq1vjIMsi6WPhTOHpu7j///hpArjpw/OOmA977
E2JotpOL64FgIR8tb4aH+V2447uzuouQ/9dSwBrvAoUrdSXn5D0zBj1qjyHTKmZQlGbC9nAO/elO
ReM5Mm9mXLgLsBKWID/+lq/iV3nwfS3hygd0CL1exKrSnvDhU1igrz9TswxRPnMhd3xq/Pz4V95V
sQGrNQwmoPHXc0RrmV6fhuWfVhkSj6YRfWOIyjTlgnVZHdk3HvHbyPujPGrelo6+CtDijNyr0moa
oy6BrHLuTNTIF2rjmM9G10r+ZY1mDFKI6mJ8I7eG8XaIlSZOK0lzeHpexVP+5iK6Nvw8F6vrShL0
/lCPwkQ5cD9ua/UxXoLY64j2Kp6hnopEQQbxaKs3FLkFiXwnsArPOh55cX+Aawe1dNi8jf1p0f4h
6sHC6uB6wZAhWHQmIn8KR2Oy908/8uqiX3w4PcSq14jZBE3kPzoJyYiz5MlXPjUASqwRTRFm34/7
7umvfGAsNSjVySrBuI/ozKJqhI2YtsvxU40t5bmGfOhyL1aYXj8Nz5i0YHLEdRnZwHchosEm8rOr
y/BrIGsZA2DOXaKbr/NZTeVCWqeGPJMoept125uiqSjIBlyCFCPo5fxP3dQrnlLHmdfccHxZMLvX
f1P4desVN1PYAmOnlboh4+nNBpozrglNgsBw58iDwp64B62MThh8YFBnMUSxQKcp6VmhkRbuCWKD
70KLJmGU8XqRPYS0OKDKKOs2oF2wl8SGxEs09tqFVUr1bakIpzXMaU2ARW/cUX3sJg28/0lM9Ice
NfEamZr8Eh9ydxHMp+SuiHJEOTP3Jo/GGt5J+HUSyUM72m84hRmofLqEF6d0XTNJHJzm/aMqy1lC
OTjluJv99/HgNVsX//JadnDeGojAxONiqGhZcWO34hc7n+EBfq5pj3rGsuhuuAGxiJLXdp5geKf4
4gHxB8ZMfXW33sCvDqdtkFmlxj+JKMxx61vK8qpZbER6e9/byHjvs29iHv/wi5s8SSDGNkeggBdv
wy6qfAjjozqhFXWo33CsvznIpWOOedzCtdfyiWuL9nMW3pskhA9URVWuTeb7qgRVNeUPH8mBpHra
I2sSI79YvbQdPI5ILYlaWa8zxsttX6p/O/BWefgt29G1yl/KgAPzqpLuiYemaRRSHZptMp6sqgFb
/Sn9Gh9aZ7NjbUfRm7dC7KGfqIO4x+KehTNw0pzyXzBdLjmVuRwJhMoCSeWAp05doWLkOE1Id/r3
GFNaDzg6V598aQ3QhpjDYmjMfC6/zbgH7OIZkEmWP99g2T/nnluZXg9WGCCtzYzJYGQFyMdYEP7E
Ihil5fa6Iz19G09z0DS5uVj/VLRyMwHmWFH8ZjgxU6diFTiHUr3uUM5D5/M5XN/Km1BDoJbRcQKS
K+scjSTuh5M7iKFdo6FPeGUvuIj6mUwhUp3y8vUwyUuKRaUHBOlXoUYaN5+gJ+eOAFdJjtr5xUWN
H6s/YxnbrBrb/uxAakfMJOBBHARNArcpZPmv6CZ837KxWnwcWMFziq9kiO66JB+qHYM9iYFUyPUp
tZTPqZforyF4D0jvqIMwOkBjeo3FDnHw5eGnjNnHfgLVmxqxSy9bA7Spd30nZDsuboANsJRQ/xbl
L//OOVd22/OGQV3I5j42g/QC0o2N6CyRzcNSmr6V0N8uA1UbyLvp4yHK99fZyV04K/PNlF6zmvnI
ZLxzLLGz0BRUbERNjP/Pp92M8g2Ay+4Gr2pVMtpTmG8X+qq5Zg0c/5SRtXMHpY1Q9k7hZX57ycyA
kKbmMmnSUvIWfsdafiXv9R9BsHHJYUknlykIBfDBdrxx7K23diGg36bPWHWUJGNyy/tG0WQa+f8P
WXYgkjlLKcXN2XmcTbc0uGemjekQ51r1KQDY5h/FSBPcTs/4BxaMAJ/23GAmh6tJfuHT3KkCNiD6
MB6TKJBgFiYZ00n+LP+mlKz/LxaakaYSJ3jbWxfkXF1/6xya2tCg4Poukm4yRRGGagn04PktU6G5
BJD/gO9HTFdTR7il4bZarxq9FPkV4IBSMicyTOv/apnHZYax9H4ChvrL5s9kzDaMtJzydXs8E3TP
DVxwdr/2o8FSjTiRjVRCXhkWEZIo5/3FCVcX0YFoNMkQM7EfKmB7NAqCSk6JHcFuXg0zz94/ysRg
zowe9cEPRnTcC2qSubhhhNoHfoqrz01c4g+ECCTyNdfXGuf2rIw9gI0XnGZ03lDFo1TVEl6qqLRl
9T2EDjVbDlvjd4KzhO5N4YRpAP6opFK4Ehkda8rxm5c+MCnP87TEfxbAM02WteGZGskMD5wv0lks
L9jmfd8eeiY8SkyerfrMPdiCwhU1KUcI4acrk/um3aYdQ4Z1OGuVounbY5BTXFjGX5D0psb1PANg
+D/ZVXoziP9MCWRUEFSgwnY/+FOjqLTK/erFXMRYkTt1A1jbQ1IMspu7dJy63WB6OGFxPATKoVgI
tnrU0COpCvAufYVKpK0/565n1ZxGKIE8UtzXyZ6Qq81V0wQA6bXGg7xSZNhAXBqwQnSjdzpGP7Vl
v5FIaISQS/dWDnXpfEH/lvPMu6PiifEDsyO4qZojdUUTeS1JvY5PugrXRp5nAv2A9VZqGt12UMuc
c7X/5fszcHzD3RZO+IgnWl+4kLgxjqd5GBmFmM+OfgLUKYIVnAxcEjikyYfHDPyTiNlub/lAcIzO
IzwG/J7DtegMHMgwle2MtDptHh1kVGQWFxmv8PfzytQhvPCVTbxvl816D62dkeQpvNP0Kox0F5Ky
6rdGeqWC8hwuu6evHDPy1tl98zd2cnjl4gpXQWh+BxH6cQHOS2Hs/1kCIjVz+RVGrVFC7kG1rGLN
PWmAvoJZzDVIIlMgNvWyIHNE5Mea6SSd4bb4Cl4ZLhvu1vGMc2vKEPIioorrdQQYIPlMzFgcK6XD
WPXCAy7ofnYG6cVaeWpISL/cxBQ2ppTyGp73Y5+fND0rmss/TTQ3Q/MjPpilIfjZ2PloR8CaFRLU
WRvLT9ZxzUPr2p3/dLG4f71qLY3b/k/nczgnZNjPIBeCxA7cXGqFuBI30CCTWnD92EWnT+ijfHFf
MIMLQ4HRyavmKlpglF18pnKi8Gnrh37PrK5jyaK1X0ubibiK9uLqom8Ok9FHvELcijNUrdAx8wFJ
g3CDMzIcZQoLX2+krTG48Y9bhMfTWCCJFOa3GI5oyo3zXdJabvpQyaiGO707GZ7kL4INPq79FM1W
4TS58Vsh1LVFovxX6WlQkmNBMY4EDvtlbxM78xfstFB7aFX3i4YfReYPNhCIuvwYIQeuLowS9NzL
XBdtPenK74KLifBN7QSA3fdtAvNcjn9BDghVCc0Q3folRd3taqr+mUCuWxSREQTbPoFvCJr58TST
vKhItmFPdY2EJIIKq+PXTy8PmI9WY+1lzlvGvMApABjIa6iVXO1odQYs3lfieayFedRxv9pZbPRs
gNb5aHvLMkc1o9iPaQYQiFuhu311uke/pz31/dh4Z+QUlgeIczyd3bqOy+TuCf0VbguoIjHKfHR9
KtfiNAvxDl0U9MSSnp5tOlXz/UDNByr0s3ysfXBe3Qhu1Y/51NQokCUMtq518qSCUOZUn9Ef+yba
qSS+cvcABbCwBiylEUpQVCO4/K6IQBKvQQJHYCyXrEVjqTQOgxQFgoTeUbhJyQB+hjzDnVs+ulDa
ybtq0pGNvB+CX6YcflLNi+xnCl7V23TUVIP7HlwkTdtTs8y/ZLGIy+9gfjNzJp+uj7R6/VmjzF9K
v+FRlemWOCivZuMRt6uDdR39LobHYmVOUQ34aLNeDuSSFLkfM69L2hVIkjP+1ajLn5XKJOPb1QXL
1qWKp08zHJgNY8kgbB3ZdUgpDhlBJtphZW5SDzTDS77ED1zPsSSXp92zHnwgd1XCnCWZjaI9j1Uy
zjndOaKu7pJnZkGKPs/KjbN8Vy0eCp7KP+lteTX/NiX4cYj0V+rU5f/KFPSnYM35UeQ6X7fwYnrj
gf9UkcDGp64jrNhR1ngFUSgmirHvy3T/y4xpRI8n55DwaVM85iCBATLQP9Gv7Pl5NZOb6hJ+/9nM
UDCnzTIaECDfDeanLObvkzGRSsp6I62wmKrQLJHa/01vXygBveiHTogd6PsoQXwma8SyO0BGFNXG
qSyZtR5+evhTw2yCn4PE+gGZNgmiZOShAo0Owqxz3ydEPg7o/IsxPHLLu7xqpfz9Pzfxg1Wx2x9Q
xeGKdLZ0aAKhIcClO+ymWRCOgOPqzTn5JyhphDDF32xv1UWujckQERlKRdfLUgX8zZRpxjWTa/Fw
21ZFBbNmFuvFxBPhiSr4yGaTWvgmNCjcniyNrZLKMzNtQXDiey1SqOVWHMWvp8YTWkuc/930hpg1
PMkrV4ICoDB9F0tk5c4Hcsb/I0fLBPUOApsYEoOL/16S1gXS99lEVxVBEMNz1LjsAP9Sj/i2x5ow
S3J8wsRS6e34PqVmooCN7bne+PAO7KFfVeulspIYvK7HbKHUYyDBoxbYT85C99H7T/FQ4Wt7CQuK
W73ZFM+TvEk0webGcoKJ/31HWAaikUkTNnQ4ACiNAXVgGIzm6iBa5fV1k3JwceF1UUFo/7hxu9Wd
cdY1G6dDcy2ilg1wpK8/9MTks8l2ZyE+DIPr5O8v+WBm03Hfyw/lFzpVdKQIpmdJT1OhvtiVX55c
6Bp/PpglXZxKirIJvCMETtjUBeZ0DsK6gsEmtN/oXwdL/loc528BvpUCSMz/cTwZVLLRdcwhnSZ4
P5NDjmTsguhlFDsatxQVzXItyh1DzSZ/ICIn3BgGyZckce1OL6w6yqxDlY0QOTxvl0uDt53jEWxW
TE655GuvH1s80KGjVBzWlcgGk6BIdTz6tNyz6ecC6Bn73wvG4Rmzd1VUWej8Ohy+NiU4sb9eriyI
xSC4PSKl0q7doZbSXwASp8TYuYO8Vz9M1FOT3D9QRdI8NZDLTCIT0gY4r4BfNqiB8czx4cMlGRA9
JERZNJ8ba5Y1MQb14rqIyBhkCM1WYsWmSbvFiUewlJnYH8v/3TrmtptRYFnSrekeYzrH5xh+ReSt
2zwrDb1VFZXCPJL+G+5Z/fBbm8rVEsYQOB+GcOGT3uqf+F+1IjBbCmJpXLkYEjTyqI6m1iQgzJvz
Q3Qas4XJOvh1zk6rLe40OiNoQuekUkRJ/pFDtyxllDfWEFNw2+HMJIh8qSxIO788CNdjJ+YJQ3/M
VOl4ffqtdd26pTUANKNUQfSN2go6sLaig6GfBNwAeSXoPZKz4Peu7yf7ejzrVgwWAORuJ7SKr/5+
7MO8QIloslmd8dBA6LNKJEUiVekqlGVXcbbZLGDcSdM5ASl1Lz/rnHTrDqu4LPAfDTURBGUNTYJS
8Wj7P5USjwq5M5BCZYB4IAxAWjz07H0tR/vnaqd8HhKECNxLpZdLUm9Qnl9Jkgnl5GnIWjQxFFDb
axm1INLjXrwXrzpcIO4rz83ACiN9cOYe37V5gLJMyBimiyR8l+gtlgmVkVeETFwWrjmBGXFFDitj
dxtCEDiTMJ8O8i7haYK2mdbDls9JHVRJKfQovaMXYyD8gEtQ91BIl6noL5yc2mIVL7ZcIexyvb39
viZpjxVj7K8eS7kkRIbZm5O+5GtFGn5BRIxKm1czrCqCvMqZg6wzyAlMGJj5KNyaXlzRJPxZbC8c
KR7WCkubl++27vC5C6IaOyxrUHj+Xnl7yXGyV7Cj2Rxh95OEjFknz/t59eu2ojnd0HaJIKh1pYW/
Y4M1ahRqXdDp3SnesChX1HIa5JJA2OQ8xhTz9F03CgzCRz6pmqLOB8go0Y9gxPHuDbvFaQ41BJB6
akTFEg6XQzcUBxKL6ab//2dN80mfY0y1vVJpQAHa4iC46CIiJslX05Y4xfZPAC6BiR+96BT2tvA+
MgGQh8wIjcHnNUyuZADI5IJqo00rQxbo3LQaf9+v3j2aGu2WdmEEPC2SFEo8SnnMOtP7YyHiWyXt
ONycM/FnTW59DhkCJVHoDKQIN6xhwBQG8d2jL/aZkITc+DWlrFmHI1RCOQORffAovHuFS+40vJHh
XTF/OjknSPZETX1u8agGnIHVb3DeRxYgzEgdktGM8c1MB1CLzJCiXNB6Am4wfujhcD9g6BMvE+tk
gGwxK0NZDddkztH7JHFkkd/iR44rN+pk8bxuAARx+tflqubJCxsbdrIe4sqhWrxKwAYi0GYH9UUO
mylpme4OIA5lPIoO7SuCsqM+/j3Z3hS0zRU3lUTTRZ2zdu3FbwobcTKjtSZUqGX82C6ppsTdwTkN
ciQmn+7dMVxQ7fMN5nEkbJ8HqgjO0FF5ooEJ7m6ESuy1CmI/pJUv3o/Ag+6KWaTXM6Ot9l2/8AOn
MwIaP9gwlDtN7NwD4iwpDGKA4lB3uTUKvJ6TI1VLXAyufRf+DdKiMKD9a9BXtaGx6RHpTuKQQbuD
+Auqu2/FYZMJ/z4/LHv6UC+rEK499idsBnV1vjowc3oFAL2+NTYpB/yccyQccRWN75K9klRjajpT
D9Xysa6CX0O/Me+jNO0KD8cZJGNlaM+IqMiQyKYpQTEnpUf3LQixUgT3QQjluRl+TxBhoM3blLWL
qm6jwmr/WneRcleQzZdfhELadHkMZWVXMAQS0C4duVM553BDU6x3BS06by/BlWp71Kf15OdEOhZp
pDGyicfMtoJeNtt7erkLqZ/AdD8ODgvXZ2aOqYhkckQ377VEvbQGQ/Q+HoNOwUT/cVQezW/c3sjv
3PoE6J2ISlAprmRk+MdUmlkmSriBR+6L8Dlp7hOxj3Jr2hrnyoJOxcgKVifc2aExzJ+gN/ODNv4U
SA4AVNOclCv7lxkfQ3DfC67NrRuQ7KEYYoyDQ/eA+vgeKsb4RnTKePUdXkJFZ/O6kKswj99J86y9
71ZbLy9FF5mVbDGPcW5bZ9qYEnv0P4HyJGlUkND+/aKEbbMteY14XM69qgeOoa9Sp520I1Nje6GL
DUOeZ1RFCG8wg/Mvflf57ApQ+oDquOPl9KorzKNiUZWUGia6WFmhMTmqPXgOqtsCKSs0FUh6WcFO
ZwPQRggSd4Ym/Wr7M2N07vCxbEkkgujlepIHrOF2HLNbM8S5ORu4ACSPMeY6NtvU68fsyUJNL9Rq
lyvmPo739nimbqSK4vB4hZEkbV96YoPzvFkie5tP2l9gYY8UPKSOfYIfS/OSi16wcV06KxqvSvzl
baa9lZOOz2rakcPGFMKLFdlTprZVCnWBDOuLnpZ2x/j9ME2n3aNlj/cuiRdXtx5M1k1xiCXN5d7u
zEA/WuEit876/rHX06u1a3NmL5hOnZynia04dNKARJV4WiJnBGecaIMlLj50ryIuJa2ozPJnMP2y
nk2ftQ37oJiXex1Lt7780pS+/GR01n/d8UdcUS8h7GttqC+R5ktjx87NTK9scvSErs/3B14dw7RF
asQ0acsFUbxwX4AP5LB+p/043q1g/rOH6/pqfpBeU7PZsRQEn82f0FoY1q5/vGISyARpJeoeCS9g
XXRvt2Ipu1Zdd0OTRanpnP6Sf2D12uBBJVsrSB7U2h1U4+NPiHKxIUJ7YqRIm924ca30EIuYgxQS
Fccaf8/Q1xywxDSp531KhI2R/GVawhjNtrCowBXdUfuSH9YsfYGrIER1IETmjm/Nxb2vexDqWaTD
fT20fYjSN4AgHWhP5SPrK3THWvV2u5VbsRzKlqjuy0cD1V93HqghNWf4YDLCIEnDX8HYnLXEmH2j
h56sDpPE4pHrsq8jyZPuUXZzMOIqGNzcKRRAnf0wdPEuuH/E0FPg2F3uWy1mIarvIPbFscPcYfK9
YN4KPpUHv1zX5eL87v8XhM+uQ0Yp9s6cheq6af/j6HHhsZ6xkVDIrwD9s6nrHnB3PBDzAsPZ+9kE
APsNq7zhe/aSa0ovDvUNvTf4W7OSG3rDxBdHuhTw8IAILspX8ykF2Fdp9hibLsTyq4P783tqep6C
C3liugkhiWtTx1KXn9/9Svdh6N7s1LmEj+LKAtO94OuGcV22qGSeKUM3kAfmFVpDTo93VPlxWXzP
87ih1x/JfschHRmGGAKSrD8ja0zUZ+rwChrvo7uhwPLGu2gknojuLSyiG3mr2NCkfHkJGMSf5ulo
/qNrCMl/pYepJYax8RIeAS/ROZcKFQYdsH+bLULNE9M4ztwF0SPXJe6tvAJ3gQT1CMqviw+Kon1W
eSBbFvZ1KcEVeCmc2jxkSNanhY87w4Yeji1i++TArzyIqDUpK4ob+/CNLCxDEwyzPt9nkh4imysY
dRs0e6YR7mWuIF/z12ZUihUsNNddXNXyMA92DsYnsv2u04VX2seh6Z5163HDy2nqr+kwsOd8631F
g7jn1yhUloeoJVSWj8ku8EwQ6YhH2V29Zmoy+TeVcyRRWKKeQYphGTKY6ch6kmb1GQaX5P9EsSJS
whIRmPebXijg/1iUe3MBzYjrbzcdBTW7qppWypAb5Ve4Ae9YMU3aMj5AvhapW4Co4JRziKvXu5bJ
7MgQnUkSx3f0EemVMpMdM59tvNAbqrzCCamXUJhs+T0ybXM/UbjHoB6dtAfQsQclE6aKeqw1cVA4
O3b3ZWYfdTq8jjTFBalo17/FxBvI2KK8saKCCzUn/yUwioOXniVHbRKYi10+hPWkdXe6FsSW1o12
ybXQvMhBO9O28IrBLUFIIbv7JucRxdDZ59BMSx8O/AINKU53tp0Uyi8KMTEv/5IiHVIH0ItrPqfG
SRqT7j0QCH7LeqGNYcgTi358V9Lop/RKukOy9yHUul8OAM3Q47mmIGfDTp4PGYbMn+ggmdwEKhRx
5jLhKsb6Mdtn/B6jKR3skllW1jq4tKMpaHeF4Vz1pFOpGSAvj9WL0qTfTJ6MkrXsnFR1WQZsER1v
PN0+SkazPe133GD6c6yKec5t5TltFc4BlRD+iKtDVzMJqehSkSmAktGMbiHN136/bkVznplS4C3z
RZsabOOKZjWpPW0KTSS8Kp7s91hRirf3sxWQRTJRiHnBL6pOnhVRsPZERgv3Yh1i9vh2g50V11dJ
DbpVkCleTnAjghfw0mnC/pN1wJwZ9tTTfRbJGbZjnh8b/qXXUPD+Gd0m6iNavG1vUqlWulkV4x6e
/D8Iz8M134eNQ0sLgs2f0O26bjPlVwoMk/fIWEAisIOM8pyb5UByb8EOVH+QdzWDyW9yfhHAukp3
7IbFhQgDrGatHPIHCqfNtslTLSV9de/oO6y/XCD3Y6dvprVYe14OuUwd5x2rfJfcsZVnIp7YqaqF
eGjp3Im7Saoi105lh7n4WkFA9eTXRZkEnE7hJ9dRWTq3vqygH65E9uqDGyPY9npNbtBuMgxA++En
SBQZhPhIVrij5Co1KD/phZzYb6DTGLnHMN99feut3E3ViO8IGUewv8n/pvIQO0oMfh+urPJjKrch
j/BAFIqnaisXBI0uKgwtb6PgcdeepNPOP3nGxP0aD9FPJRnoszrzq1SY0CUPiVTCQ+c7hAJjo8NE
jJPlLjVKibgr2FhlmCh0olVO9+9chBv9HoP6aAXT2x83vLw9xcpawEn21xmSVbQ5LpCjqVvIfI/a
3mglfBgHoGabELBAdqTQzPSCCDpKOTWiAqlXJ504z0u3ECXyZrEzHdT+KGiSKH8hcZG4wPXx/SrU
CooESY3PmgCmMj3q/prRQZUKX691BY1rqah1sxBsDfTO7AsuzIgTJL39ETUjD8EOF3/tdgHQ4XP8
VIDUtIsES3dGauavdwrNeBNULx8l0lthV/VZipYOubLaPsbXMtsmPXEz0BXDNqCz7iuzykrrCYjG
GvXTCBcUehHqmQMipoL1HrWUpfSJqug/pH3X19lZl2UCZPP9xtjgAbCCQoqfUvvJuSfLx9gpQUvv
JnaF3ekOPTn7z7IU5L9f8L8MePcw5V309GG/nq+ect+GTWGLIvJaT6Lyc3WoQaLP7G/GCzEEiCt3
rvB5lPYKRnJ1VJkY617PxklgfkbAsU//YdLNxR2LhKd7wtBy9fDbP0llSdTHwwmq2jOijOUKxV8c
4zS4Z78KstmOXoJP7kk2eC4VVeZKsCPDOjvxArkt5FLVktG8OYoY72w+IxLHlyKgXJYia1U0466s
t8N19NRMjNib1RFK00bANXH91ZGRyR7u7keYM162VWbl/xnjuFuCilZBuzvrhJfvJHuny3VKSMhr
HlheYOCIKvRzpfTzZ29ghi+VJ+NxG0/RVgk4tdUT1MoFcsbcwDaNC78lNxzj3EkScTIfdu2Gj2TJ
XamLe6d6x+IhQIpsm/VHf/P0c8P56gAQNXUo0TtnLk8KnxfmVGN3qMElwziE61qobg0rYU8/UQDX
7eP1P/FciINjl7YffnT3c4IBB7l8BjPkLmahDNC68UvQg/3ei1xovXW4VypD/q+1NznmDbKztc/m
I2G1GnkZ5+BmVrWW4Ey9xyOthfKleBgVYdLfrTdBcwOYf0zaOGNvCL+RZyyFIL7orDgoyWxIvOCX
unWiUCphZErF6RPH8N7NmTH3kE0vx9s7hrEtuMs697RMO7EMCawnpm8nq4kEu2Qy1X73TeIp/DvP
VmqHmmxht/tWFoaKj+S1sC66WTLxvEwcoOrPZipBxdAUZu+cfWxRr3EuzIueY9rC+9vQ/m6J9WwK
sU13Bd2JfBkiKpPRWroICoulV1SpRt1SfuV8s3E8nkcFeshWnINyODmSz34BOd3NLtH6GHis5uwR
xVbxnXzsrcrNsXBU5ixH1RQuzfwjk//UbETX7SDpeP6ena+8iV708nl0Fn7tDazHLBm0cD2xI/3y
Qc486onYDhjC+umNBCtcezrlcnkom44yS2VIWT+hxy339jVJvc/FecKO4nf2kx8sOirkO3CjPPP2
V+d3tPxGT7rb6uFsM12t+flNAU1dYvmsipcMHPOUH+FrtcEMwHsuzYwYlMX6v+vlAQ/ZmXJopLhg
jeE9QPenV0VBR2k7Vv23+BmBjDE9IfNNW34FQAmV1FcLLm4Joy6uB3P9yTpaScIW9n3jtVXn4A6y
/lyEO0wDTPr5Vg8fakyfUx2L6s/jrKcb2Q/KME1/I4vJXTJHlwHCRb/wQdI1GB78PPL+AXz8mu7/
/42vVOHVyXoYNKTG8uSHKCfRfwin0OitozrHU3tEDxuTwZw2RzpWCeOo+YA9Jr2N158Eq4QWtFmS
84EeIoZkFKl3MfbY9jFH1RZCBQLaoVWbY/OxU32u25voMi5KAhhNJE7l6Bwnf0HYt3qEYoy2X7ye
80ZMEnY/vdJXz+yzfwbR2WLjfC1XH9ipKUma8qUl05TJ+aWE9gejnZib3iEGwUHlsoKGUua3F1CQ
O4OemP5G1K8N3Gnwu4mjeRsA7OUIO4QlvjI9vaSz48v2wAjVuEE5n32cYH3F+K2cbhg+XB7Afg6w
pwcB8oUDHLPiBQvaonZVEQqGajvWZl1diLhkPeZaS2QIf+EBlm585TdkpyqywHSPzZLoRNxbWMBQ
sBREaSIsZZiVl+Cw0kBlHz2zqXBKTH+LGk3odCvl2QgWXOm5+sE0qwW/4X6lN4xWqPGxL4hia6CU
wtlNg/Q4v0g7N/6Z0ppy97j5qBeIkfMChWG5RnRYnkG56TuvAn/P4a6vT+Gfrdcseoj6UaFbsWhM
7/6LsSGfkY9sfuTJcxj0mZ77RMiY8iTQfKOGz2Ox+i92mUHkXrEZNzDOIAVRD+mKAHk28Yt7/ZBS
6ly53I/PjnsXTyX3W2uBN34WHn2Yw87XHSo6hHopMjZAolrMc+HA3oN64Y19CEH05pYrwT3JdlEy
Zw0UuTMMX7/1nfWMM3JJlnw7wLPByqFHJVGc/GR+zVBe2G+QotMbUkRmlMlj/NyN1dL7uPA17flk
aj2WQ0Zzx/lzI4rfV6y91nxaVYhwE4uNw4wZ1DmJXmsJxl+oBu1px7zo8tTVoNzEgcFPVDDSk0MP
iF2IeZVlKVAX6jgqoycChlF3EanV1RoYpEsIrlcTsJfsEMbT48OA1QvaPrBRZNeA30kU+dJoS+2X
ybAEEli9vkDseEbLTHu1UXS/nuMdgEsL5Q5hftfQNTh2HS9nKGeKGjtFFdcbKj6DFMVuLS1eqOgr
2m0yeX6w3TUMp01+lOj+HJYaU+4BUXl9C6Wl6lFWUU74KifEaXgj8+3Z7JwwwZOL9eY2fl+FI/t9
ALvj/OEpS0mtTlarPSP5nJI3PX1SXQVBr/R66/8VSEJjI1hYTnUMOqZZ7JxLnr0ymI9vYOnmblqT
HNP3fiiI+tUORXPyfvwh1Imt3x6CaJ7o+q/wvhGhKglgfLWu1jcXDxZPtNwVvL71MjOvapwJwVal
eF4CBF8x1+GAIX44OxgnARj79Gz1YGepWDPswAjc5LPyvGdiOyKVZDElhWoQA8DwIXjjD80iL6Fy
+NLQAphYgOw6i6HVSgHkOKan1nk7O4KZAp9RLtDJIhdAbPIVV7ljJRC+45mma3tLJKBQY9/xP/KF
YYCYLuMfRJ0V7EgAcs8cmmpbGhG5eWP4a0SkOJnmXNhUwXZ2GAUeOEIOyxE3GOnUIY0JeBHBl80Y
Eg7NMnImKCQoPvwzIvK5n0BNZYvg7GAbH7C/huIO6jGLGqRZcWbGa7qMzr749s0XqjUswi55Nit+
rIt5JXUB1YfqG1m1lpyyU/bHGRLryUeybKqZmW3xSZqcmbRLFoeY9kZ6Sf0LVWMYtYUC0HC4Xl6u
XLVxXuEvqcKPEZmhAoqFlX0yZOe6G2gjDPaIMcLnvPcU1tkmVZfShDV6VU4h1Tm4clSDcOHt7Pjj
KPU9fab2EsnYPBPEcNdM+GhwKp9ikMMovtdO0zD6XeHYRTnNCKmZ4EmB/gFPVtarSm7EGGfuE962
EJ3uIt8oAUSHyZxX3eA0QL3cg2XZLGnXeZq/jgrYYhy/lv1VEwFRmJNDfLDz8b7frRru0+o9tCg0
ikC5t5cEv1WNlgaj4nR7TT5l5xH+HZf3vnQ/z8cIb0+I3eAB3ey2Ow1XLphLCrHrBk/K2F+SB9Cw
pSuYjBNp4+KsuZrU8R/lX/PGl0SZnBeRs+Wcyqkmw0VMHSX+p6eq84DZIDJOyQFHpIIhayJ5VkiV
NrBryIyM2LnBLJxmMZ1/nw54hi4tTvzpoXPfH7mpVhw2DkTbCogys0AmRhGRszCXCh58CS1HZzVf
3CERsitz9uOf4DRfaVhcSIM8BH5FJsv6Ds/bv+lw43xDLDfFzGkMxQM2/4PyE6Asw1ZIB1rEuYhv
F1sz6IX7mdg7iuSxlYpLZ7SzkPvYxpyvXGSrMlXMPnT9FVuwu3OnXsThTN5HSET8yKSXSaqeFNXA
sw3R7EHgWupkSaZ13AGaSOl1ieYi6Xnixb95oGy5g2Izpx2q21vxPA2knw5HcXtoGveG/yiFRro9
hTfxYtDns9A5swkObfTbN0D7MLuUiRYKscA/sdc5ckVlV18VtK8Cvy7prKw8VICCllg7QKGmHu7V
L4rnf/qihl2uR1MZvqaHk2ybbpalteSfUFSb6j1f9DJ4xGRgL5QbgolMnPeZTmNdAoQSB5mb91RH
mciSdXl+9HR2ZCNq1pM0qf7yKsR0kulqW+bYoy/gyfcP73/IfpHJlf0X3wfB6m4rVR2hjo+Dtsta
bul6svMJLg++XZVaW24UDGIVvlvuyysCldkRVY11rh5z0+k0btytVu0vyl/to/NUWes7TwMZStlK
ofCrrJQr10BENEM5dnEYFPanWWcsLOtqvBhhDgUN0uT0G2JBDIHkikZDEbwL9hnA/if39tKpCML5
5UyrBS32st9FEOdEGkS8X6DHOsp4pZYuEhGP8E42lro8DxelhuwoVyOAXz/fYk4BOOEwhngvRij6
8nmxyx4+fLF39zIJXxTIi1KsqLmeogFs1ISd+ClQi0K0eWN7aG28mImN4xcmzrfA2A4bzSVwv77M
XW83ZNTL2xR1qwiY/6Z44EAHYRAT3u0vBmTJ0S4v2jD60XOi+QbvuevVvI3Hmrd+2QsKFTInnRBa
yxyLI89Lz04luPwU/CRXZuORVeRS3qn3A9xNH8xuSfBWudpwu4/6iV+N7G/75PPMUqsdYkMfgGoq
JW7q2IRnKGywWco+TxmTCFEGaKnYY8WkNQ5uysimLDqz/ElYHYlNnJ5maXV2fpSo+cdzVyUqR8xb
OzeOwKDPuLhF4O92sUyG3ebJDpGKOeLUlgWvVNeMS0j/LMNn2S+jGHSBOzNBV6LEN5ceRlPKsQfM
2RiGKZgUrYOWtCnzx9jW1qISaq2snyvw1FA5ssXGruwMwY3nOANnfaVqtbmLm9lMyRSgpZR3xAxE
3FUMpPWs+7qhwq+PbJEsVXsQORY7mLdGi10g+IvoH6+fccTvZIhmX8w3Dqm8Pzx/mjtoqwjzssYW
MwcOwxUw5o1lQVB7K4maVxpip0SH47ogDlrLJaElOgMpTUaccjkl/PyOI6d101IV6qbsh9UdWS5g
ux6tOzuyK3/H47mOzQeHYm+owDmka+PDBJ8heXytDXcgDa54OD+yqmydU7A25VSSZd0VwI27Mpo6
SlZ9tWq5A07BsbsjtoyL4RLZsp2pVkquArKWX3cGAkzKJUKiHv+PIdLn+J2KD5haaiTSyP9ZKBwc
+PCD/F4gFxYhLjYAOIBo6SR8v7VzE0kVVnXoHb87L4U3s8L6doQNhclciNbYghl6fgGLx4VgWgZ3
yaOvZvMS3oFwkD8LcQfHohjHWPJmEky5qYU3pd3ZDP5VejJ1SPchBglnYaxuUDSGaIo6pWvHm1SM
FgjXUQeUFdcHf98bU2BFwaxyiw22V2PWWXja5k/DC1YfdPdJ1tEicG5XIjassCJPVSGbQbNUKlm3
jL7xVvzP7nLY5Mv6ex14xL/FkzkKwFE1N+6yEEiaOLUurN7ZQptLxPzpxS2VUrfmlE6mCNhdRjnJ
X9rcGFkxvrdY2hBnLNafpnk2uk+csBmWuLD37jk4Fga/7PjPVPifunCo48Z+fuLM+a1wKfIgUfdG
HVqeMkB4VX9co+K5+wL9Mfj8F2mhdD9N5kCxVsd07xlldUuUYN5eQXj1SQwKHCAJ16HwGbyYISjh
5RB5LBGgtAsI4HIFQVNo93JUm1RpivImYDB4pG1RL4I9xgmac06JuCDsgvkDapB7MxSPhG+qwec6
bGkUNlnz23oCeIyRwLMg4iSN1ubSQRlyeyE2Rzieqo0zx1AjOhCIfaAPNGOF+LJr4Y/bvkEdCM1g
j1/orBl7NWoSmUeNT8voGeAH5o8pqBAElUZWilGOgzx9o0AVTZJ+ZdmfMqKg967+5HzfkQbGOehC
Uiu4UuoeLODbKQGP+94yRboz+JQIoCyO2P3dgRbhQJPLhzIjqbNCOx9dNkWum0LjaGCUOgawTUoz
Bh6IiyGAjhOW9uFOiVZw7sFH6O0xG6up3MAK7wBho2OC9Vs3vbvz5ocSFLT8Ic/SlPwOVuI+CinY
fdWj0+8xWYr1Yi0xsMZb791FAXQ11ec+r/5yto/g0cTeG6JfeWegJhYf6P/LOYDW5N6ITSpLq+N9
NWszYEoO0i3vUhkTWL6iAIwtpkVNsJjB3R2rH+g4KeqUUnaF50iFOsukkucFUie3maDd/ZMwbiRL
wdq6evSo/49QJ7yWfxB1rncQqu239qI2Wjp6Z+hbLA9m4TG6tPgmo8j36dXIrjOAs73SP2AYLrr3
8qVsDOKrbVHmrZEpyGqq1jU4VDP8nNxLOZ6wtFcyDsxauM3ay+U6cgbzj02zAodFXhXNsY5fHjVL
bZNPOZnXRrG4hUWDGWNHkbnMoSbM+PdfO1jCR/+w4JmV15Y6Au5e5vYdZlj4pHdoUCrUpYC7r7ly
4QkZ3NPtBFeyjbIj3hyxWPT5kOS759e3iQ22WZgtU+qn5BdPqFuxCpM9TXwbS4cfdbuFaKhv27Bo
0jKdpbmbMDiPwc0SIx5DkFBhHlYOQbr5lJgO2P+Ye4DSfTHrQ9LWyCrWfCJW/Tt1YeP2fYo2gmkr
X5oy3PT6F13Vl++xvtrf7xgn19PBqLBfUqAYDOu+cmckf3DzhuFlc3zVkqZHczRuRAvhBRzox+6B
Tgtub2+cnaM/N6Tf+1ArpWd1O+zE/7LTeMCQljAOFZHd3vhJ9odSs71/wpaxkbLuBLt1gX9GSSYz
a09xu79lqDNyJkhXN5knHcnL53RvbqIRT8B7gdpDnMrYTZjYGEaJFMHyyx1zownPEc4/pfbDWTGm
n7lB6tELG6lIFI/z9DFymTNhQrdWFnrXB6dQ7Wey495mW4X7YPk1LZRWqtyWOLj+4bsOo30qpGFU
yrzsvhu+gVtNF0ra6uwiyjx1u6KnSv2qIdCa2j921Vu6qOjRoKrWRhbu5LlGaYYyqyXtlWLTQuVV
EIO3U1f+o7dZ7LRjhrhCzBHoWl8oLdfT0dXDBqj8m7Pax+C2YSfuTSmsR/o5VfTcLVZcFJvQpnI/
S/+ShpyK77z8ws1Ox1EFwlyVEdF5zo7jzTf//ccuQ2/XmIaO6iBey/KAhwVzkL/NRjmoo24a+Wms
3S4o31SAdQrf6/3gSq4fP8dpr76H6NGPU6GkvrVNxxhjapuanpv882DzQSUGlkbyEaWyzesJuzGX
RG3f59o9yN4+qyE82+Gq8eYOEhzM9HzfJJsUIRxFR/HKLU5XBv/acjzySQTprBw43UgyIoiRZMZY
mFredwtdDdnieeA1VqvJ9Uj9sv8jQszCf5U86qeHYw084S1GBvOs82AQYOTe4JRpmGybzuzVJJA3
TPQzteHCluvr5Se3mN7WnLdcMY+inBP4f1Skp0ZCpGLS3OHCLG2G3QcGQ63ll7LzNlijtNUxyXWt
yhutiHS8JgV6vZ9+4j97jhE/uRQTV9LUApny2ZPHTqVzo+W0ToImxYB4FXHeB+mZThmnQpR4rJ67
Jl3a3xBBtLut1WzDhYhb+ozoEkpEZt2AMDcwP+MMXEhowEmclNHA753GHctcBJDCNUUVBp7WBAkS
u+qADoYYazSzdXuawSIjNPj24qvVr54QUWeggguLfPcQgJPDqGHZJgbTXeI/LWLbbUitcFRztlX+
ksOM0inLngdQ3kvv+hoeFjKdt25HHwdUEYyZiTLIZebc9KZ2t0Q2o5P6gn26xO2slqVosx1nlG/M
kJ4ckI0S7C8D9qNjKruwoii2GtwziZGDisHh3FF6nXiPjxJrQ6o7HLG9w6gT3ogxfcTeAMDENQAH
LRZVV5PrgdHA7N/uSlbL+qFFyq+cnMAjrCCOeSL19MsGpqKV4h2oOHKLaAzx+yUEYQIjoGVyQDsu
76A5CDMDr49+FpAV1bZP/8HoF9Sc7bFwvgOb3O3hKFI3akJLhXR9Zy9D9TSg8ZA/QIWXR5yeqh4m
EyUu9gvkjIghaHuP6bwE7YeUmKQFLujuw52E8RG+o0zxouDpXLBnJ+HtA9GI2UbgQWYGkJBRDMSy
Yd1ZBIAC3tgkawTEpmxUzQDI2J9tDm8+7v2e7tIsMZ3mR8MNUsIncGVThtwsMcimErbEj3HsA28Z
8PlAgBSU4g6MBJQeFxOGjvf5Mc5JRdf4G7EZ/3miwvbA8o27HZMyTIQe6lmgOFZBRXFsotyGbM+z
kntCKJhYK/1PBAfPzRLSKtHPqMYLjHV1RIXj15uTkJQTNLBcKp+2bzP3joUGKH0zeFFhkjaxngDS
XtXEITHDkXAbCBCTGYNz/ldaNl/kSuNU9I2qJn7EDW3IF1x7Oa9x1hQq4Z7yPr9OoRUaWlC8Xt9f
Ggfp+r79xYzzXoL/TKJuXNrw2xuDFx/s4zzVcmqm7Biispc+DNkMLq8tJthBb0E/vRCpZqqtsN2c
CE+tcIybtQ6bocZgwRBQX7+HVrjDtUVNSmzOvXJJuPe47lbM/1yY4yvaOlDX7Tpfqioml2xD8y+/
q7AEQim6w+W9TFPC32MrqCIMUB303t+VSlr5arVBpU+Gt1w2X+9LIg6oVyUCXNVDou6Taj4j4lnC
SxBS4+DSD9KYjeF1Hlq2+8tywFQyv2fsEGlQoMbjynmJgY1JEGJIQNpc8O5ZnsJeViM6+nArX1qj
A/xOYcgIwUTDwtfcd3YXzU5P5NZNaoXcjPXZ9+38PZTCezkc3Ue8xeTOU12auQiJ6Jbwtg7oFqQx
Nnyy0eDmOO/xqBj/GD7JSm8QD/EJpaDrzmjwb98/7e2prEfrk0THrfhIgM8kJ+Isar/HizD5GE/Z
/ld3dvr1Wb8SgkJ+47gM2Ymg+/dXFyHBhlPtGEPL6DzhqcdngkRdnecNvRwC6Iuwf46Fihdp8PDh
xDufftPSJ/bJgSdFIAeB/8+EKZWOO6Yii7X9uW+3yjZDKErsN6s8XxSj5aoTrT9cc78uHfpw6PVI
AvUxF+VS1Eg4kmhKfv+Qk/49F41cNyM6wo3tPlrIqGex8fHJ8bfBVytrvSS0ly173SYr4H6V7oUV
2sBfr2hTwtunakdtcUEkWVqCrEfCQA4hZFPIP4nnfUmNszIZFvBdopL4tkwqNlK0744GYUjx1hu9
ferzfobLPeUGzOWBYe91fssGmL7+y9Z5tlB/f+ssiQs9uo9sSIZQiVDfwfeWAdoNYh/1BIAi/2HI
e45tOXlgg4ws+qtnRdtv7QSHtFK7pRB0+wBiWqxxTfpxtqc0RiE6dIvRnhaLJfw6VLYNJ2luZ1Qq
VCCEpKvufyJwAY9NjvmfhLyfMtybPn/igPOL+OpOaRduOumbRCn3CdS4z+TisFdskt4VVgph4vD5
YnB0GfVZ6kWfoiwUnN0oW5qGrYU4xDsdLMPYG/FkPK0z+5Vu6fkB286oXBlZJKSOX9IUgOrnAKik
Kq3POltyFWPctSTSIPFpx1KUCBmaIt8DR5m9K3oPcccro455bMAP8afluoK3IxxnZwy4VagQ1lGH
sy0alZMV+lAtxyk5I7OZ0qw/7MQfmAfbflGE2ZRbAP5RVmJ9WtlMZE+laj+C3E9yyv95yR8I8lqH
AcF13QPLQJ7r7+lAfTl3xGJ6zjWN0PNlWZzp+YP3I2T4EYzGQgTQknq4oqaYa6At826NCVFbNLGg
1CfYQxgcb58mici6weocA3IXlnqX2zjnwoiOQfh3LoA+R/2TmjVn40qmsQ4MKZBbGNIAe2mrDU7X
E53scGgtIGl1gXfbnH9RL8JNUMoGwQRjWrwV9JKa9uGYFQWa5eL3iXOnCJad4nGio9MSIJ1R7dWq
ulwPwyYGVdjvdbDKPEB7TZnxemTdeyRSd5BCFoCAqkwUrzWgWpLg9FW7sk7LWRWr0DNp2nujenuw
mXDlhcnahPUg6+/P0TOBiBd9wzpnIrFNRophQ4HtObhxSxEL/bQ42EY7DqYof5Ox3L5oZjMeNqUu
jSVbv4YL6fxn94h5cZisgCTqJ3q6zJzFnflrSA7m5b7/pXkEScYGKIz6FfAsg6gEcjZu79bCjAt1
aY0yM0MEiSIPpAiYc2cGYnHEcDzFzIZAhTusDrL5x4gpfZW1CHsVfJ1Ho/1BYtJdlL/KsEbYZSj5
lDSBCx0kEbaSMWBqpTkhGjGIJ4xYbjVznI8LBnGy72TSHRffRXrepLTpgPpmfv7+o1W3oERfvPaT
RwgQC3RYy5+WG8DwwynBnJOJzfmDfgFZ3hO7G5Y2H67Auf+/TDJqoyy2L8zvITnLNbRbJJ+pHroz
8apLl/Ux3g+Ya+V7vl9mR5/bj8izmEmpRM0rcWeMtwcDHyLgjWbCdFIlUMsBqXm7bIPG55V5tiCc
OyAUPwv/EaKHfJoD08pDxtXvqTVm/FQKB5wDfgV4UYzcXGItm+JBlYGHEAhdL607Bw++Ii39c1Ei
v88wIg9KIPkm4fWbkaHnTwvciohVHn9S1fm8m83Q5hj+C/F0NXL8OLcYlm/cWKrmdo3w2tSDZStw
2pbrU0CkiXo/Kfl+aohPIPvjSbMahBOTsEX3nieh/1nWQVUGbrudWTFXdFcbEP/4lnYtXp20TedS
B30uR2zH1+m/evI3SEKndtMpqU69/F3LE8qijWr8TGANl7Vti7UbydDnzsTv8A6gCrw3ZtRr8gxS
m3OOXcAuZ91WMAeLXc9sw7Z6zp2H02Zgp9dS1t8MJuptXbLaXvVSVSbPUvdPljJNlLg7W7xzxDZc
wOuK36p7YmVJpgHX6UxYFL3hyOckeIHhGBUK8BD1vgt7CHxTZeWYd8+3C6mqkGGFN/8ht30TAcAG
DCpaZKp20hUwVi4HJv5Mpbas/ULoLoT+r9GDnsDsX7V8dUp2hgpWiWzSlX7Vqob+YDVFO77s4M6S
kMIXqqdVCTKMZEGzsYtl9PsAZKVOFKOxDn5MjC+M4wz/wv+nyxiU/RL8WSE5LPQTwduqLw7FGUrE
tvlErGE2MP/XpPur8Bvu09OXRAJdQhxui8GYOptEhsf8WuvG7O2Y4Sn7OA2srH4TmfgdUlL2K2p2
Llsbe293IaUDYwbxsQAamKQKNxZ0Ptep+ahESSF/GjRVrEu/6O3nyERLtRo91fcCQuPZ4Z52V37e
8AZgAtn/NRy958tkv8dBs84Qyr89Z5nMl8OSQ/PLiz4wY6aaY64xSfOAdqe82SF6xlGp8dmylzli
X4zi3kh8d8wKfbpUDaSMQ/pQ6IMaFU/RrWKKjYekOaOvSP5SXM/CVX1HLwlykUwI/E+QMbPU6UGJ
2IZNxgsNEomkACxTMpenUFDPtnt1xN2mKiFWOkydYBjD5LoQL3D//fs0pvZuHesDKnxGUHJ8b+cx
sa8mYbnH2SCqSRmBIYtqCwu4E60kd4QB9BnEKCszl4C83COUCs1kqxgudN8sfUApOisjaX92E3Bj
Z44pQ5cKf3HT10kxmZ3+uOlc40+nmXLDstglMgeTa0L0R6IEG8MoGdGjzG9kRdSrU7OvQRX6Wkg2
RjBTMUiejQwCrCSrao6dbsHcUstOvBbOJ/rcGjqBwGq/mDfRj9mhPba8cibwMXMfDXBXcdFsnY31
WlcgG3QX3ifqSwXc6m3RjUZ9Y2Ki50+p/hJs1ET/GeBQbyPYFbdL+1uQXdGJs0+Ikioa6DLozSXG
Z2UQiHnYkwjLzKE6GkebDw+OUeCeQ4GxDskx2ee0++0UBW+qq9YWMJbk9y+d0vlMD5TjO4r971yX
US3eTnlAEa6hJl6SmhPgL3QLFxB3jx3fM02upXmtdvrUgZxa9MAUX4GIZ2rX+IaePWd9galBKtOQ
db0mXbJv8bPC9O43qBrVrxKbP7iXgAndPk0Q6NWLOHfwYMgaJnhMaiCygSidcBBd9JJNY+RfUBOb
zM50SVuETR+uhcyTaT1RX2Nv1hteMfHFg8H4Je3MYEfrA5RUMhdh6hckYewTRMFs8ovFGq+RPbCI
/EtPcGlzOIKfQ1PCe+lgPdtx45yQ6yTSPgfZ6LlanWXs2Tg9hHPJPFb/MdahB9pSz36XG/JKDoD3
M0bf6vDtAmU7p3NBvOQ+X9QMKKA8gQpADGraPUgFpjEnTKTZpW6oKVUyu/S9hDNxn/POQZPvVOr6
aDH0xpgvqsl6hdTzK8H6GqResF5Abmhzx78udUYuEt+1Lr0e19sGeG1hiYrg/enkbPSoGUNqDJ5p
q4VSTo3vsuQMW5WqB9MkyyZvoT6PoQNln40yWgywX422NliyHtn7V977kDxUIFFS/sz/2vyHFkYP
AedfQwIb4Ov2Pfu7wcfPdR4Dyk/loS3062WXGQIoTZbLNJSVgRhp44aTZL5HcYU0UvLfq5IZs0l/
koACIYPn44Tiy5i3pwnhNXBxggVR3Ix485klsKNfFQeQObpiU318R/IIQMz5dlaGNqMzOpdzrcPv
4J5eJ4dZl52tslXehKvGapOSJ35kkWsmz6gW3bnNZ70BVdva+6cNnIwmU0De4BWDeY+Da+RtMUJ/
k9rKKKiAgISTsvTtnJOSCzTlCcYGdRjNyv/v/X4D1HksRADKPcVd7n5KW9NdSDGdSRu0XkEKVUfo
ZjaSEOtxyibTS8kZwp0k2yd/3rpZ/SlVVWtPW9VqHulAtomZ5b9XjKYTPFrj+lVflOBRXkX3uchq
yxa4MJxNxacftAxC7We2wlv25V2OCikLyQW8HI648y/jvWcc4mfR0tOgYS90WsB+dQnM7EciE1uR
zRvXo6SoobAZn23qzm8z8HxY8UtQMZs/rI5EuNW69iQ2/apOqgYCwhhY7o0ENYiSgnHOJOMui7pO
461X7QJxE5NCOw1/dCBC7wv+kXKQL4/U89eN2oFClWtybL5HT2Ft6TbyjPI+b3fWg+AURtBKavJe
l967yBaUoRM8G0PC4/By37toLd4orWZpFnQIYcgR4Hjuz9EhBRLzF0EdWrRu/0CpqoXETJ8aC6Ie
ng/Lo60YSCq1Qz+HG5kClgTwyVyxFTuJ3mR4MyOWkfofr91g54YZwZBoUQ77fOTj40LSFgDblTBz
HbLOx5DIL65LdCOmXLaeoGaKCU9pR69v+P34yUFhVsfLE2BNu7yNRe8IIDcgQy1P2OY83T1XqqpS
7QkFxz4Poiz6VJTzOQdaLrFdpnkMMB67hjdzk5JJ2htDJc3Tr0lD1ZLd0T5hTM57RjAohMB+ACGS
OhhWle00ORtCz/Q9BH7f2h06XSF+QfiQiBRl5bpWWunmYflf452BLY3h8CMvyANercWQPR53RsCX
66a+JPYaFIY7fajKOboytA8+RxdJMABRPPQBBWmlZSJA0IopnXVCGLZF5lQA61GTbtV95CGigdSf
MGZD5ZPSsoeBwncP+AJ/z2ZDSKHNqRwjQ2xq/IeIuw1aUXJu9LXLrU3JZpb89zMmogdOuIAdAy/j
/MKqrZZF9QuJeP/JkqTZqhjJmy25XgACjtjBQaD5Jzw9DNodhKI+fOjfKt+41Qkl66UMc09kB/vk
Y5a5qLZfXIDGd1m+qDfZo+bxEEhrwafw/kZH2JVXddUogrox0ueKwibe7mhQXRJkCvnwAfF8vVMt
e2iTzwOdKMQhXCKI8BHWsF09lf0QyZC5bOo68QxYySoPH9jCQr8pkVVZY4/MbL1euYjpBWVay1V3
x4ytgBVJ5vBInzEq3GMEeMUx33KW0TiKkikgu31nHQvYT5IK+3OqX07Hp1sn47nXgUufdLvvDrFF
r5nfsaBa4e1VQeHozaCpJtcxHZgtE5M0mH7eErEViLDWZ4ckpS8f/uZgA7jA6BnzkOJFk595/yVG
fH7EzsFsAaqJUpgzCxtHFZGiDnTuiolfbu9mJ55vYoMYq3Kp3H/R0AWhx4ZpysC2DL1qgldD70vI
+s5zNaLGJe8I1q/1MnmcIIMN0jE1TXREk153WM7j1QFOocuErpCJC4Diz9KqSBEfF6OMGJzthwbS
UFzkFPSnlzmSDMKjWFMQ+xcsrqsiHxUcGbTI+0pDZk3bG5IXhOTPFwT9SR+RujqbNnC5rFP7ZKx7
ruqf/uVmDzkUJyJc2sKcKF7m9L5PQk5cHoGzyNgdOwuRE+VUfANXHxvSa+AwOiY5mzhp8tB6mbcy
eSTMyey00p6xTmNazx5zM3wxKppRimR7K2/2YPqFFL+afso3dtO7xMwaeeMl4/IXJq8xkPpKXCMH
JH7gf8V3zBOaqzMIuZHJmLtHGnY3ooqGUcyIK6QOs5EP9Vf9+3LCeaXiV+FEXv4X9/++vNxhToLA
9YEpaUHjta+USM7cQEsapWBzu6Lpa/CpsjwWEdw/ThOKg4zy2Sk1HtACT9XCo8RWHgGo1btH9F3k
wTfB61qNajjAaf+98xo2eOMvrU5fC3PVGRvbv84iC+d56nHe+wcW45jtmVS6Nq1Kby0j7AU7gEY/
FKoO4nVPk7LV1VL3yf6w8ZhKuJRLRbRGvQv8Mm+k6BEwlkMMx4YJeUZJMZb0xXjbNz9fJJfhcb82
d5Sv8b6eQ0m7Qvfbj3EMIu2oXLNO1oeNu6NRpVDDm/vYAwqwYiOy8o01pRTKFCebIzUWJ52XfPTU
HG/Od1FaZe68ikvxX0ED+Fu6Qt17FDt3kh0vai6SsA1PolgFetg27IYRJOmqWky889pRZtjMfnL3
VYIgwZ7kH6IlRLOnQCB0l1sKusb6kdw9j9iUOaHMfEdRK3u/6o0FqQluAxq95nu4jH1DSV/QrEyN
pMVP5VcTRH4l5ywIFqIC9kM4B+l0q8sOlf2/tKB7t8SuFLAxB0Ra+ovhLlquzEwa47UlkdQhlzDs
fiZZHITSlIMckzo9J1roO1YlTdzbK4lREnBEIffhfEXy3i8VUKJ61bE9fDZEBnRL3i4q47zzqOEh
S8hmbJhc4cfMWmKPJp/fqH+j64kzKclCTd8LYx+P8dpykw4QrRIciZ7PGMHsyF0xYd78GY9O4Hug
3Nk8bRWVIi/sCiL95suHqwudT79Jq4hYnukDbThG6dwgBvG5LfqmhzST4rHySIyE1Ck0pITf6fxL
/99buGDvjYRpRUOK8JMkKUKd2aRppkVEgJNoDjuqqBiam0kI/Fj1XebiO8PIznxGgXTVCKNmlfG5
v72DGXaQ4aVLKsmJwLCMV5I3c2UBgmkqWlwnFew75+nZZhrtieZiMvWLbgosQJYZ+W2x/MGlKN+e
rL3fZvEwZfZzsUgLpczAlhcqqnu4Ata3PkpphxrdpOMSwHe4jLG7+H+PxHhLA4vv48Ys6scKgzsM
8cdS2xpqbY7cNm9SMpZyfAbfsuIjMdn2nC/0oxq1cls6HE8jUd1z/XCm62UuLXSOCr6cVBlbwgve
ZK5aiWXoHbapU7T+urb+Rmxf9eVkUSxYHxSN2N5Tfuv3QHBIQ8Ipp0BXHc9s3mtyqKi2nEXIqRjY
cZxYa1eUlvnHoRmqol//HV+QfkDMfqjwZ+PM/IvjN2Cx9OjxwAsE5Cz5T+Iok9D6T/EhomC9EQ2R
aiSxRIH4pbx2dMr21ct97BfCzssIRi8RvkZuy98u6bgkSNlnuyoorpjEpsu5cYyifKML1iGATYwg
3VK/br5HZvtBtrcQYAt4nrFF98+CAurXPijxsH+7gR4hYVvYfW096vl3WJJxr7WMvQdBnUr4/V6J
B1BpGfKWlG3BZwFDAnLgbGSvZrCaQRDHalUmKKRLwCIjsSvYWoeL41lVgzA37erIu7rZx6+SzgaD
fwwm3o1wbPYVGwcLq9dV28rTulI4shj0xBNIcYu3lM376MJ0zQvOhnsadxWK0Ze+i5Ufij3kZqmX
0AKuHlnS1G69A/EIxAEZFN21lNdlAIWnXithpPGXsHhALR5wEfT185EZX3y3u4EMRR31lN5TektI
zn388M7qKw5KJJgrmDL6sVd91edFSqav9xagxnJdEBypsFg/7ggZXKwWVr+PFW3GmFe6Zsb8A2Il
G8GuqaKHLU5fqZcHaRXnWLNHQABjk9i/Akz73P8cWYgCihsu6VEbJCUB9YWcYtSDHnlUJp18l2kd
nKPowAtswcWR/7resqqXoi50S8cMs0p/7BCq+XkFX4hcaO9VCp2Rsi49o54CEc5QBYBAmHspYxlF
4xMuNSu3arOxZmQAUQ5Yh0+H8sUQ8n8j78qFHB3ZrDc67lDxR/n8cd49rlWiNDLyN7H0hiLLkoDz
cZVzojGCPHK8nTbDAuH2zZ3YCIVXn3G+YTDOvOK1kyjdF0EAwIpAWedLMuA6nOrmK+YvZInXIp2T
OR8UreshTH0jF0YRqo5gBFFswU0tnjA/zDnek8QNQ2KWMJFdfkcuCCZbU1AkXq4+1VXA2k1Ig++m
myCzJVEaeEkRtow/d2sEWp3pavz2e9zjmKKsoJoMpcKAN0RdWUJDK0T4NYBzTjklwZxGFGYXy9ML
KUHZhQ4P4cog05dYIFWss0aw9azdPX7VSltjhKbf7WWvnxVlRVkOxpU2wDtvYwz2EclHHFZIm2Rw
uQbJySp0TxMPtShhaDoN9ewWIRekcur5Jcl3/bKNeaRtK9EwcP6whW2l0yyulH5X3kS8wfIJynwR
e427FsqBlQn0dhlYyMfdlnvtNsrPDGt6I8ptWlDP3YGCL1K8O1RqsoNH6qbh1WrEQVwM5ZDz240l
h4NF8u37lDS49AD0kkB+0ByOLCRjh81U5E5w8XPn99vztJSEZxzaf/xpwSSSd/mg1FRqX4Ld6EM4
GknOQD5JRxWeZq7lgxLAckiTDXu57KsQyMbHovhFrA/y6WlHCARVSj3l/ZMQ/F7Igrs4Za/Agls2
BYw/qHETq+CYoO2jD60JTwCSy2j0PCQrQRnWEwHWutS8s8RFdIOTq8332Zt7szoMb6wQt/mE/9x+
99z4m2jcPsb6aigXFKcszmMMh0Y5gkTLjhWUxx912Ou+ccrongGC4KAUmjV4Jc+cSCb64PxuAN1m
pIUpJLimoAhw9yfJGZHrVtvwQ0iHkwau2ZcE9mNgat5v1cS8EQDGtWRR3YJWowRWSJQz9rJEHJQv
5ydJsfTcKm8REAM48xXNU6PFMDaH+byMyt941TdP2X26ugjX0dBCUl8YJ2hF862yUJG0EpSTTtx/
KNGMwrphFBM8qMZasRr8cUFcsAUZTfKioJaC4wVWoq1yxhb294R+Djh1ISClFf3Y5p8RfQK8IOer
P+0PlUaiWlRHexcyQQ6fAD+Yo6DHfj5+sprEhEecd9WzcDoSL5z21o5ixU+sDT2tNuHjeOlijcUz
0FV0WsPV5uiPm7BiCrdWmql2jj8X3DXtAU66+WBJdh0G2kkpyAle/uhGqUwjXzUfih7v7QX/mH8W
dBA+y2/vTksOcd9Tna62Dlvt5rC1WriHK2EPooDF2hakKHNSAZWIb2V4FFczJYwmUz5V30gHYwsW
4pcWdS2HQk57Poo6RsSjQx1YKW4rLH8Kf56T8Y4KLvBkedyXjIlpTU7cfFZ26FzlPFumZmSVAqXC
vuZF5H2ayYwuwlH/QYgGI8oSZC44vl9kKX6aiVVjUvyjBaX1NKppWwmSdqobo/L6nI+R9SqY64Gx
qa5mz1uXvf6uyq2SUdyaH63E7g3/2OeDuS1gapVbLdd4aUm9TrLpdugAv9f+dsoa0ObIIifdwThg
rTn8d8WAw5/Q+oclVFQdLCxJkzm8GvBQKr08E7QFYd3NntceI/DbxxKA1IU63GUa56vx0T1NAPCa
p7L/TrA2fWv9TBYMmQKdMRz3iyybtgnsZrbIZ73AE4HRg47tNeRHEhDmMlo7lF6RaKF2Z3jfmzuI
rIOONYfYCNdbGCH9kHQ2NsDYWkyUdEHyrImxsAC6bg5opZwS+O7Gr7emGyg/bkRvruk0r+c/GhkJ
sQcBrXvAIpdE/tTx9uU+9e8+or04uiS9UPylIzzg+w5Hzfflyy1/h38V7Vt9Cgix9fnUnPk/rQn1
xOchJaWm++vSE/6WEdiIWmesxZQzH64Jdk3aoUgW2f3tyhWj8WBFx/w2zg5ByuwYsJVD3F2EWCSr
FiOzp1miywYPwURlhOpZx41QkIrJ4kIXrP8WiUUfrtzaq7N+NrzMyujpOvYs1plsqaIut41mo6xe
AjzdWz7ck2H4hS7cvPtsyojEeC/RyKgRpCYBKHM4vop8NvMEGWLzpJME5vUvolsNAPcv4eX3h0LJ
sshG6dyAs69e3Ar0x+LW/yZFazCleonEj2EwNy1NDFqvVlsbUollkL1gZzIzs5UTv1XyPHOtT3XS
wI5YkCfeuvkmR4jIa5aZUirLdU0sSkZrCyxVOSvU/YrSwiyFgGus70cnm3azWKSuW/16b8fx75Ey
ShSyv60TFqRWnI/Z9PIkrx9YoVZo5YWPMmZoQdhPzYKPxnYEr9ZnwZkJUtHlGuZbFauzGUEfdYXt
IskR8Zz2OeXel+l39GZMfM00SAPdTfvQyZcgUP8w9UQGSYuEH+1RlRwfkV9sloAGyzHMFaLA9hUc
1mdEMQU4smDa7gReMHixUdXqgx63Ti/TxhswVLVuYQnbNUGxmZqXixUH2gh67KqLYywhOd+mCZCX
yKXUg9NHqrimVe/uOzjQDnKif5XF+dwUSBVB1fvoXEt91ipEOk2hdoEw6QcpE2Zguxu91GE3AyIt
CkkApu6q3bIxAun3PZCHxrLhOQeAI31xw48KLAyi7JGlG/W+JQNWjYn/0nlgtfQU+Y9d3ttMy7c+
jGVBfJJHaZnmiTQU6quL9mjNhhWzH+2x+VrZSbN3XFjR+JvTw+HOLMrw4pj1O5+T9nRoCYPbHKBR
zgZEMp6pSk+WwoxPMslmq770PJuAnJlqp/NGfigrMUHtX0zoq6gWne6edNTo0y+vNW8PXgI7aF5M
R0kpfLbecbLtmfCZDf0hdWlx+GfXxAocdfUZLDRsUTC2f71F2Bi9bY+4smqjWcSTeM8t2IMtGkVZ
FFWxJV8YStUuivkz9GKjiWzvNjp8dVBilKvJF2aab6vGuNYwH8k9HusiWdrbV/Dul4rv+lx+Amft
qUR5g1U/BWVwGwQa4pWuH/9pVqYSrBIPVpa9tOAdrDz0OFFkyXji1wxbKaRe1rvu0f+NCCJUUEku
zwNQYXdIToo+xOIKa5Sbatdp/bpFFEU3+/X+tVdqfv443x23bLxUfEA8BCUd4j4M+zURnQUY3pE9
ynLCHFgKCtzz7kGQXW4wFCSIOiZisjRC3X1aXuw18LK/rGuSw/ry3X6R0QKIoTw+NOVC1fQnn3z0
hi17xAF832uD7TZYeAwhfgBKHKvtvAniYRneJImidzvs5xRf4pzVwMWRNyFPAHN07EyCjpuef4nI
vwhC2OC6Tf5f8XccSD8DlU66rG1dcrjkJjIPVa4ysTricR8km4SABYm4VUPCLUd/l2y8Yu0AhQBF
WmKh5dnP0dv03lbHIWBL+eBx2uGNooHHKF/sgbntrr5OhaqKdlTtvxBXn7QIQaX3lPivOsbg0xP4
ElBRkpHe+jz8W36uk2CFIen+Gg1jUrsvAH00kNYnBioFZfs91Lo2ZTpFczT0IusrD4qemXjLmTHZ
7ijpBpToCMpXi7yLQbqqLr5TcpHlkU/sgxYKtHqlgbdiJCvcT4DJq5HPjGE9OAy5dnpX2dSlMLks
8GRUkCmiAw0krJxtIbfwVeFdsV/+tJSSftgRbWLIAJZCmpX3YGb3DOc+71+pS8wx/X/s2hbiLAae
t6xINT8Tk9m/JzJiIRjhBYAM/tuoZQ6mJiLMBR7ItTf4fT/4RZ5ZUrHJss8stfktVlQctYilD4/7
rmMapJZstEhbMIVr+9+heF+nkM0NHv8qVx8gythaxef1Aprwp+m/4l6SY7KUKk7+zRlhi+LzCw3k
PUQAx96q82TpaSGcYp283fWgwZ5Kzgl+q5iPMma74mOPD2O8J/4M0S/LK+2lk3XUSM6+XyuBiSA3
ja+1j3Z/TqNFItJzQDfnct8pBMnbFCt91YtIB+//MWfClyD+v6VrOLhw/Ue1hK4pYN3Ye2p07nVM
WCRQ3lsIKSMeikEyLBIWtMdtBjF43XlOe7kGNQKq4PZHFAP929DlSA+UA+tHYaa6KZ0YlLbT7KW0
OeqkNiG18iWwmk3Zg1UcttVv9ZIHn0EWHRWRhNfpqBrYfv2PhgfB+JQ+lvbRD3dL4rpqjGRCmUl5
KABktzMp/Ztq6PhK3PjLYG+1uVn5YCvBaTssrBfqs0U1w80Bk+rdUTHZIGCg4xlhCioBDro8DYam
/V9KDvsHREWpOo6T6vJMBpA+yeeAwQXxFCyB7UvOW7UA3fY2QLgdcQ4U6U5Gcc5yqTKv/oOAZJGf
lvWeGgV4iQVq7GbhD9NnuFXOC9Fmhw3CqnCgGbdhuppOGRoXgF3qor2qPJQWsbN1thOAPmUHS/oL
vq61e2I2JVbvmAwbVbKqYact3UiUj/qr9yMvcPUZ931KqvvEHGgXKec8SWzjf8HRDb4TRcTiGRJs
RRZZ2A6/u165xkGucQRFwOidGAMe58pbEXXLwu8FE15WBI3jvoO//lzgMUEyP5EISbGJpiEhW6us
zYs7aCiHFomaNiUjpTO3BQ7KXf8rbt9KQuIWCv4v3ptdsjXG/fyv0BExjqWbO2VbR2kAvKZgbDbF
IoWK7g/zxWjlpogOT6ZSmdBvtEkkRVcxXiH6sSR7Dt912zRlYSTRk74WZd/bpCtjdlbEzAX9pcKk
rGIW2FrkibuCPVaW/ISkfwrtWK6NEfBwKDGabCJhQZGorT3TLit1mXM9UI9Iuzc+NxYzDriH/O7O
RlbpqSwgCI0zdNVd1LLLJDStvGIYSQaDRpePomga0lPqs5yng0D1ej8fXD6lr0RLzPbQWcCqlx7V
OoDeysbQm9aXgw+kz0Aj1gqdcfz90BUbfOXWMS9GpMzcv8L1fZKiS4Vbuil9OU2rQlFvz8n0S69h
Xa3BaRytpiHXiYePLmMJsVhuwMedeOmd/oh7veMXN7XTjY6LjWe7J0UyfhbzBj2AFftiIlpevO6s
kZxpmWp9K/Jdq0ep+O8abMK6Zw/ivBRBy35Nke/ANqdkn/5L90lE43tWXdRB2M1Xa72yIxYrR+VJ
98/o+PKi2QIaSBY4Iq6BqbfJ0uXrldWdklyxc1eNlrYd8Xc7xpqFsV9l8LeJDQlM0A/b8uv+RzsU
dhFDrcCOgnjOg6SHDXkxWYkeMITtYuRLHkp7+aEZDO9fNv1mVBP2HKiPen+41ZOTJtnj3i1RvL2J
vbbxFfCFMw1OflWzZPUum1a80dDDaxzR8S+L/JXW0/k3F7nTSNiJ558VJFI7yO5GcY2gqV1EC3j3
7bXuZTyothkA9Pv29NhDjgbigiP3oEh1hcfPi8pfnLjkgcd+XJQ5ctssf7aBW0DSrD5L/FZ6D00+
534ytvBHd9R7Bwxgog/sEbXRqymmY+azIkh0BcxpU+B8NUl5ZkBZifTdCKwt/m4qkc1WK+P5Ewgb
BVR5tMDX63F8cli2jZqGCngd/sTtqdEYbR7WV76CVLrgkHhReb5pEqfGXGsEbhU21SVQEJRpXdOs
asQpmTRqbA3vPUlR1m/WhxUjunrd2lYRVKErqxVmYac10PwCTca7XPcfWtu2QkI8bkpqSxUw4cDc
Els13DICtK5wAtHOniln9AeIv6+BzlsIb+jBNmHOilLiqUaG7fjErME+p6+VoK+yFE1SgkOQOdE7
UHjgLrcxjEA+zXzVOCJR7k9yAU0SU4M9RVaSmUiK5YAGmgv5W77LggVmXzQxF6L3BLfw+6yqA/pb
e6UsRd0W+lWpqh2mrUVwp7a4eZ7ILy08vjfV/45Ik1GLagLdFFRhfgPiaquqSNs/0SxIoTkSaxAV
n9bCXU0X+3Qw0JE4A/iCAbIQvbV4ZOZuVQZlQsx0aFUbCT6nGcreCgrNKOm5fzA/gm5YMk8iSm/8
gNZP2+LpqBNEdEzklJCYHZkxnthbX+B9emjlI6j9O73QQTtMYPvY59o+ZhDXd6V+ya41SUF7zcPk
HwM0f6xFmHLwW6+B1jww1j1Zf1Wp846mq4x9SCz7Se/6GEGdIP7B290mmWx3eEv2b93Yb+Wi5RrC
xGBdEtq9XR9WuoxZWjYq5A0eVoQ5KFO6pNk1Xkd1TiINr1O48qx6elt28SjZOQBcjIpsEqdq7B8c
pPE60P1wFR6WdMSDUY4mLejB+ahK/wsw40UThHbvxOPVcF3QgA4Xe/wJZgPFqT5REkQCO3jBMgRQ
vSfhBD+bicMnXtMqlWsLgJRq0D3ZLwlFppSNR53iFU7FNWs3yElH+c1S3lvVf4I3gRvZ4d8d63i4
etD4L/osc2mSRDjFTJnRIqSfEbJ9EaPB2BwG6iZbpSg82SiqbI1ikJGXqb/sobBGelQE0FFG33/a
/BSJZ4gDGIiXTjiD0/xt4qA7K75aMxosZS/BpeRw1bru6IqsEiMygWQtZ/AP+ujJwRuFlVqFYALy
E5wP1d5blfSqstNUdfWc5zO0QswLbZdEDa5+ZbW0kSnOUnjVlywocGBMSdTPccEAw9h5QvJSgVQI
9vt9kdS3+UtgiAeX8KFpzEA1xUnCUKzfgVigPPxNvcmbBzrNn2UeBMXibmHynETNgm4kJxNAWg99
Qe00hav5OugTkfr3bYS40F2hkhoJXNCG4BlaGP7fxeelYbffTshjDEahvPfOPNDo+gQw8DoWjL6w
h+5DGhuGFM3mDKRDc2YOKwrcDj6HjzFPPg+33X+5eNrQinKl0Dg2KT9KkglkU+91yX33APVuB0Mx
FqaHz+/e/4nDhDb+j8u8Lw81DjsJ7dx5M//D8xodMfbxEl2x9UzAvUB/ymZIHMZeWn8dNsk2sa7n
wIaHfUEe7uEe78Ti/A9afFDha6cS/vzaSV8DQVtvNxMCwxXNf3Mbm7uvitE/JRNBTkENOQXbIple
UsOxg3r9CKNaH/VVV9Z56dYItUScQrU/b7SMcsbI0EhgSSN4oUDPaHAPapt/2x+Ara1X5cWw05hY
jYH4cmvaU0zhtmLZV1Q5EjGT+oYnzuFZ07fYI7iDhhLRNPKFoeIpngigFoCzmstCsG53kHf83D1h
r/5sKunRS2HBzQCkl5JIJzqBj738LslHVfd8Rm5m3dK7M9pr8hz7kZXOG8pE+aJiiyM1XB3GTJGO
N3kIoITO1upRb7fVGbOr/mlaqhxko944DchyHRotnrLcUJGSEluK8/KjbkhZXNwY8PARXljKrxbL
n0G5aKnjRhOcG+BomEyBDdaDhn7vIRthceowali/UD5xrFgR0qjmUe8Q4cWABG4nm1tLmNNZ5tij
viD+NdMO22efc4NnV7Hl3XNs8Q2SEq6hyCeZ8B12PqFEvQkF7dGbSGmlZqAHayOLT1V1orFt6Mkr
JZpW2CgyjONn9Pu3Ic3HtDbpIY6rlPspHuDOhki8ekbdPrAWAC7CF/2Y1FxV5JYaC3C/N2PBvOu6
aLqvp5mSu0wcMEfLn3KX0d2J/3dakFi7uZq091R9BFKglnXqdxtDC4yt7mRFGGRUy+lgnqXkHDuP
myy8ovzmySniWLVZdSc9/I6w8hYsO+1JzWVCmaWzdKcTF9vYoCGVgYAy59AL4ZVHIxeo0Y6tGxpJ
Ii1CyLjUpMZXAmRgSenir5nnmnjuek5H8DuK4tdP+UZ7i3IXNspVYppP7awQ3nYpDaOtS/SoMD0d
b2CpiZMFNtG/ntKBhVTM3fE035KJcaRcGnw7Vrozb72vilSOBBMo9eY1aSzVa74uwVWEebEl1/aQ
C+WTm6NRNVojqyPzDAKgQ9KnUeO6RzUV+RYr3JwyY7d2zgOnPJcR0WSoiUwy65mGvIX4LsA6bICC
BQ2x7spSqKwqpkZ+V1S/lz6477MdF00A+8gKQLVUlJtgOfcosgrrcm8hodNV8tDOQxxuGehiDttF
5ca8+/pyegWR6WQWY9Cner3QglPqo+dzzEcKshD5dC7qECEkrQ3Q/U75pEihDDP0InDkQ/vUtFir
qhYDL3invrMepWj0RieWzfsiiheExpjkrH5JOqmvOo0JydsZSg8UIXyGlxlAxr18b7kkZhtY1hGL
eiC/Pth+bughcP8xS5ArySFFrN/c4I5TypXfSFlq2sYg1+rvJD0fNigCw+y21xWnn2E2PC8VMWXM
BRgBdAdwJ1sN+ZO/SK4WHl8GF0LRR7HXf/tl2mMobgWFrWpdNojdtmsGX9FQtOL5JciHdozoJrfw
8TFx7BhmYeNljgWN5LA+AdLvnvuvdVHEZCtP7B1NMe8UTxol04y6Lzkm5eEB4i8r4a6pLRNgSqC0
A48n4x5SRo8MUSJ2VtVFxkzBhsMqKki7N+bPRwWkNfF+fYpNgKrd3bRQ90/CJE0dLkZ92pJH1LNr
quV84JC6UVowWn1fx+h5+SV2iThIUoCc+CBEyh7ZOPnrjs32nC2M6tPcetJJ8zaxSLf8ayFOXd6x
a0JOYNsb+MlHS2+Q/U4ygdAXfRLul+W1vkO0zSJCZDDgkM8GvMtu/nY/l9qyJx2QvcvC+m7Umjkc
181xwbcM5iQa3e1vARDlhavW9GqNca9znGWyElruy6dVrXEwZQXsaW3XaOr/uM7mId7t9vo27uB6
eg2A4BssPU84GwiAD92CGhtQQqnLdozE8fD4b4opK66469kHgW9WjsmSVKeJlcozfMoNmrdVjTns
wpEvWUz2euXGzFyJyW4giTzkcnj/4pgZ9+JyqVoyW0ixGYIcdBH6Ld45VswDW1nPCVMgHgXr5bOw
15zUDFlj4WTlh15+/Rwk+j2pD4xWiPLO2OSRDJLkmn1d9XRRa3wGsIr4ygZMVWMAgQ1PNYZV+qRH
C9buP2tC/Hm4f32q7SJEYo7BdDYbMudBwipwPBCogClmfvjlRgwCmdhmuYC54Dcfr3lbLQ7YI02a
3qto4510CcZG5HEhvZeJAUPn039gAC+JzwFyaCYArBQGSuQyOoTdHHkn2yZYSaKjrEO1hA171YrB
MNRWM5h5Ly90msHkcNdz+RwBojgM5aV8WsT/QYilOMvE+q8yRo0jDLQgrBi4T96o+OGZ+Qd0gIXT
VG9IzUlhMotB5sTn83/a+HmHVNrOpPVvS2huH06RNrfkpKZgtuGjY9fiPKR2DmhCwBviswOomTdc
amjHCtLVptugiL20pk1ZaTig4EV0h2pcC3GQiCWH69Njm/DZxJqa9Ca0HQF81JG0/KcFS2Ds090A
M9oPu5PQyFjUIg2dzi/51N/6txzAEFD/rTK+8HiUf3MWaARBaKnkP5glpOaWaHc22F45ThgiCXmO
SZV25t+ijVuXUxOwY43lS9X7Qtp50HG6gikLLHVW4hCGJIJbSN76BI86b5JBZHK7VPhNm3g1FTx1
SCLd0PpLTTpaRlscD+ZuWHwtGdjMgCssqvnxAwSx+ZZg/HOLzA8NuuyZIT3J22bgMcoTFMpSAT4A
uEs98f9KVn0hRinPrhyHoBr1klSzBPEQWvSzeiN/yh5dlIA7SLOhIfPhRe+EAxXQ9Yh44hV7BCW5
fAWSmqaNCuhQUZzDVR5op2AAkIHctzjUAXDdETEMYm0MfQuk7R2i4oBnWBNBgktWEcJbzLCjUZob
KabhF3rxmnZR2urOlSML6O4pt3rkr27OArnyFxDR3sWF3a0DngeCnuS5ubCOwH5PP04zHltW4K+I
uTfIsQdAZTBG4DyeycmjMAU74Dox6CdhOlS0B+rH11R6k/vTl7mCkiLILFEwu4r4fVwb+vCm5h9l
ihJPN9jodkciuaVIILs8WJn1MqRiZ5Nxk3+BMrANhHjBzTzYyXTSnSA0AClWBuyO5aw/jKVJ5M0y
0an7BFlPUtVGK25Cj5WXq7CAUmoPsUb2J4SkKsbk6MVlpt5yQt+egyNl2RwMBoepO7QXiH/PKWm+
FD0pLnElpGOHduDtly0kswsHQoyk4Gs1XHBrXjDt7lFAnKsn+LlGTc5av7n31W+CW3dllCzdbo/t
3X6p6PMSqb21epE83FV8EnB0tqLw6Z6xcIPNgG3aNKrewk7cm2weJLgBSsDDJEwtWzkAop7+hmIK
wc2trAF6FPgFkINUw0tb9VuWpBtsDc24MEptrSgQF7HA0VmzTzYVMaYh2IIAZn8tZFN71oTMmJTm
x/vDGJ62R3pqNfguy4P3W7t3gvSRJQ+6aRcV3ATJKHOyBBNQn+OjeMCdSoaW0bwkKbisze0Qsfpb
/fM+uvEC+g0k7diTS2iDcy8DwOZO2t0BFAQogz59bnotrmW41rFxgXTJglKNAquoT/Q24EqYMln5
3t4kibAy7fNzMhtrZX9YAQmXT30PPoDkO6jm3stGBJKzYX2Mcn/ozPcFheWFBAChUoyYe38xgNav
jjmJf26bdt7CYfrxWYnSrpFsrAeKopjKcuHgJb99Ep+XFAFzbzknT2LzCXxTeOAgGiMp0Q9P5613
qRNMzyeb8TRlWU/T6aIbsDuiwU4TxL6hynFmMBUMtQG1/p3a9nnqG9gkh6+QLh8hJHx433DJFePQ
xqTppHNQLV3PCw0JJQpWTSz/yVy4BH9ssGN1bE8YCb2QY8/ZzfDsvEFvxOoUXZUTR9OYXfgmySOz
V1eWteK4Pk2spFxfjl733XRa9ijwtCLQreLASgQuHt/gtRu9dILvXb8oKGjA00kAUs90b/IjnWyD
Tm/XL0QRT+6pKS6jLuWrfnbaz1NEl+Kak89n0dCfDsWlUrDVamTQ1Lu/7C3xv3kFrdNBiEPimaRr
2roWidze5EGV3pSAN+MG6GoGW2teXP8T1xjVbD6d+wmh2rZhFiHMPwUXD/zYeqoran+DBpCERYM6
LvJroZdudtMDZj/adBDNQ2XxgExVwZTWSp8IGYGqv+JqftKZFH5CPyS46b2HBDsodHv9goYd7b/H
G1qx0ET8zLhTNWzwKwnBlqwb3hnSpwXcETA9PgWVjmYhbdnRiLhb5nkVo4Y0hAFhymcy7V+s+5AQ
ui0FC3rt6mR9vgLMqmUX1v6bviJIO+O4naVNc6wUtrjL5kZ0gJ2XC3BYvgk3MPaEkygk2AeUDUFl
wzA9XGRyr2SFTRzut9KvK0jppcyaZe8YWqorC8ZXPAM3CSANcgeNGNdqpEzp8k0Wlphpl3VXmnq+
xHbf2nLqW9/Hd8rx8YDIJ9Z/30ebjvWibsRZczhu7sPqr0+Rcflr2PoRbc1T/OBLHxvZGVy5zXSk
xqbaYpG0NmG2UAt5oitJqOdk/d1LREo+b8mfnBAY8WpYtdqiPx8Gag7vj160LttVeoLxFpoOTqBb
DQTDY107h8kCHqqbC8gR2GF7SaLakeoP83u15PSQYiyvV6Ak3m1xiuYn+r1vVpn9ry7yfvaF6dSq
Cp1oYqL43MUdSIobfZRj6R9EuiPWof/DgqlF9C6UsQOY6tgcfVohwt0nVYD/ufxnCQVjOvsFmO2V
dNyopZqsgP0VhKqP4MTRS8lil6rpOKeq/F1ZAka21dn0SqKtCxn/123Joikol/BLK3nF/yIYX0TC
JsqY8dOx9nayM3dAuA4RH07nirPEYnY4WfQAmHrY5vEi/O9nVqVtrTDTq5Ei+6iZGXHvAjE96rCm
W7b82Bc/AO1w8fSsnhmDsf6AxuDCNf/NvQSztTUd5WY9nBy/HstRk3v6mz9Bs/Ua5Ovs729MO/2g
TTYz8WNy/qM1as9dZMGeOo99m1ntHftGKq0OcifWRverJZ2xTmotImhuGEPKJVGpU9TfbDz5rx4z
WrHQOFv/kInCv75JMrVGduSAVpzlWNWEiXu8XQZOGKgG3VwhneqBb65QHG9Ex4+FZjtGzqNznEhS
pih+qGBKX6/5BDp7S+CabHTtkSQy8kyBTFvn2PuX5KwwQUPoi41I0H0mF7XdmJRTZhUnwe1S3QG9
jFAlHKCo5t5Fj55xoKkiqEs1RcvghUWZUUa5g/tvt/GRaRFPp0h3M3pG22ZtKQe3yyFH1DaVFMy/
0WA8bUl2HIEAtJI7lSKIE6KlT6h+sIp+XFJ8S6ZA5BwemtF7XI3KdKhJdoiRdajcpdh+m7MxSS2y
Uz0CCFcqWeXK+54VvLDUNyrGe5xkJnj3Mw/AnT5PIQhr8C+BxXajW896uhc3z5Klo7QVGllgvm0U
WiBDe1EUf62NclkDRPC3Oebp2Yk+Q1Oo7vG/zl+dMkRiNhYWOhFTyr6frZHsq3xAgFuQv4B4YrkZ
4z5o3e6zSnr4FkHllruffofnknrr22Rew34iK6HnDMlfE/xZSGwGWH94GTFzgggRHETqc1WG6zez
g9C68d/n6SVGFp8OcHK3fU6WGY/a1IrdWjRO8bAB+SEZwVX9baej4xE/i+m7AU4M6jjB1iOyAoFm
5IBZV7+xl27uMqQkOjAjUrATdteX9LdBZBx8WGQbf67PKfv4FVfTTaJrBmZY3ub8cJErl+ex0m8B
U6UmYLwrt8pfkbK4qX6rFBGATSVOPnK1JUegnaCDg7lqelImmC12fgOuhTXbg7WvaQhhk5a6GTfy
sHuR57kHqla1D3pqNvwxOgm6/TgG1lX3fceHNOR9RyVIG1qaGm/VmMT1w2kqEu8gSZ15m7KEAErc
3a9fcH8LrIVFmx4WAsWSUZQXrxKogYtT3qkEJtkyb4g9Uu4AwDXlLoLJaq/d5zH65nrhFW4LzCXV
VAFjmH7W9TGiV/VF0YxbHEMStFEt6YIA+5d6p3gL4cXJXEyB0Du5l+5UeQJ/vxcpd3Ri0kJpc+QV
tD9JK3eDu29KxOWLowrqNiIcwcKwXoFC0MGCn0g0565HsAJ3He+Fyj5QPr/Vlije92FoOYE4c6xs
sjX0xhK4rCTDwI1yTdUus1hkqEGj9HrEK8qYRff1dIlsg+mvICYYDiCvu8QnIg+iiTV340/yAk/H
vPfFjY0jZfXtwKgXHoTIzxY1k4hKZizFe8QeQWacuubpckjw8DYdk7g3msW1/4Fv3g/g4wlsbnR+
TvHNtbKzlEF6+4/cCliCVGIWwDfodVXYgwd1H1Lz0hdB4/uIQaRHnvsg4cEHJUEpWu0KhPRombQY
CuXGkTCCToiStX0sPel9xiCx/107PkXVFKMugKTBOasDXzEZxvPT0gOahZDKq2ErnLboQ0DbGQgJ
WG3juFhug8qyGRWImhhHzvS5RcJGH1YQeCIMEP+DPNjbEbMtiBs5aLp4XzzKr6pIFL0Bg+AzVxFV
ZiJQZ7uw7B8Xd6VFb55jrtTIw3UsxH2bPbSXBDlKQzVwkVq3jsx2Hl06Ebkmf67L9b2ekDaV6hVq
6q3H+urNhvaAG3KarobfqdsIRbVRraj13qnRwaiVIYjTSmxhb8K7eoI8Hzigjy9Z/kwh/1/eEhbC
3FqnKK0/U8Nj8dhMxDlZtT0qKhTniO+07BNNDmeBTKDonrQ3VVqkqMxhm181BBO7vIiGHEKXebDN
IoVo5dw8Q7f9z+jc0MrjApIR30NDYX0CdB/wtBdiV8H7QCyID3OIqommT+h8IFcg4O20/5Y+0wIN
XKBZrV0gMUDdQr4CbTdTPF+SF7WZnfP32qL06/fKTFAU3q0Xp03afnFv1fP9vpn8Y3NOceufUBOM
T5E2UnXCNrD20bIvcsi3rugh6CK/I/GMG+t84taqiAqJv2LimdHW/537Fbk5bbxlKRIDoPTQETHI
p8GvmH0/vgYVctXarXrbfKfICqlH5kuh2t9piMq577LZg6HPSrveg/GYF5oKCKd9kKmQ0A+BUuxv
umDKA9/FfQlul8o2jJ7K02Lrv3+iE50EqbimaS2uPstdYQpeMbE6dLfyWrKSlEClw2U8l1M4ZsAm
Wfxegws9m9JE/9CcOZ+5QM5ieds15+eSc5Zu4ZonG4UxQjJNGGa1yZgM1bxTne9dnPC8t8lzQfNK
ziSjp3yOdb4N8Z3WXjqAOGpRhKnFQgxyGdzmycLxxGP6QTk+5xYbGdJNoA1UWSZmjBgVnZ4vsAn+
lJyqFcXojKzUBJp3czTDN9FwB/8LGrGZteWkyHSZW9OcvY7IQimRr+BjflaMnQET6cKPR8PtouXF
k1jbQpA7y+2wNodDGJIeTLyBwi1iqrIxnErstKN4R/fmPdONBKFxTiTWc/hORlB60gKf/GuWtoyN
m1Z29/IF9ThXOZl/epnfiFpx8OXZdow/Kn1WgGyYSWlP7DwON3S3BjlDJt4T/PTWlIWhMwT6Uhkt
jtP/mirRzqImRkZ8ElNxvRIeFEnt8aAwyOWYoQ3sQHKmD1oN9yTswMRzoocRqDuU04aTzKu0DlT2
5M+xfHP11DuYPq9o6vgRVBmzNWK2Uv4LAk80RbktEfb+TE+FNqK+OP0aUS6CCGLKjXaKJafd100/
dgpSTUyEXNRBkYp2aN636CP3WkgbVwsaemDRwox7V1d73Pood2s5PkraSvn+xzgnZB3ZijfzryIh
S78i+Qvs6ljHgllhufLi2LxKGhHTWGvYd2IwcZwjq+1xCdWxx+7s7oj/dIzwuOtGXS+2iwt5OevF
J0wxdYh8PCsWbnGF23mDtIm5ht6a4i4X1CR6p7alagW+mxXudTkNn315HbhGmUzFCCwTJ+7QegPn
YJU9d/UgKccLec7n/wWn3y7ZueV16R4i4mHQHNPhWYGAYBe0O8AS4rzYkpThzjDhy9THkPsXxEpU
wi4jBKduVeriS7xVQVhtRWvY8KLEPCXSTf6pWuhdFgIkS5VwhR7UB4CVC+oPE3CsXCBhRVRuRJxE
9hKdgT5UfKXessFwLwLrTstM0WECpBsHnQJY7WV6kBOMIbMNoRpAn3dkbq7b0P9eXz5woF2v0Jvm
joUvbs/c9bs48ELqWL32fc+vT23t7JLPS6kEE4+0Ux+9jVUD9eWRwL5VV9goNzuHF1ZDrozzMA6d
noZqGPb+8iCzsEayNacB+1zr/qScTfAyAHzhEv2NN9ykxYAjZwX0IbkhgusofknvaMMQO1+n5HzQ
HocNcLCmKiEPi3k5t9KabJw+Nh3jJSn1Vggl2tDuGTBZdFXKaXU1m9NwTFzNqqspsred1qjEMgG4
EHRR9fIkYMnD1PLPZeHjvSMwGtiQnju/DmAzDR5pFNKAJcKKTEzWT8IaExornUBIqAErUOQdolbm
TgopfmvVQ1laeiHbRu+J4suehpapvxlu+6vwIzfXynKMvqnNyxWEw8d3J9MlBl9aVwprqO6D/Lm0
oR/9qFguxpi+8kzsFo5gPlR+iWvB1+2XR69EqPRjd05g038vN50X7JFcklWr3aDRU3y8nnwnlbbt
S9NoxbsZ7tdPGHETeLdhRM53GRYCiyitAA8bNEoHlNJOi9MszXuD3/R+7JxZ3FBkKmbTYDS4aDv2
BMRq607KegnPzZ5NsGxB6xASai9WsTORHgqNzsdYPLxSWgyaLYiwcG9IC8Vryj4IVAuprKxkv/yP
5GTELeIr7YtiZjxb327GKoDfFHWYsZblvZxYEjRalWgQJb5MoHNPCrVty60F8cKdh0JVQcewm9jj
ghGInIqJbyuB54dqQjCsk527TZAmcql9CvdWc6kairPk0P9KgERz5YRVRWZtlazLvVS4naV+OZ6j
nPpjlkOrCYbKw7HtGoDWGlCZb8IAOOC5ycYT4xYyGvlDNwYF6BNcDNXXk9GMQwRh8OfFkQCMP5Eu
VFS1k1I4TK0KG6rTOjQox8RTc7QscZ/EE+E0O1P0Yj9ReWmdHcmgHrHebJiMx1iuwcmxVBNBc3fU
bfloQlvrQ7Wrga/zuZhz/m4cMrjJEDQOC6pXZ6l2cID6tXQX+CqYgCsE5MUQ9UYyMHHDRFhS0iL6
Sv9y7CA/7Ywg4pEALbunJAKQ1v8UhyFGFmzo/+kgpfLAEBh6ecRSx405eupdPzeC2a5m2DxeXM5t
xvUBDV4RWiASKoEo00uQtANB7y5azr8SP4SQaC1kJ0gsH3fOALSTOwGoFEKhy2JVNO5zSVb6vLGS
eKN0wjz6Cpw8hJBOuougB+ADFi9Gslohv9HuUFeX3qonoR5yXm/2I1bYrPJfMHOXFiPB67DWIGXX
1E6DrHU+QPice4Eu+sSukH1VQQSuUeM7RF1D1NC86yoVMBOHK0iQBm9ztl+Q6lBbniNeBy1xZ6ZC
2eTTD/7gTkPdBn0KsrjOTBX89V+q5Pl6i2Kp9UgXgecSJ4Y+HRIj4qZ3bxLuComM6qZGoAIJ33E9
EHacNcaFwlTcefQGSIRlO8gwE4y4ZeDnzOVEe+sZ/A8OyXpj2q4UthLEwubplahGCSWzpstgsAN+
lSlw6cSfwHYVZ3XVvENR4CW/afZb7jaw1lbZH4YiAJOjugkn7G3gIq2TUMddfDIsn3AO+MnDpdz6
0baCBh9NvhNCVvh5CC6FKa3HhC3c//yKf/LKnv9syf7DhQk1nXizdAm/Sqwv6DaEKVTwrYrmZnw8
UOWpd7QLQTxKcpLs1Mz1DqoUgVePMogmiWZSnzouHplxlS1efZdOnFnVN/r5Rpi+kR5W9xJ4tsbG
StnRQnvJehGIWReg+YiI2E9rojNeB+DhHr6kTFulDRZCWJGgGGHpPQ2EuJ6fKyvBdcprRlrOeU6A
thQriqQ1LL2mSI1ND/A+pAA5YRzNWvIRYYdMrMNQUOaZQ9z41hcITqslz2jQyBasIIVvqCUvK79v
8I7RbrUslfw8cI6tA5NSN6KmC5Sa6sTHHKt+xiyzCGv385j5bzxFRMSwPVqixVRFkaXNsmmc6N50
tN40z8qYWHnuvzOYdUK0zvMQOIPNVg2RwfMX8GnT0GHn35vKK4ln6w6L0r//bTL13xNIxjqiq/tP
r4nzh3J8XKBX1s0PCEzFU+GySxiSAuauFv6N59ltYnBV02EpJB6sS1pL16PGI2Acc3rnz4oPZfPn
ojgqf1/xojevL3j/9zMd+piutZSNYq/pFHqN0z2rEargM8nHvP3+3yUDRCw28BcCcyo6Sojg0MHm
k+sf04ZBul7asd7nMnwBWMS8Prhn65fHK757Db55adOkgJUJJd7w12hbZkMlzvJ2j0kUBCZMpaWc
x00wFEACIE3fBOivJpJCgP7dnvXE7ck5WURnHHJte1gHEFkZDweoPdqQ2wADixtI4JNGSNK87itw
v7142c0T7t/zffJiknxfZamfMRE3PYZaR/a/Fr/VZ7Q9ESqD7UWXnv6pQ3fM00L9j3udUqdqtL2I
rQpcs9opZJ1vrIwe43R8xRRvBrJ3C8imVIyiVwEV014iakCjUhJf+pWJ1U/4yutOytuolsfjL559
41LwgcUcvgdTPAnuzik+Ic04HYbjIXZ2jqkXZoDB9JKp9Qw1eclBrpfLavgW1/DMSxxvdtxxq91J
Ayu8VCpNamm3ZG4mt4hSUJATG9tMzxa76Npiqu0Ur8wkP7YDu8h2B4y1bP3YQc4ptKOMd8Dn+jx6
3xEuNU50WLCUbVwGfvM9TkmLe8m0BoPq5YEQWi6agprh/zR23ga/y1FuPJA35sW8JgEcbYvjORj0
hVWsRTageTKf22GW7GQdpk9EBxIPB5TB9RdYkbN8sOkcV2RuYommqc6CeuUT8Hx6JtV7wWsTvHr5
Fe9Jucn2EGMCIek9W08puWnt6vWPr0c39gvAVB9uDGzYrowvzMbcbzXyYjfv8kIIJNpRQYkZb5MR
4Hz3mNLA7v+FE+lB3SOkGyXo5KfYV/UXfNnaECqY1y72mK6S26eFprhpN0ahlLdDBrma2UDlj5Ld
eixEMOm5DzVfP2KqEaYPb9n9B1Cg/b+dYqt39WoUAEKcZeimHa3PDPOnuxtZbThhPLwWlJhCL2o8
YmAFXOxW2U8rPrFdIPRA0mLGEJvW9LYjL3VVcBxzGRzP2IzCBEqDNGOkqmSc468hLeqGE/gRgH07
qeXa8lDgVtRAdyD2UY6pn1VjBGE04m5RjOD6zsUsoEUkLGJ1/h+txHXj4jQVMZKjcUJenq18TH0M
hVd+f2xinepMKooOHAB0x9KBSHADK3DwT/kXJwNeEBVSsrjh9XgzUlyerhxErO/nB0YdrNld9/4B
xM26wRwhh/iDkcwFRohslgQAjopvwjEYy+3V3iPil0TjF2OGAzWfJ/7PmjH7V7G5ViIizeQVZOLX
AgE8O5um6IinPsh1QnO582TCVVAy9O4+6FQuuMBDKjQ02rTA48+4SVf2tpZGwM+xSafM8PFdKkIx
Q1a3Sv1UnrZ6WHt1uhiCqWa2w6kJwNVMjsQHkTBZLv+TNT323+wxLNcpymndQ6FIuZyMRQPUREr0
lu93iTZfMETasyjGVXvK0lAdRamBIrVnTx4+QehdEx4kk6rzPEQP7AwuvTAt62RbGcDyDgRSuZdv
2q8aUst5a2TIZObBuMF7SKuq61Y1cUYLwFm6C0k3vbtmcnQ6Q+0fxK2nfKRW9XeBPNZzsLNYIa5O
3mI+kvQU0tFY1kck3UGtapWG3YDQbpz1gmAEMHhG5a+koBlufFw3WmvNfv8a9hEbVWli+Git3fTO
Cl9F0PWndZZPbg0mkYVybsIO30AHfnC2wu+rtu4wVZ1g+wKzDhMSYYrBHNYYt+0Q7m7g7Q+JKIMO
kTH/WQ3CmN0AsTe4j+jmsPQD/ZBSTXkDFDUFr8jvtph7I7D8FsulOkjDjK5kFE9puo47RQYsKj1/
zadUCThpUcrc711/yfmc8j1LXqSFnDqTwxVFXFn9l8m1WYPWxHjXEeWAzPstlhJkttLvLwOXvaqD
Cd6kiyKW96EAHEWuY0qznLCw2hBFHhI9AWNYR4ccM4iS9Dv5BKLBq4D2jUMf/uvkpUoAcybNUwwv
peikxPiPcrTCytkMktYmrmKreqeGCcsb7gg4qn9EQw7IuJcUVDpist9uY6EMjCYvlxr179WHdsZI
1AbrbyDv/II4U2+WvAfXYM0FC7YYxkJxlFB6fW46FOxnhyYV5lCzewJxTGBHi3eDiADBTyPR6vX/
uX66z4y5N51MDZRJrqZlJzb3xQ2iF5cdQi0BYvA7221F99aeki5NtfMYchFQGlzxazl/9x8lD0jj
/11lfFdXC8b3FvH4feIQIXUjoClRisF33SX6+Phxj0N6A6SOvdW7TPTLkDZ48YFMmWddGauhdUTx
xooRwxpjB3eIJWVqNipF8TYrf/WdJPeRIWdcIDbPr8NkxvdWVLCyhWQM0RIODT+QCi+xKaPTEe0x
IPNBlnolp+FYlmaMtneXEOfda8WqbtNDke6IY70+8j+dfHujWsIM6zwYRyG/bctEpD/A5ObOFV42
PEr+vOPxSbeDCo0bndoRDEMO+s1duIhR4w0JglPKnYGB9ADKb5+qCFiGbGgYdv+TSS3h3iv+DFLm
55RvWHVXQKvkQ5O6Smnql+LWm9A2CNTBavyJgf3sOkE54VaghZTFiscX+HrGV2OgDJIULL2KfOFu
uO6CJILmx682EPNm8hJFXiLWLAPQALb/M3xw9ETZU3q0+Ihz+TbG9P3JTOEKYDTqsmYOpLk/zl4I
Hw6HOURXEV4nHDh3cqODFnIdRLSnM66ECpJdK8ZjRpDPzc0FJMjRTyHGzI2pIB8Xlfs8P4Rb+gp/
Bule5ad9bpWPeXFZhASWzDGvFK/9b/mqgOWZVsk3/Zgn0rIbVxSGdoZVQb3G1srWSBpiyYQHCsqi
aFmkMYTmrtwJjahjVkOJU/M3AzdyA8rud/1OMavMEp2MwxPcElyc05ARkaVa7uOCGWHeLLf+fB49
sEEcA5rGWb8VilQRyS2atA8s+fsOl7uMJMyNUYsNW8JZcMSImlR/1QyFsf9rx74QEPMZqqa5YX2x
6jX0NmleZZhTvlbhV6nPS2IvgOdFemzX9A+j+uZZlVqDe3yFpmW3YyssK3woi3eYOdtKeLZMUFd/
XGNDNFZHKAEFrC+MWXjNTtpMPL92+eyEXFoi8UfCmDniOhyBGLOqh9Vzmj1P+O+ooNBiU96S1Dv4
G/XFYco7gwuugyTz/O9y76I7gefAr4rhgn8PttYFW59blEpMsRvJfxkKVznRov5PUAgiz3DuhGSl
VJ7tvpEA9Ct4bI/zRhPaXDgxkQWIg38wecqNlqVbRDK0Z7rMsP5QRo3c+drAlzdljuGdZz8mDMsn
zc5/D/W9PiACFvbkcDsddv2WIJGL8/jR/wF0xD4LXhjrsSmkBada4yevfcZebphadCxbudcXS5f5
vfBWF7BANhc/8El/WtU42bN1+Ng2EzzSLUXUmoxk1ugFWUi4gBscxNxLZa6VTJ03bKeSpwoQ1lQE
pdy+BNsCXyfpkJ4RxPXvWzTFpGekOyUP/OnArrFZR0LKgYKi3/E8NdEsGDR+XJ96LesEhSm057am
SUiKxd4WUqjIawTGaGMcuoI/VB3oKnCYbArWnwoqp5WcdkV18tMa6ej/vA9mNPWJq96V2+DGy+tC
t7kw3xQGr7LdINUiL/mUVbOipLSFAY2Oi2XNNWWqbSpVA6cId9gC/COrAntjNoPYFI2OVxDuZbxa
VHf1ZNBku/3sneCsz3xtWSfEHZ02ZQhk9VFlx+uLhmgO+aZi/QnXrLITM3f4SuY1kG59ZFfDKABX
2VF9QD6HJ40ijlxMt2C9grSJgdKGByzskRuDJWnLw/te3xeviidlYKQdM2NLDMfa0oAj8/4+W9/b
8FDU+qBNYkSS4RlLGRwYCf8VhhiOvBsDKY97dMW6SK4SkS6Ppy0+94/8DwgyWVoVDiSK6KILR5E6
wDHqp7yoVdFlD8XfEhyQ5obDRS4v+KOkJM57uNW+S9U92NK6sdXTSvALRpuufUPCrIOeyPfKZtEY
NlnxBZ9mUORnc+rnacLKhkJemIdqgVeYW9xsgTWgLg2WS2stE36Bv1/iwk74VdNjkb9UjMjotXkd
DQxRXCmffL2ZUAZfzBrrc5y+ejB8v+VUXi/tPbQk9rUhHDkKkieI/NbCtxFd6Borzt0APW+/6up1
bSsh3wcm+nH9CIkNbig1XOOIMi+VFZ3Mg7OOCUsOjostzIsqaL6tF3Vp0PyAVXoEdZq8jm1vFUyU
mmLgRNq2H6n0V/JsODgFG/cTDburtH+8DCgW85WIy1QYf+RnYqIMsC8KP42XgINHjBtNE218Km2o
1cNaVWYHpVuNxLvUI8f2L3etWkH2um5QxwsTdxtGKAp0OUS7k4EZN3OxmhnmJMQiJKvqR5tL907V
6bX0LK9lGR66E+FBKv54d07bmVd0xtPFGDwDPb0IkGLwg2OhnlXUus7hWL3tWJpoKPv24iGliauz
1Uesgyzn1BY9IcdF6GMKTPk4e0OZ5cRolFKejdaGhbIO01kI4F7wHR5vEyKdeMmfFwPYHLzOiGPE
wQAuKM9WZpOlIESJmiOnXxMJXeGlBC7mUd4satA+41TPNUOvD2yMmmqHG5rcvvIFpAm+ZCI965Mq
T8VXr9TyOiCaOx0ZGeFpCH+PllZe89t5Dl4A9aAaroW2JYYVYGIOOzqbGS0eJchHM0kseF5fpWPe
wV32+itzg8hE+K/NFKtS7VZT8JXm69YtRmyxoKlr50kkqpoVx3Cu+TbTatZiYo0E5TfQKFfSQhFL
HZ99XcyMa7MW1UThyvK2KcNqJNW6Pqjoo4RiUiKoduvkSZa7it/3GrzWJ+lFmSHktqbUK69z9FkE
u7nL7iTyIVL67MkrflsWROpGKamS1WeLjxUBzYmSJny6yjxMIa4QsPdbY+GA7KiHyl9lxGgpsqUC
lfmR4AdksWkXrfcytus6p68OuulAOVVIiG1ZA2D7GQ1Lg1kaNvAAcE6Ey7EP1THU2xyQ1XzGgqrF
AiQe9E6rQPJkyGVWUPVS6Tq1EOeb86utOgjXmp3838eq1mRtfJf72acYMoG2rbMX9Nzd81fkAUQd
Of9RXMwXS5ZigliTlPZJzcE3HvEIgHcDYP269Q7oGj5eXESfxDyC3nu4uHaWMyInNaGuymJS4wIv
6rAiO/RXuutUVj4KbUQR9dIwracVTsWK0HkXx571D2TpzJmk3qFuJFMfbR+1hPK/m6mCT+pc3lV4
1eY8TsKzd3/XjJ9nHvRxjOR1SjlAYmQKX1MY6JRFPkhUyN2Wybky0XBiaAbU1ViCtdc23ySt2B19
BHCzkC8EwPNqAZlj9bLhlyjokMoKROR0BvOLC8gvFs2W5NGbPHdn8xRLE/zjPtga8Pa1A0AS7kN+
O1vBZmyvmnJjue3099spXUB4mz8chW53h+hqaN1d29srVVEhATNiGkO43TsvJOlU7ROeAsY8zH02
O4XDRqhF2EnqENWwrG4y8pro+5yMSeOCiMZR1dUJowGG1utexkg6723YNdzzWC21fkfJ1XuUYyFc
v8YM5u1+ompYL3Ho1SAXH3fhdV7e1VmO8LxPr3UzY+5OiK0WOe/+voIp1FgviEAnVsUpRzvaiQfA
CTxxTjzD123EtToxCJCBu+YyvDO4JmQzolLRvI7zsABlrvwtOlUlF2C3/lncxotmqIvjYBEUC7FF
ggOnjvB9vqOXyHpBcafZPzgysCyLnRfhydJjdxAaVY4YKBCy5d00K7KtI4nqNlPWQQGT3SddeOhG
tW1MPF0+LuyxlbD5CaAY7gGfaYI4GPgGR7Q4qhInZj2EVeGkFPeQ+IBxL6TcNuuHfcRH7pFhfxBb
oWlU5l5/IiqlZgTILOQu0xIFmJGqZjODavVifDee0wWZ19yRK+t0y+Fwprnv7VYimmIx1LIXkwfz
l66R9BBb1a29+uLavPMFRH4jl1lN/j1x7o2byOBD/QKObTvQXSoDP3W0JkFlWtfTxeuZeo1njhla
E6vxB/U6OoMugn7nvABZo1XBaxnaQ9GDMTc2oAF6w582cYCe/ONBe6TJRPXGXSZAZRRy8EZP2yMQ
L4Vz8JfigcgChKwqgHcbrEe5Z//xwrVwkC9V0ttZeKM4MOtfR07wXVjQjwx512VuHxLKPa1eKYcZ
qy4kNQ18N3T34GSW5JmIXRGdtTE/gTa+OrJei+LZWx+xT5F7BGVWEqdpj+SKnyovc0qyloM4xcgm
j5/VEu8DPGTW4J46RJpjI+Xlb15voC4GFaf+THuythHgBOPmSPEI20s4KVDhVy8J7qPqm/c1MjGr
SkTHpyFcLNCRHhZ2QPOqkrFh3gg8PZGHdukzK8pPhIuP4e68WNbf0jcppjJT8xttEaqUvryf5MY0
1GGKIVGzAJrxvA8WOFwdpRPFfjpxxDjyOGb80OM6Mpk5r4GzrhENNQnuw3nlFbacW3zCUPArkmkq
5QwQKMtKuWCu1DxhpRRB6l6Gv1TA1axvhDk3hWoPcM89sycvAIYG8Z4NbvnBCsRqz407D7RtSwNC
36x9snZjJOkk1TacICgQn1jNtVvImauuliERu9dUJ2d7pmD/c5Atg+/ij7D7Km1x6if00b1y+mUH
ARzm+lFdtkiKsm+sllfMMBpp3TT1u7n/BEpteDWAU7Xs59j7j+nOblX4zSVzpwKJsgPyuu54D0GD
I9BPfpV+5PoreM4TIJIBYmGVwaEOE9XgkDyHcBx2culg29GR4BsHXSbkxtNq2zs9VzPjDKYHOhC6
oMUPErk52yQnwpvz/suPpN8LaqoJcVI6blPlv9sJX74/9d0TA4VFQGKvqe7xgaYhvfDlo4dSKGn8
Q1D4DGJCoivY+2JWwn7vTUFW1HYwGxcS18Y98B0ycKzvQJ0NPLgIhXU+CLR5x/kqPZ7A5GWliInV
MHHEfeZ4dpKKx+WgOattU/a619dQtezfcLcBa/moAAWp/fgcJ7cxibg7+sHRMaERK0zZ3X64wxUO
nAYEUwl4EhNwh+s04hUJdG+BaZmEX+sgFQl0uZAK3qhMjDDgS3mafE6VnhBX7rB3XsF3yAd5UMy/
xZ6YsOIDT1WJWzAp+QUfE+QL8unr1iWdjgFS+PE55QbWS1IAR3N8TdFoENM9dC7+1FXylqNWsADZ
xsxI032nHbSxlg9PBzrVyDyQcBe6i/2anCHDfSk7gA2B8jAo1MPLnlolhqUPbfMSd/th4vFWIcBv
BJ5lTxXypNa5CKw/fgsjLZ2uHF6ILOsCshThxT54PxVCXhE7skTmuvkEcZq5WXLg9MSEk3YMkFZL
85dqlI1YKroMp3hlQbwlFty82ioMjMQjgPmsGv4+4HOcIg66OM9UhOIbzMVYV3LuQCuIUTFFH1NC
H2XkXqIvtBZJ2ssiUvvgHf68J2Dh5tvh6O1PgxcP8fcgJmtp6FrwXIGpL7WpsXW2+/+WWD9+luEC
ALssnExo8GmNHGX7d5+jJ+eosjq8fWqtWZkrPrWCEjk8cE2bE3q4/gqyehWYgvoHCNHAeFfJ83yj
RpfyJXrc2n/NIeCvt4yKNTvrhhhjmchKtzr8J/B9AHl8K6XckbqCFMF5+2OZxrA8hcwp5bXEuQez
mJ9ATc/4ev+EtNPs29JTlfWvecgOCrYt3Eege+NqR2u9+YECLsov1ELuBgZDAxqYwNych2u1JbGZ
5vJlSv2zoQJ29cHeU46/lxgAJ7tKiIibFyBIziacPdV4rGtIseLldOZru3Y5Mru3aawdc+aIOezz
pargv7laFKpY7Utu3gAh7+lREg3EwB08KKDGMr+cNYsSZvz2YCk5On0TaAVCHLeZX4sSo80NnZSM
bMmsbtXIJiuHV0TYiD13xIQOr37a3K9rO0NruYDmF0cC6nSMbavD0HVv6AXR3eHu3GI+l3F1Jc0k
an4TkNh5Ns2porofJLK/Pzhg41rl5b6WgxeSbYv1XVzdtf5HnbVm8qIJXOTVHqw22XEAp7uZH29d
VY5OMFJnX446ig1EQ77vraFFmwrAAvsk0vYX3VfWzkr6JpTY1NCcqGAg7Le2WEPDBg2YcvAT8HT2
X7TIO4+p7pedN0Oz0XJ4NPhBgRTXhL/5dKToFwxFbyzW2QXXpwTxTHpqt2X0vUZ6BIprnSYGwe8E
MMqxxOMMJsJ7oISuLl9hHVc2TcZTwCxTj5XFuX2OuHIyYIeHyL8WwM+e9AlfvXAG7GvRShTwhRKD
m/PCASl57eH3fp2Ce7X0DMPVAOqdSXyFBgmhSIziSnAhxGRXuAG8w89DTNQoNrUxhvdDIG5JyxAV
GCa6+woptiLpgQ/1hEEyXdnSSFPSflI7t3VJkQLnn5xKsNMLMy1Dhz5JOpD9GXGQrLHf7fAZ180h
LL57bbPELlDg9PT1tgFurzGqC5mZ6bFlsYhMDblhYXvqZvTzlb0xYWtXJzcG4Mqpx69ioE0geo/C
mArLepfjs7jGKNu1HdZWsRI5wnooVZ1hJcO341YAx9i6kXlDirNGeB1MN7lczKQcmjE3gY0quCby
wGKuz484cP+Ro4a2DktKA0zThlk4R+QUnD+RswsSToHdZ/l4jWN5xGF3+IRrn6Al5zi1OrWBTx4/
r3O7aaEuDAPgQUF3idY5f1x1Xm3kouiyFinwEeT3WhtIjwvmqbI+rYUFuJHVzY856CuJi4/YCl6K
1fKbYRsmsJV6j20ZmTsDgRLY6uIhxV7JaJXuMp9g8wvhQ4VPGImo/NhwKJeYGGWWzX+joUL+rQiY
6T3fU9WMTCCFEAC0x31QV4znNInfNiR7HPXyEED5jpdAelDfeWW2JEO994D7/CfAlb4oJMBGQKNq
rIIHtE8+xavbbVGUGzS1Mpj//yKSBHlgS/UPY+h6lqrN5s/zQn+CUzxttQS/sTCgEVKtrjGeLrMP
lytwtgaL0foRES8KPumKL0tyS4U+2wXd0J6eZp3B8fZQKZLd3NgcXOU7BSlxi8kNlawKAmb0sItr
/XSxTcBUd+3zNeJKaXyV2zvI80kKi6kZr34sgCUri4WiRJe1/1ONBm465NSZcUWYN86btGSPD+zY
1NdhKCbDBYcFG7KfmTRceLdY3/9abcqGE+tSW8CvvYJdGBDewxYjXKy0q/d1Ai8NPWQtwrkvBhh2
96oJkhBm9XaJpIi4XbKLRyiGdA6nuU8gzlcujD0vhmWU2RQG5KXfNQ/Mf81EbCvNymJ4mipNSJTc
R2SFH1wPo/Vfwsmy7ucOA32NTEvRiyOhW3yKuXF6PDPEq+ev6J0rrf82vlLAEvKWb2qdL+Nl/6uA
Ij0IabA95t65sEOH7lsR7rzP27w+KBwys9KtkLia/+RdWV3ke+gKtPxMLUg+ufAMp7YSrtvruDFW
U1JDakeZ9nI5R9rcf6UvRhdWmw8KGQwB4sUS2iZFX73QIbAu+1bORUeVglewMq5beaKcDIr/3Kpf
M/jnn66GoI4oX3J9EaMvROw4hZuLbmoez+6MCTpMzkWPTXb+ty4QCoKuH5VmJJWZVfoBQIGcFD4E
2hmKdli2CgZkukgrKogKkRjbqBdleu6ua+N5GPpZqpPIBqc2gDiNbc038X97S3gw57lF5yd8aQZ4
cQApqiY/jJ3IsAnpSYemJTXB88dTfYbMmMKYdy7/Gf+YnYAbgzSIQUIoAbcFkjT73Tc/WaCyQLzL
y7DoxgmuCj83ubJfchvN7r09/pBuczNvb8oGkzsf9LQm/gjpukmBfONRRh/lUpfTuN/gkdzU+gTs
5s/bQoiV4/WgW6kqEq2NYfh/Fh7dHtfJBbQdP+yMn3WVgTYNdhBlIyJnjek4Elft/Xr6FTTieWS9
ZtfE3bQWxOwmNHK88CjfXliP2yekCPTOMYvlpmn8wOfShva+6RgQpmgfsjbyA7S2Mg/WEn5jpQkU
l24vEZrE0lNVm7DiWfbuu7s0UfqvTjiddfHyvodKfsk25fasEFyMMTsjAowqMyac7o85XfPNuKxJ
VWMs05bKX8ob29Pl9w018sAzzsxLP6NAarJf68zKRPiOM99ZcjCdxINpbRB467cFsKC4JsFBqKEb
HXJwEMMqbbCDU6a7L3LfCZWPHCrXfjmrVoCSCC9N/IRCGW5b0//FfYkteccWGVXj6oZkUiYkyq15
3RBCjghGLz1uRNBe6TTTu0F8FKtP0UPYK9UKazm4fy6tmOeNrnOoEx3qKOKFCSYV3GO6+T03kgEd
zNRCKTaaYiLhn58eJfF+l8zQl19NI5YpBnujq/vYjuKNidagY5q3smqqVL+bJO3TwmNSJOjg+I57
7b5PeNvbNRRF0lNUoFTuJ18YNjNUvOCl3UXYt7YM7W7DL5jn6uwoTc5VhFpckcwbbHUk5rQG7QVC
uUxrwj9LI0T2A8RFjWE7TaS6OzeMb6C2JFzwEMEETfDXrMKoCf9X9qXbRRuTaAilaF1eWSj4kJoZ
3OFsOyOmBDlU6gyPNJmVi4tE7rv/v83UJpkgQK6PNRZj/mkP/Y+oyM2E0ocD3K4za7QMjwPS21Y6
5t0d4RFkBgEPdAz46/NABTS3bG+H1e/O7VhaTsl3ADV7mHbx9YR4QY2wJh4c0xgoal2Pqkanacn+
MdI2xS820Xw6p3cwuuP8sX4sENIlzmt8zh3SRoaurbjF9m3glNB1b72l2ZOEiNJ63boYGrgIPCuD
atw8k0mqmwJ9Zxapz80B/kEAKOqIgE7dV1BVmBZDa3k7M1edY8c3zzTLQtbbGUcw08nUXpkU6OHn
sXuSUiZDzP5uYHN4DtBfjKbJr0qEl0uFGR+lzZGqIghgA+hqoPNlLewDf/qjWeVhI982BFFtijOl
Wx222P2dsjp9zlP+5fj48thUBEaS9jWipHu+84Dz1xwQDk1qmGyaaKcrZ/8P1PC9TiqqgCG/KZSY
e4gJW0EpZEM6JY8TdHu30avWJjklSgFYalnPkIDF4rQHf4a/JBpTQXkny/I7evl5E68VDOVpIwEd
PXxjeGM4C520PaNQ7qlG5S3ZXhrUDNZs5wUNatytS+bhNBlyEW1Lr2YDODp6p44GTQBQHOI4JVNU
cQCGZTwzrkNmGs14XOnRqqmaiIudmJTWP750JZlXzpYGkipZP7Ng2UFsOHafJjA0aezd+VaXg/Ao
KKux4PrvWGNfZWmzM8D9LbKlDL+hrXa8CiZIQAmMo+ZWM98pcu0tldVlEhbb4q9LlqsD9po/pAga
o5r+OEhjU6ciY+qRpmH5KSTer9KtfARpa0tZTmNbXVo9TeqHUKMg10mSJVWj5iUjDDxJvgn1W2on
AQlPBoNIQmc28ytBqLc9s9n35qR5MtJ00mixAKf2R7MEknE/0Gv2MkMQ9AMOFs2OZcUy0/U4AYJS
8oObZStYZH1B5mog6wT1su/8jTqqzrb3wHUKX0edAQk7X4DwK+x23Eyv/Y/4bsb58nrC8+Bla5oP
TCm8aU8y/oTNIKVjIJaAimh7y5gCbdYzWkQMw9o3qP483NA6ttUJgyEID4z46EqQ6RjEv+2oKHzC
8UNTCOtMVntueOxNomSwdqErPJ8XF3DRUoMty+f1DasRjJftb2/zS67eQBxzXHffyVZAQVk2PbC7
8MT2PR7ncV346Bg5HZEW0KWsOeamNqO++O/VQpwDxbzcjTaKXryNEZ3ZY8g3WmqBP9Q6QIG9hp+2
z0CKMNBWRYVG+KN+ObHJSvKOIrb58OIxG0Vz7EReeCtsB2lsFqEqH7Bh+rf/0n/r8GXNgwYaOqo/
HDRD5uNauClrLHVJAuRhWvtNguNdxJVdsGnaHTLzZjJeXGttY4T+vYw4b++qWHH2aaY1bowjz9OW
ETbNZHO8dEyHf2CjPsAwi0AHFkJuSWotX22w6XIba0r6XDSrz3lCaDW7pXXMNeemfXWlYmb9CWLc
e8wsOjsK5plQAdYukyUgCD4MEdEKSxXl7xMWriCKK/4HQ1R/1297Qxb4RsHuFQSeVJuP1qLqXfbn
29B5Ka7bCTogmGwsgCmqJiinG6xlmGJin2e/p/hw8i9JY3t8DfMsAMK4BbgGHULh/UJp96DinQIV
nLzMlAdloDqywUgFO1z1cHNEHHNmV+3EgSIEOvvlbsrI93eh5FusMgohZ8ls7qHi1kV6AWRnLsfd
Qc251Bf34d8awcQRT1OQKxMkwzvPayTvloik7zhrKeLlGKzrOXRS3ImKRlpyeKNGHqvnRBpUgF5g
YOx7CXOy0TZFetO1LG20zzfPUa+N4ikYoL6Tnetcwc2kaqVV3gh6sVNimFIW0iDu2IUESZdTyN9q
3hhMy7ZskdMXMVxgYt3llWlHWji01f9c9nhWjCX5cnk/RQJuXMo6RtC9i9PHJDvG+K2kIF45xPq9
OYb7K6PtwoA7e4/SMMUK83cZPZ1458Ivj0zQeoO+/RmeiPWkXbf5NYgl/Rf1cmxwcuKHZLFPU3ZD
Zhe7l2oL9XWztcQXIzBvKC23haWniBCn9hWWjmLO/TwIC2C5QcaKipOgJxMqv20bK+KGYgJw7u6X
8u6gJvSPSceCwAP7m13y0nb6Ib71fDL6TSDw+/RpFCoaa8MD45ZPUtdvM7sDKzTvA5dO9BbbfVcO
B51KgYfeoPlKp+yOP/zTBm9pJWwRa/M5dy4CW7RMyeU3pqBctxNK1XLU8OTQZgmIKVApEH5M+PoD
n3s5xcmVoVcmnWB1Zjprm5OaF5EhtuDlc86edamibji3+f8sAR0Gseg0Oe4cyB4YOuPFUFS4a7XN
ZESL+3B5GCsWGyMmcXnqJc8HH7Xbp+XQgiXeMIQ5GDyhi3oxCbZDsOBqVTBFC1KQe2alfrWmSL6p
fnApkCbQEQOm/cj+YisQ/qlyV7A0tqBSxcp4pZdChPvl532Luy/+NcWP3n83WlxYmSP5m80gr7zz
gQxcpqN7G7NeWiAsWZgbkohXIl23wlLxEqC5utq6nPrx/FRm/RS8y+Tls75uXUmePm7ZPyHGhe4j
LPPOyPm1uVgNz7eTHSUfu6iTSS6SS+Ocys5XIiI2ZSuZvUIvifyQs6fxSd4dOW74EBTfe1FHY+oM
bVAnfNF4VUF/4to5RoLJaOVA0ocFmC7BjoLs+an7oYdlQFSDVPUPts5H66VTgeMNXmkaoElEkVhZ
Fg76tL91KwRAWo4JtPZQrNpUqU/z7ZLpddRowmkAbiaDVTk0qt5kO5xYNASFQGfsDpri+PZqIp2y
B7aJnmwHT++R1HkC+Q6BQ3XwQ5R/FIy8in5BY5azXWDNEvSnGf+9VrsBmQvvGTAnoj5KJyiPvpE2
xO7SP0NQa9B1t1UpdNjyqC7Lf0dZ6RDVAsbnBeGPNzAjJSr7FD6ri2J8ia0RzKW61Zf183QbanRn
P49iN2Rvu9ghuLJqQP6Ngr5YgnHXdgH+Kt/Aw2HOCSxYTqMMlMPzjN+q3lHDeiXi/dEBHzAeFgsz
Ks69Zs/DQ9xspDEbzheF73VrR1BPVzzx92Bd2cWfFrnyXY0hA71ByWmd+RSVOzvS1iycnj/Mm3xA
IHJ1t6JaGyuwcPAqlxnAZwHm5TlfDmckgfL8fT/EiC1reHJI1rsMXb4OLuXXlNb0Z2bSkWuetper
FrufGpu5x7Yk4wjA0k5hkCFdq4Ex0fz5vvPP6JwWhhZMWfZPTDGRFxVWR5hinFm2o3Tcnrl57dT7
z0ZQxQJItBRJxHoeFCEifuAqu7HFnJklCUkfPspkF3cT67xvoFXSyfs3fZgCo7D/cohVJFYS7wws
/J4vZzykG+/5rzKHAjKV1uB66iEsMNKjbcRszIpyhHTcZRcsW9V0X1IPUJXYazKEFCm/IsjKzouX
gp2RS2pAB2GEe5te1/l3lyMcHOJsZw0G3Jr/KIqOzo+nbmnkSHffxtbWl1WiLFu/qFYkWFlxLm8J
zMf3MOJhig0/hz3YvwoVWJKi25BJL8eDUAkm0ETs5SehjCRxnKEBblpOAMas2nRI1vhmPxN/LoOt
IWCj0qFNoRg7m7ZwtlaamCmAs44DwcMPzM2n7mHGFOGAshiaD3PZWuG5n6EdTZXalvY6a+wSNSKK
UfOWP2mX3wjEKIHa53cxVrVCyNBhc/irgKYq+PZd0B1VwPeZlkkykj292nYBseYmtv/kf78i8YMk
qqm+3ZUSiXB+iRwiE5DHplrKtRSzyGDeDaY/IvMu5uuz3P+ynUU++ulVnpljpHoYnJCWbRs7s/HB
18aUiFhU/iZEN3kazNANXxw0c/4NIWcGoEFCcYXs8sV8KpHh3FIB6uU83ponv3BzOGNMAanOeedC
E66GHZYCDUDF9h79fE0iKD/5mqhGf6A1ryEkyjb+g49IBjBRpU5PDVokoQyJS3TRrJYL2AY5df/B
f3rI4xSnfZuiKZbUKkqyJt0SnTSIQF+w8/t4iXxwoZQ/6kR/kqUOwFLiy2EL1VEtubydv6hQFVWG
MfdzhZ/60jNPZ/qS06rzN/m6GxWNdSukKVxuXW9Z25xx4qkAGtli0p1qP/+Fy+nymTk2xyteiyjm
MUWJwpYY/UTo44RQXRcOtsUqTHijmUjjM1d345uKNFAb+QuRU+qH5E1xBzsAAvxpXLBxsJncIn48
Wzg7q5bLcAWMO1qPb548hXdUzQFzjiGBREETUnEaE3YBY78plFJ2vbAMoWKqR36FfXbOxgV0CO81
i6GoU/IJajzg9fBHBEs8W9PnEUNFpoB/PlbcM1il9pbb9hsSIBpYvrrvzVsSWis/LHeQdS2+mV3t
V10ahPqbMT+Mq+gvO172pbjVYA50mNKhks4leJvmXCkXUkPi0kx/BQrBFE5sgsF7glotmH/mFZmx
wjFZLuJ6Emq+FdTlW0/HgmA26WgzyzRO4V3qXSYEAAwFQCYHGIXBtnVV/sqYskh8PCVRnHR2NR5Z
Zthic1o8Ih6x7sn8qvKP9QrUv5a/EuZg95QLQluE6t22EUBlQKfk16lRsjEBS3WN8nhlGdpedMfG
Mbkx0y8TuK0+MmQ6yB4B9hCPoV60YJQ0jePJqa8wcT6jLhaIMKd3iRxHLQobiGUum3ZiMJhSHD4y
agkWJPZFnDmgVISOoTYiPF86Eyla7Sl1Y+BmaYu0Xj5zACDaiotFdQ964Y+zuzpRVg7DceXsmIUh
7HirQGaIGvQf1uzP87NTuKCw1XpgdFBQ9PrxJ6vBdacqTPKfBV8mYYTNDJCbEBOxN0osEOTwXkxN
r0GVRrmF285leXQBbR97O36nTsPXRRwVPlHrg5SioNSbuo1zvCkKXYYX12kDsHpzvBT8qHF7EjAi
T0+yJnz8SUbR2SE8GBIEWzMRM/JjD/RJ8VUmH0KCVWTfBtevcS9tqgPaz8iCMzV36Hsl5CRcvMbm
/A7ryuJzKx/EdAIu0YhohlClR/GgHeMwtkdAPJh8yqGiLKV5zWjUewXnWGJnsZz10I0+nUXKLWTv
tHIRT1KkFSD6jlH87ymUIOcHMu6auuU1xNKWoW8Ng80tyAjsIdBcpBKNA43SdcMi1xQ6Szh7NEkG
YKFyxw+pXGGa0eGc8emNUvQIdi3ypkPWf3z0wiVzosAGRElj15Gc55IFmc1I+uJm0srfIIZxuTfS
q4H+ddh01VNTdaWmWfRddANrS//gO0WUdTqxOJJfRsFKGbnzf8i1iyiqe8RnoduoKtB5qVTd/yZj
cwwKwVEzwBLvq47KnV9rF1tLrCdSQrUeFtm0QC6D08sP73QqzM+nY0n3jx9rLgFqNIitcm6/bwub
siD2miCf0AZLLTTIe1dNAkHGwefhgbhGLea1Zi7OBGaeRk1GXI8doxczp6+wuYzB65PmV4qjYulU
Vr7q0MGjV+VndCVC4fJ0tpe2yMr5e1oaVuFvqBrAiONHMeYwJjEwh2uASMjbyux41yVfvwNKOr33
gAcY/9VCr3h5/rPzUkfACqB2K/5gsa9gvdVQdZ732800aATqmedGJRS++aHuk7DmQp6gQ3YEzZns
5ADIlI29qj6EDsyyu31agq3GsgOSBeEJcToSggOb8RIBPWOFeM90EPw5rErWlxF3Z9Bo/ZC0g9VO
xgJnMxiTYRlLLGGB60R+f6I49zhFwjcgsj4f7SpZzZzwsI6dEpP7sOOXoNHlRttAjAvBmHPKgNsO
ENojA2R/GvB/SHe4UZUQi+h8PVBtt6LyxSqn+7y+F2RdslcWugg1XBO38kOTpSLtCDd0DnZ54/Wn
2yu7jGI3GNR5f+CKpbbujjiOSwUCCZfb4oqIqYK0s/blaRP3vfWqBMYMg7QaWDeBahF02Pap5vLG
LWrX2eakdZ+9YIQi3tnlKMXUtiLWzAAT4q2K92iRf5QU/CQBVQ75G27ipxMBhBzJJV6h1Pz2G3eW
LMWQbTGctYBV821AlRaXFKhy3qeDvOkje6qmXbXCkN/iP7HmwrlhbnLhnkGThKqe00YIBkYLZair
2fHwYCJq9MrgGatcGkAmDxqKY8E7WktbPNEG0rISRX/gZ6g9dXVjic4l0K8ceGoJmPUAlGV5x550
KG+HETj1oZxkf/zgNutNQF12XCLRVC7NUpD3V/56tTONlwAXMX/4CW+H0Mr0WYgzdJurPp4w3K/e
09/ZRF1UITxhSA6wWYT+S4nC8mNFMh6RFWtI+bD8hUw/Dli5YonKXMhY6ADczoro6cHxlCeBFxCy
h4quGYuMs3/71qqHwvRzsG/LSRjcycd3QRlJlTFPSIpQT5UUR5vDhKUTLkxilrnCF8uTdztntfZY
0KzmgbcsuR5nTRSWLjeoyR1JB1yZ7Z0HQlnPetwi8CGQn9fbMg502mTgaGB1RDnqUHZono7NxXh9
coRh7hAP7/UyFuOmya/MtQP6izy0s5fnq/ukeNeeJvg/a3ce5zUj4QfZLgKEuvYqeVu8mscvd4RU
C0jmrZC8m60ahv8mlmyVh6YMUMz9PuQfyDPfFTZR3V0E31ESvh7O5wTQPAg3daxpOiwsnOI8H1MG
TK9ox8X4sCb5jDn68cOP7JDzh7RXsmDkJJWpmvDALcUBg9x2HG7A+XgKQWWrVBblL3aSLxxhVwqI
7JVWa4Zv76eNAGdKqIpvYJ8r0sgCYPoGRQXGWk43yopISNMqPIX+hPZ2vKunv0wortZ9dW/bSq4M
FeuRzJ7znHX9HnF8GYYE8QjxBoKUHCS1q4VfB1rNwt0iDEPAXsv0k3m4lpbZxc7G/mdlkHOqn3tx
z//OsW5gfi9z35Ar70xPnt96IkXAmKcEDrQSN85PXGiBCEOJBCE9qF0wJDok3Vrw+0CcqLjZf/Yp
ivixr1PQmiJtgP9cG6RvjoR1amau7OPSFhCCLvJT1Ljkr0hMvbAHExlVsKh2eqYngiqzCvcZIvUS
3SpEn85EJTGBpK+B/9eSoIwuLBdWeHm4vp0+/pJ1NQFdUzUU4ZMA6dg2XjPdO4gybzHRCw01GAzJ
AblDjpzv4DMvsBHfeiEAQytcEwKXAzyuhui9hLv8t7OJXCH0wHoNR95qV2F5imuS8tPosbXMvMVd
A5Sxg6oTfovnzqFRZ11oIbZ/9mlW73e4VcnCwXvk3UuuSSBK7U7diDbQ7h4CFCX9gQq9tb4qqn9J
5/UKVTn0T2YXB9qxXCqofMJrSzie8C/iCUA3b0LDou46J+FDQaLu5y7/Jl3kXih8nnlrBeUE6AYV
gi4ryIGa+Tsz2U5uG5hVroaffI5Xc1FijqJtyYPAlCfBS+JNGN0HkYgdfiPhKQxZ+b/9R+ARSqTA
D7BH3fyVNhtA1zi4OwlyI0SoSO6W5E0l+J3DHi6CfH3no5g8chR2OvyRtofykcb7YL+vE0SOBBmI
N5+GkeOfxP/jtQA4YdJStbNBSLGD8yG74Fd9fE5i2J3DG6Sz/+dzocbeoY/awnWjtbx0wGU68nhQ
vBh8wMtG4QzFYPCXoItj0REc7wD9CJEPGeFP9vxdsyb5Z1dxdOTHQe4jayQJ1zK1IcxFsAgYmas4
70GXKJxWntN+7np1n7fcQJcB/G0nPuyAIPH3aeKkMdRkkNhdGB/gYU0mvPLfWEZONiGQhyvkLLY8
JII00lXmcmVcuNavaVU7K0Rmn91EssLhDoFMlLxhLa6HDU7ZN6dokjYQCd/vi7IqxkDMNi3n9khv
qzsgF869M8hjwDYH+XKyyEekwvmthUK1DJflx8ZZNt8gv5gWKzkJjZ9uf5ge/FiwLFmEL+FkwF9P
MFe+//aPfvfR6FzU+xFmsOuxfBzQrE6FvWspt4Z9Y76oCKMLGppjmaCENKe4SOaD2p5Qd8j2Jzal
NAlOMY+A7/+Pz/TwG/bQ9S7dj/Rx9nxvclTC/wN7gGEBCqHAXBjwaJY0qeRSAbeEdAairW9ieA5Y
9Mrs9CiyPZWhGHFiJ3qhd5WpemUikTangPRH51uMUYxp3ivzkftecDzXmNCXTnzwa6jnHe9Cwf4T
amcZPO87al0+C179h9az/lHu+2WvX/Vr/zUzbWdiA32fJ5ZepJqFXliVZY9M9YTcVlLXPCi4rmZi
41r8yyHPqcajSry7Un380GpzfNsQTUHln68J5el3YibkY3zx+a6+FboaWl+sEozvw+wwmmORpDKR
x0VtxDTBFdiMlNi9I2kz+98LpnaJkHVYjrGDP2U5CKREzKvO5IZe6CJSp1lslGLN2fkPpyqLqLgA
kFPGdDg0fTM6pL7nY5vMANNDaeAuovurNWbyIakTBcqlRBOynIGFPHW9fQhBBrd/OTfrFuNXZDzx
cuZEb4OO3qf2fpBQ568s1rd61VATwmM9b0X2NmtRtRgiOoCqV5EfEwe8fWYjSXeOFRQ8CHVPRqgU
MfR83nj0Iaa/PHMSJtr6cJvA1bnfJYJ5NOdZizc8wtLQDDkb0WGW7JJo6Sfbvf79jp6z4/Cvusb/
xAm3wSzRxzqIuLb9dDb1vsFtsCp79eUedRluh8I/c3nTrD/HPLuR/Pu6aea8+p4UXxe1ipiM3vJP
334ArtQV7FEjaB7af9rFjBWSxOEjC0c/7k+qOQN1qXBSyQlJ7++b/yI9fvrt2jdxEbHp0uCc6a7u
tRxDy5tAq3PAS6xIn1Y5JHbTVBAsq/hVeVU/mr7VN497Mswf3TRFJM7xvFDx7Cq/dQ9D7UeIa6h0
OSDaqTTWxra2SBdqLcjn++ypjaw7Xrtu9lBu8U2BA5rFmungmrnAB+gg3rVllA58RMAcqVgPTAbt
J01EBPPEc3B/Moz8thrH989ixuJH0srS+nWi9JnMb2DPSa8qAUwmzQzokv7DyEonga81EVBUdXxa
xgNk1ODzSf7LG1MKqarpk/OR7AjOUoTpaBpLlxIe887n9mdYCRoahguX0HjkBeMJ+xzwkMX1ZKw1
TKRlSK9tu7aGlPfnZ2cYuWbPL1LspAbreRCo39+GWZuNMCG+2nhQgS9p/MZ/Id10wL/GXXmaKlov
7W2QfWInBwc2+q+Vi5NcutJ6ml8q0Cde+qjmfJJ1a6bNOKKNqtOsABDJyxR+IXx1erV248cs8x84
uww8Kp46wrBTRfOI3Vwakmq9plt8hUY11Su0OSJ9GvsBUch2HIQUFKIuCii5tY8CeBg+YAqxUlRr
LOITbUJFuYfR3tcy3lzUC4ZBaSqP8CyC4IHkilmToWmoODH/YZKqZnemDSGcfWm/XBRg/OkN/3ob
epFLFrlyTbzSeIaj48045daQnerULicQWG6Q1gCLmvxgycMuW4ES79effGfOGMn2hLWYrW0ttm2Z
iPSR/csX/BJ5s9QIlIoOkZY9Y+oeCV0pZI94qXFmmNe4KfnxBaCk3Ucvo3AyMcKxOwmKZ9LSdQgr
59Go0clC5ihCPTjdt3O1ReCpRjqOuoCu1ijYw3HDgEFu7El30JbDdOm9KJVxXiGZN17sAoWEXUsa
DdciNZ4oqBTpeJX+YATGFWHDjgGxpJQvmsLfj62zUBqf+jfALu71gcjrzF4EnjAcsS6HQU40DFbj
LjievMnq+ABM9r0KFuTyJ7ue/Ir+Gzg4iD+esA2mQ7gNLu4KU96jbJf3NVfEJ8hgU+ep7C+YSv37
Oin/ufejxK1wvcyna0XWS4inHr9fNHeANgtiArCgbVJk9zRUTNQhJnqG4C4G73NK4Wr+VCzJntuz
H5IjfRSXgIxSK1syvwluiJQPq4Ejy5Ge8fgfut1UEZgCk0TeRW3xGci6dFs4AiUgvu7t3wyFDlfB
Mq+6UgZOUoUzKOj3ZYp+u/8HFO9/9QAVflOhSj6UxBLTiuDeuVXdO8odcI2ayKQlYoIOZmJbSql7
e6L4Geo9HsCxF3OzETI5xe+dWWmulXsOtkPxBujbYJQvC9sAUaMl3aPlSKuvFzMI9msGW1OTRAA4
lMvSCKv6USBDB+DcjqhB5IXCXGpX2+09HsmRGS3yuvYlQQelgN7VrPTTrS8EyWDjSW6yZqrshGG6
A5Wj48fLR+8g5Pw21PdGWCFPYq1wYQiuruVqkLCZbDQABoe9OO6CauZtyn1rEDjUVvJ8/IoHkC//
5Y/YrqnjXtEg2kEe0c+SoJotaCjnyLME54XQMJZNViebyFwDksWRDFmGFAiovI7LesPjP2WuYU/9
Y4gYh57e9whXhcmlSYudfN7+z4b4V4uldxJLHT8eqcd7zsEajIYIV1Yvdl88nnqsfrr3Rqc86Ueg
3UWxDme/wxzgjxPR/1AtWl1D8pZ1na7xXxUL9v0yiK1tZA4/u49iiZr9n76RBbbAp+4rGySN8tY2
hB5zyi+7a3GNK7INAiKrIexr3o2xgrsGDXfsRgq8NQEgyeK3wLwaXWbf1RwWmZ/968qDKqJOgJK+
qbewhrNa2ypdLRMp6jVPAg7g0IZa8pH+/CocOoZlm8kqQc31fzN6bKp2u/NmfeU6/Krf7K2X8LDf
IBdCw9oQSo97D63OFiApSlrUhRSJ5WVULJYhtUDz6BNtXzsQNTjDp6hdkxohJmkUETa5c7Pjc348
NmEorHviRTK66Me9/+1mnHqNVIbUdg/mW/tRn1D64cgW/7HTktsfCwTm+8+ycCLtshLL+hH5ND9U
85e0R8TN6aRT5yA5D/Rjk/T3f7cw+eA8sh7T3hEVC9HbulsTZdSsK1zw7iXgF7SvcWqIDdbghgcc
Ie4EVV6xX6406A8gzqrSVV5hLQS+lwpqVf4Co0giRJ4xeHBnnXEUMJMaCRLzF1f5YbxEzi7xj93X
EvJk/KzmdllOA7RBSQFzlH4n/HoS4ZQzZ8T/TZGPS3B5rtiCgb+l2B8e7aQOnwZWNxXq13l+t4Lq
wnlaW0sS+8tH9iYgp4BZ6z95YDE/e1GIyUfrykbFYb50jaG12bPCpfenAV/WvCmCWfXvq8v+zR2b
SgsdudG4XFNHUQ4CejGw0qDeOQYFVQ0k86Q1qId9BSPl+L36ft6PldU3pUZFnL7z/jlYjp9Wq1jv
KvEqYsJJ8/L1qeJB6BG5NGGxbUerBiKXYxkPWWKpKnJQSxfbBNvifemUZhwTTYWw/iH+totZxYXB
HSNPtnfY6+wCxlzdG5JoTslLVsEUdBjhUSP45tbMDAB0tZboY6DLmhbZrKPxUwVxBwoJYpyIioCr
agq9rqblURJKm6Ywf96bxt4HVeKE/2mmwUuttzvpyp7OXD5kxE7wVkjrX/O1tLZwXgB2LuVzmwjH
OOOamkLdJO7Y+UACj2YDNsj7HDv5vwxFT+I1fBiaFx8S0EzYm3oG/+J1m+AhU4O1i6yyzMOGkpuq
Hh+mQHJ2ASzQdxbPuAq/e2h4GzJnpHUN1HsZwC/0QG2NtjzebnP4THVjR0Uw6t29OHAdxOq21px7
MkuPm0+qB2coS7o5LZgnS0THlCk/r/vtF85UTP/hS23/cEr7uWKQWUZGL7x2j4JLm+CdktOYsuzv
twBiIvwtbc+6XtSFdsi64MpDnF/nAAA8pTmNkaOX5n1EFXwU33Fypl35sRAATfcWnkCotD1Whmfp
k2zCqTIj+gxj+Dx0ws7InP542lsf5Kwthkw28OMLD67eApYxKHmJL0XOa92CLKVKKikjRvCWt68K
zQ1PaKk9d8TXpI0yIgjd5To+6VGwtn7rrQPiScWuniFYBzPhpIgBn3ZI6queSj32und4cZ4kl2FB
i9Q1eD6DScCrsoMSUzAGhm2aEWJruq9Jz1iWJOwBRjoGTrBaAqzR50VMIQY+crUYkk3cvCut82z7
ZMo4zG/IwZbVOImp0O4UdiKEjIuVtPnZkGO4SXqG/xTVN0OpzpxRSUwoFUEzf4csNeykYEQH2ek2
y7Ki4YZiGZy2ULH9+qv1RRgqhsoDKH4/g97DUtgfkgeHwz4SHfS8RAIQ4NZrM5ZCrUKxj2apyRJa
UrSMIeyjIRTAxYie8OK7H7DPtow6QzT4UCDDtz8H6i/elNN/fJzsiBYG3LqhujpuQPikrOCvmCfr
vTsR/R70sIUxTnTy+cAOzkJOXTDQpCHnHGaCgY6hQh/mFf9mRVHKx/5czgjBcfAC2GF+zWWZNxax
rHzlKLD9SSnzRJVgbsMwBlfx2QreaEqYlFktt9U5F1Tv/9LqASYOrRn45lD2sU95u1IvcRboHrxl
0qx3pVcYLW5k/8rmWeHc2FVCRaYlqV0JuzbxwlnhBLWuh2SZlliCu30RAAaKQuYRQ12qmQ5UAyVF
UNVQluaNbQZyMOHEmbGmEBnQ7DuShoihZ7+jID58UxDMOax+px5fMXwaN9ErG8/++pdrmAUTAA6n
prTxzjhCiNR6Xtu8jcq+kStZXmWnEm5Mnf7LeSN+ZAGyGBLu0yM+hagUkoUVZu7K1vjMB/wLn7Br
CXj+ccNQEnY1FzeF5/sfHozyYL/MmPItvb6fVokqN+dASC+s6qQhCbOMEHoidIeicUQ1YYyVf8yI
TJoaRfGUE1lo3BCp5ytDPO1/TSZmyvVQM1VUM7sx3+2zqri837W22C/RTlikpu9uUAwGZIb5YYNV
2eToj1QeOCw1SaxbYgJD7oEdEtDmKU4EqMdAYPW4ZeP+L3zZGvfzsG850VYouj1pIPa2bVOpAzEg
OYFE67mKGbGAPxnLB0KZEQsYUQadVLr6NPgMcSxsS2VZd/2GxhTyRV2ZQHqrhcBCjwe+G009NAym
baF1ZCGiEDPr3F/fIndU255c4Wq6nsKuxWVrl+DVvGUD5NsWgkFVB2ixL3BcBLrfpMyQSrsqG00G
K6Ba7Tg+KyRQDLrNlRJkvQUN5GQXNnDIzRTGorOgOUi95AuNLUFLPukPYLFWIVnFf4dQA+B4VAkz
V3lRiw+XKaGtepnrsWHCUzsQSXBaS40tllwRIUJjo6SVuoaHwlUs4eNnqK3UF8NHrRDoNZhf7XsF
U1eOswSGVACbDMixN6k1o8Q/J/RGAZOWZMWpbzlDKqa+V0EkpMVDdqJEGjF5qDZyBSiXm9uULR2Q
sWuTcu5YsJkItrh2+KIO3BlDErRV/TCNMTH4I4H4b3UmFc+NZ6wbjApPq9yJewaP1L9iPQoMONm3
YWGG51fewxPcB9Ku9wd7WS265U4bz60nWRmgmeZiEkOv0GMXwYeKHp7Bn0f4V7lOPW6ehDs0gMip
B+f7nNvvFVpgmBE5pmHMd5ls1sN+Eq2NE9oh2F+ZHM6nJy4WvwZbaLqJOj+Gfys8ZpAChNGDDWtu
0rlNkBOh9wOA3YwyINh5a9rPayGEuaehOIoLGAwyFFu5oPgwc3k4jIUeD/TDm0Bt8jwWDVmhDkFo
MNMaJ88h7O/Mx1m7TgJDnHYYwXk/mWA6bGWdA3UgrDpEWtq+UUTQH99tqCV5mws5nExeSh73vC/0
s8aApZhhGpixDcoM9OJufqNIvrQDVC3Nf4HXA1VwSlAhtFMzXWrzBnyfGe4OWvzbBUihcQ7gayYr
JPFSoUOptIbKxr4TCCqhR8oGVoXjRpspeWKLe1AjGx5gyIoQlQ4mtx0QVK6luBrajpZeP9STYS4h
L/izGCVn8deDV/qvjKnL6TwM6ybvys9Hc8lGufZMpkHKH5WmQ2RifZrZn80xjr5UR0WOnPWdDpfh
92fTGjNIs0UeDf11b17TrspQuPiw/VhzAApibBGhq8J3mxyqYivTs5eawIYg0l823wdLcpdCyfBf
kgZbsnWXYftAfuqzDH+TEh14fSbpThdt/ycWvZ0wEsgSdtSyFYsBdNREjRAtS3Lr6HbrvCA7TX1W
sz0EziyQVWVtW/1MKTQC3F7LL7pUs7njbtLtbPSyXuTF720wKMIcC1lGKe76xLDOmyshzjcemFjJ
6f/u9r22iTuqpDisHRrOv7J1la1rA5Bo6Y8H49SWOXN3j/iw/+btjgzV0LYn4M99DUN7Sy6qKAaV
I3AfS4AkuzKDJc7AMQIY+nCcbJ+cmB2fbrVDt1laidu5Fsx5OR6TJ7Va7b74rfO5SoDtQ25nAcDp
IpxgoSlCLr4jxXZ1V7nfz/YvscmIhbnsB4xV8K/QUHplPeTzPNVYVMelEQwpVYtTdi7BgdoNcjc9
sOTT0mH/Qi0Mx9gDGY2kSM1/Wnh+7ZsR/uPNL0I85HNi9Qb0SL7SWCCoY0AjCDF5JRy8ErMxU2iM
7QgJKXgWNazNwC7Xn7XwssATzyUf6IDpcwxLgNYmKVWHsN4LJ7dn2G3qxMpx2bX9IumXVmNZrMGJ
Mh9kImMeWrKEoQ/SyF/1onvvrFIPO5+vnFO35TaMhHwU5oSyMeV/TuruZ5YHa6zoammvseOFKgCb
/JQbUGTB7GzTd9L582Ay7WfGQ2hkAgPPb4lRoLG2J9MV92oxTdLlY32AsvgAYUk0Vxz9uUXhlQT/
gV7JQPDCcgbu+dOcnMwUu1bREv0nVawx12CPPXIqfW4DzJNje1KVza1jneYPykJ4jAHZnbCDzLCw
Li0KFz0TLd4zsibBZVXNjxNzR1yFQEjEHoexe9cIRY5Gp4d1ewrwLyoulOx4EnWuFjUXdFyIbrqz
mYNWbp4jlxzqA1ig8BGZMYRxxyLwJ9BJLw08+pbViW8BA0jnpv3dT+I+d/SUgbg16dn54nJ6/yzS
BdtfFNZe5ebNSDM3PlB2sSvYD+kKiwDAGBmG5AsEzrtKup0r3kCwgXY0BnP48qf3Im4O3WDAcpMG
LwBHbKgcHQcAcYlloHQbHW5gsVjNyUNL5UQNQKZZ6U3nEc8dBKcXMDZvsMUrCPCR/NJShN4S/Wnk
M6MxQU2O4Z2HHK+GJgayKhSMtsJKtg2qop7o1beOBUOfv00MTM2uTK7av2O64QjKKQGIDMG/9bs9
9UG4AcPyOt6H7BkL77ONEmMXKW8k9/Tj4AzsA1pSw5W8Y4IC1fiFIftYisfyptHeZDWasT+VZhr9
u7SX8/jHntWsugQoXydb0ZHUnN/x+fMbxfkznSebTI7q+qmJBjcHaCjZjel3WBaGkwGSTXjFOT+b
tsKRtR2RdDdhLOztNU1VAy5NjLDpKhLj8x/N3XB2dnip9OUJbxjWzurSy3ElqC+bivS33WmF9Dl5
mOhEPPZQtBC6FqcyoD6vQ1i407hFypSrdUMhjxehwXKM6c52tMJ8WEK6k4B/VqUjprLELR82wmMY
H6VaGrLlRtvqGcrNiHztrO6WSpiAQrmqwRhZNcRpbd7moQm0Aa4F7XTyYjJ60CNDcIDlVbrnY/md
Q9Mq9U9h+q0n/agK1aS1A31JZEcMrmqEAh7W22z2eFvhgPbaVXAr5wZikz/e7ZqdcoZNNzZla4ir
qUygzbZeV3JLEzAzmHelLpKqGNGy4HmOE7aGQqz1jPMLsRUngjL9LfNAdiHs9nRsFjWkThEy4gyj
7rSw0LpVLv+FSIjaDZD0y4WomdqgYCyQ/Iq8rvv4WfGf7LhFpSwtY+rq+iNK8T8q1+Qwcg5mJHYA
sZviBGZdJQvwAft7IPQn+fWV2YjcHq6pHkH6UYRJkwnZHssPa7DREGIc10FHtXGAMFvgY8LWTIAy
pyaIeOOQs0V6IoEXKb4guGO23JiuCgqiLuDESuKHu3dR7/dcFaBVqRT4kQPEtJs+kjm7iWWzQUZn
1q+TmZM4SM7aC+HX2AUv2cFkeLRtTylcnvylqdwUhWl81ykDXxpQDwVO1xPhQr+LayWnPVeKd6Qq
Wzt3j9AVxXzB00Stqg2DeKkVVV8YeriKP7sYhKiqoGixQ9I+EDn2qCUtX3QsvhMh6j5LvIs6gSXM
JYHehSo6wxy3w0YQqAFMaQAIc/PmYgx1UmEXtOMG7sGcapkN/rLpQeYKbxXuRp9m+i1q2jk2mXdM
Qki6CsJESZkG5XL0i4I2ed0q4Z4Bkxg0BUEJotmkVH6jt5Dur6rOFVS+D5c58f2Yvcqu1gX/M+BL
SPhImrriwut52Uy4B4pd75WB5gqwFh/ZN2cJ4Xhr4y22EgctrlGisgDOPSNQ8IODtk1MOUx3L5Ny
jeG795Pl0LHgtEr0iWkauQCX2lAZTQTY9F+n7y+kZVQ/DRRlKk/a7/WNy5ONCe7qUqONj3yqVRCm
AdooBDdJB+c8FxMyWxx/rWD226Gw/226YYs8C+ZPQuchlzGaGCyoyMxvSZg2hx68byld6MA/5PZb
bzsxupk3HncuNes+7s/p/40hkLUHoAzOnrQvs77Xm2hREVMaj6ZcE7VJfMr7VzLNpkb4lurWI/Y1
BWf5mKiZw6IEBSdcNGZYdQYQxs3q9sc1jPqhC6QKMleO+NLbijoauwjjXROVXB2PUor2CuTUcxw1
/vTetfnzZZd//GKl3u1oS63weJ44c5Hfe8LEQm8F+jO5fJT7MUpb0+5rdgVFIiH4nisWejCnSZKH
dQEJSKC0IVBw6QTuV38xlsGDuRuNccaiE5iC9DIWQ4GFbP+45ccwt+l0dpWhgT8bM5DgYTPNO1Hr
nRJdIaU0SjfEMlC8sRnsrQ8PI+I7xBW8Aeme+mk1CBQLTEbBwL2mhlbooDfmGuSgMip6Bc4ogF8Z
vWxRyKRfpEh6Uu4WPgV2IbYRwRwaaUXkTqM6FCwQGUS+jsxh5CblaCpi1y3m1flDLJsORheSWqUQ
G3A1L1gGRb3Duk0Tsv7q6+E3RvjBdcYJuR/nY2Nb/RJfWF1XP9mT/Q354prc4k21ehk9GkOu1HLu
F6IVO+880LqRLH7Zf8i7rZmzfbVZ2Z55kL6t5Z+Ip2SRltEu4QSFgcowa1N3gJ3AgEixT9ZVxBxj
ASPXlgiX0G0y45eAbxWBBf7BxrsTRycIu8yFAGPuaNn5sIaLByS5ib3Qrfob6Tt8Mr0gzsQKgcjS
HNf7Vm4RS/ySKDu0minyA8k5n/mbwKkfhY5vd5lWZvHpm9WLWXVe7yKFVy/xJoSMMzXVHprh3fnZ
i9nIRp7nI2f7FgBILsxo3av1M80+ZH8PRF7Kyl54AFBnhaVqpm90o90RJMozK33n4Pj7YqoqnOqH
9USppfyvqK21LLEZkvhq0NPe+c141EZxhF/J/lZWsezmqC/1S+DWDl+k8H+OR1PKFHIzPfU7EweS
StAjGmysmKmBwpMUHww2/kOqHfEYhNtmn21xryRiXJzJRJfwNPqPsK5jGOTbUKaCEd5ILHTUv4De
gJj8ayjJmN4vA9avxB+k5YiWKFWu92ggec35xQiqZSXvS3g5cDU108kKOw5jyK0XH0No6er9yNY8
G2IBzN6QpLntTyQtdLauiPdcaCDj6SCzcZNgn7QydR2HSUBXaYTAd1ttdUMibR0RQbPb7bJUav5x
UGuqlRRfbNsme1wGIXPCUDfkEyo/FFfssI6RkpuNuF1H6MkvRWvJLJpTX0M50fQEHgfwPdyc76w8
QZeDox2Iv/LCd2CXK/v8Od/XLnMdH/VGqmRBKflBviVrJ/gEAWCEBSTAPhFFXArrOB5p4+4ptnPl
jMu0Rdk6F1hw97okIZq7qgaoCJmNfKLkVyu7nVwnMCB3ZFXByYDdH3ZUWPITQUXXfmxsE7yAxucT
fr97F0u3dGPu/HPBTiRv5lhI9o93jV3T+hOxE2yM4pKHope83NenAwl5XX4kmwPgaiH/DrZvqdeA
EvCl4RiqU9jLFMv7TGcPaPA0fDYK4MV7m7c1ElMGyTxQrVkYDiMMAk/Mi0+6laWPHbeOg3zQdbgL
h7T5NP5HVdIKGfN9AFzGREF3A3kkUgAVqSB5XJXqmPUr+lPcIbNCxIAy7yf/s736It0Hlj002+hv
aJx1bEUGZPYgOXJzNjBO0UjXE9asbKsde6pyaRnJQPN2yMpp7C/ClpNGyRbJ3Dc+iD4WhEo2+/5M
RmukqNe7MgV7m5NeSfPvx3godCNyYyYIneiV4nrtntDPo6zUMPzjQHMz3/BGGi1hv6DW/HVFYg5q
3ytX5iw2Mqw4JnUVMfs7nEZI/cGZ1egacgYdoLlgPsXwE3oLivYr5x27J8S09x25zlTcW++O293A
T1/XhyWE/FxCYa53mMuMnSqeSUL+uUwFE/6yUpiCGM8OVDGYBY1BnkC2OOQ15Au/Bcb5ryGlRdRZ
NqxS0wujpTaWrJsWzo5CTiw33JPOHl6piZmt3UGoOdaMxcseL8lEy+zfYkPcdqP+V1Pdi9sYSi3U
YJUotvQRKbECswk7FL7MAjQcbb1NmA4W7Nsm+Px2JT9kxtq2NHe5Zo10I7Bt5ZiuSvGXt0x5q6Lf
YucBXykx/4PsTw77glAdO7wRH4S9aRsTp4JhIk2FJIVoykqE5UPvAB0q3kxieKs4TaJAfPkO4aUh
eIcn8sGoifHu0sxIaAqbCMzpekTvmm/QJPhotsvLBYQKiJyE8zLxSl6kc/03N30uc3JFw1QPPovS
qE2wedgx8wi1zBpl/xPSCRGL4QdjsOnuZecTIk8O0GMtlUQgYoBM1L5EIXJ8arqzouNbSaxUo/4y
E/bSBPOZFVA2HcsicImtoXdDlwZYiugyvWBevMwpeT+XUqXrvdP5MKThRe+C/Tiif3nE2ky5+X+a
KqTlBB/I2/77axSdL4XQcvbZEiT+/aRqNoYPfgezrr6GOAWb7pCotmCPZtc5MYTo/yaz2e3ZTWf7
CnedkHm2vEB7Uu3L5rZMAYCFSO58CEKTP7ABAN6qJbDG/oSDCrXtS+/sC2zU7+5nT4KqC9TdxAv8
UfqvCMKRGTHQIGR2WlMWV388zC07+jPaDWN8mp0efgePueg34T5v9fxSZPKS+1CDDkQ0q+4zvu/T
EVpYAdH39KJB1gQ3e8efYQ2HCAo1VDXhimw5qJDJda4LZAstVQKfGlFT1/Hc69By8WS5ysNNcUNo
/aQKT7GOY1A33mkuYs+p1cp5nF8o/kuaiKppQbacUM/MX4VASiph4QNx31GsCLpcdiCwLapZEBOz
wv7kpLDrqcOV8mmfUJxms4gb7g3B45nq1bqsd6ocJaIJ8/oi2jD+1BsLT8ykVqmhvW3OrglPEztw
jHIzCjsT8Z1dKjcmQXy/5N+a7GA37lnuq7GD1wSNfD82Dq03jl3eMtCrKHmIzaHmHElTuu0si/uJ
QOK2riF14rRYBcJ1cFaXjb1tU5Shnm2YHhar5wRew7CGHLVuBvP7E0PeNYZ8psz6PHD9PP0fuADS
uH/IUgvlTt4iVcI52aryiPowhtWUWfbEufLmWZNifnVwd0HaL83R+b5Asw9RZVtP2XiJE++T1BVA
ySmSqqdk6zTmVvQBi/aEROxxntVe468q88xNTqstzePMKOjmZSHKsL6cTebSL/WJ4wxtPcnsWTGN
kSFYrRkr89/5e5IAru0F4/2p+9r9n08x14l49xZ+Vil46C+OvP0LyxgErQy5I/C6N2PYyfgG2QJT
hl0KMn9wkJVwpPWVkVAKhZXt6Z5cEo5OS/s6SG8l9t80PM3Buq1oTCYSAFVmnLcBTuzlDskol0b/
7diK/iWzXrg0n8ja1DekPqfL5Uzu1WAtUVm6kXC8XRsKKiPNaHZGqWwlz8i+GHZj/KGJIqb9OrYv
3T5EzYQvKYxZMiM9+6/Gt0uCGK9LK5osgd6lSGymVdYAGim4MwPD6RFdertLEpbCRSosZ4Ocre7g
kNZeQ5stfUDEGMFP2IXJ5o7qyqFWtTbi0FFi9TnYkLDbEVdqWMssUeHmurwR2NxBHzhRYQYoatKV
9jxppMjU/ujeGsvzxOsbocpyDyqKAwS1MXa6owEhc5tQ8nEvEWPU9Wjd6J4El59ZnkE1RlaApmAs
Hpd/Ax0uTpfKVHVECZAsVYe6vDJEWeMIG3d+YtRsfPzztdatH6ehPANFGIgJSVJwgWEsG5jecqDG
iXLIQrYtORYTyats43JAEfj8JqZ199L8x+b+2ev+4TAbHuo9g6gsiF/1ZCXB/aHK+xxcBJMJ0Qym
Gcwn1o6L2dbDASvqMKrQ6DMnEJb7/8uujpWuaGEAiUbRd0CeqzO/S0qlk3DnlUEHEUZLf/Ro2Nrj
uYAcXsDMMkdRRhuPBWn7sy3t0PSffr6iKwQATjwUcQlmctNjwlHfaoGsCrl6S/aJ4drT5/fbb1IU
iguIGBCwbzjYp1IY76yuXEcvr1JNSZBpGWZ6A7IblY8zYoeMwh4UYj10xnZMIv3yPJedjJQTaPzh
Zplgu8HiJJmw7eVqaKAyJ04JzkZz4wQ7/P3xCQ+nEEaofVCBZsk3YCh/qXFSccs3mE1S33QR5jnb
8JStP/sIiZBsKoXDSVGsZZsFhR7eeGlnSEt/9PBIHXo2Ig0Bndm0b5ziAjUWC0dPQOSl6Q/iiXMq
yoW6kb6VyavuMaaPT6l7U00Ssmn4gX8Yty6ghx9ZXucvZkSi4JAWf1AuV01wPxoW0IQml0PyUDrx
z8ZDY613N3uGUPKwIpBYw0XRXeZjWizAZtEvQ5So5N9WKsYJ8QDUouvZDBSldFNCmdUig2De68t6
AGhr1NZy68dT6VTYu4IdLyglSv0ICGBUHezc5o+DkKnoOIQqivm5Q+fGLSWdz050ZiV88n9vQDGu
FP+nzkt+xDqNWea+sDc4XL4/6St00BClkLxfA7ZxRKLGyzz8rmLtemDZJ9eMu839YGBjO3ErPqM6
M94a8B5H5HDsBfxlFvcyDKVoZaTRpRLh0Mkx6Kb6RQK3+JmOkfblHu3fnruQEXi6J5GXdqsNTXh0
9w3iePWlUJDTYcig2tQFuM8AqxaQ2CS9gAWQKDi/XZgeGuZ2B2Un62XLRqPGArDttYVfyRptoG/v
rKbn9DjWAqI+wbaLhF2OZt11nOgElaoxsKUpCC8rqOywiP3CVODPr00a+jwJxooFGyuyGMrv/h+k
BeMxK/MUJgwLex0tIEKogcxBfWC4QEPREGGiuS9Uze/pXx2+9NYjTRPk3ikjWszh8GZ5mklZjDDV
RK+Ap4RP7yWs+yTmTKfQPWXnin/5AapOmg0jveK/AL4VECn5gkpYecdZVnfhZV5efuhkhQ90l934
5WC9pvJf/eyd2JiamXLW36AC0xL8wpQbCf0QGTULWQKov96+PatuZU05aYbrbqrJOVfNpRurgTXf
qG9dvA3KAPxqXfz1oVZnMRnmjydilBf1wWYr3hmu4BctR9sEMH4b7IM8z0BOpVwbXNzby/Yya9cH
6LYmONhKP9sbQiCjQvY7W3bev466C5xHGhduJ0fqJiqGoFaZ0RRHS76BXtC3r09BEusby2QCt3zW
0ZATL8AYFZmtOi2nyiwi1O0HOLkvyAzQe84RsdEiaTCdhf6ZIZdWrWQxfOh+vUVMGh92q4mePP3e
qdduN5gxIbOYRD/+uGzBS6rzKJrciFvda4EQ+aLKUDRjMR+D01ihxXHTR35iLpUVgW6ru7Vxc0et
1utQiq+JcB0jC9qBpu0VTLLiDfrwmOKA3heC5dLI3ggqOMGxxw2g43CD1P+6nGfoSEVJDwq3afZ8
Uge+wvkB3iUJhqGwR7DNjI5wzRUlu4w/Q4DD/33mZAyLZjMbnr/lfwHz2cCwBFd2kLy6B2BVSdd9
tv9ENVpz9fMJRs5UXiTQGQv1YBGGoTZ0rOX1CY12HkD5q8NC2B9j5PQax5ch8ET+iX0RlYuTAlo3
TwZR3DBxblLm42KYRL16cZUP4SdOEUTQbMKGcLy3/oQSrgXG6oTKgLr+O8TEVXsxgFHx4JmnuoMu
wTvGEp6laCcMUgN3J9UPHL0GkMDPL5jwW27FeBJMEcEuL4xgv7grHW7URcvBcx9rzAC97mEMMkaF
wVLACYjxNV2oj90aK75aPqZSj3YoROrJlDNEPTrS+A4si8NAFI5fDIGi/wT/1edIKdBcJP1GDks9
FswpyxFasTs0lSOJoCtduBMshL03a7D3vNEXYRWS/QOTXw67jZIT3JXPT1QxxEOTRXVAAmFyGhTi
QIfqVmK0MCviss84ZFmJ+8R0h4rXK6svijyslKkCh6QL6ybecl8CKMmmxFI+3Wox3QckXJC3vwUR
8XPWUjbu0yBh8eQtgmpdblqA/z/05ZOlGUQTK1bN/qjMUy/UIrOa9R7BBh4l5I647ui6S/mqPfcg
UDc7T2bFgOkNSwEW+PUvXRIfoAHUP+iB+l0GYB4huiWMKQNYliWCcFpi4o/FYmXKtwhw2/CLbb29
hDUkRZKv8q+q/xXKZqfeSQoSdKNX2kF7vEFyMAhRpLX95CXN6gG7pFfR/IxfX+HRfhrr472PfRXe
jZ8ueAV5Iz20fDX6KqbK789sKliC/rfu+NVRmzfIwD22Q3D/k7JH+w+hUYCivglKHSwrUCAazlpA
SqAFhawaHJBhqn/BqcyyxrkEON+9LJr8Bl7zoZxdLx9TzDk0MEpCbDOn0iilsicY1viXgzQMk7JC
HFswAogs37RfEF4rmDkXskEndywyY7R+S9hch2ZXGwS3r8tepCuBcddWyVSLhcjz+Hs8p4npWdG3
ry5DbHbu5v6Ro4wKBcx+i/eJaNc6zEQSywnLJABRvlOmQATO3uzdyzwPl+OG0s4g9gSiyjZlBVkg
UN/a+GLxjA13HXL2z9wsYJBHyx6Ebu5nGbtYM4p84ywU5cEZk338wX9GBxfcx87AhjKIhVAYGSss
ONtiTH6jCYTW3x8YnorXXmgo2+Pv1gPobzs7AyIkO9qzhIvUTbksCrp0tD27BjaI6/klaN01WmBX
IIY4jmVZWZJzPttiZAVXtz+lQUfHqe5mfyjAdqpBZyf37Xx0EBOWeuPJYfY30QioFgvJuvsgA/mX
0L0XIGpEphA7+AJHv4HxSVtYzjbkoDdWqEQ7QMDHSWCCESw6HhEO5m0NDgWx7MV/+HJ0CGRlQUMn
A5PUsSA8iQy3OjBLII5Q9PPHKhIxVeyQN/ANP88Qkm/Us5AsnGZh/fxRMj/j8nehAlqkdktTyRCc
7VCxXHEGot1nVwWBqVlD2nEN2dGqJ833zLSchjl0+rYRtA5KMFTOaOr68A8SR1LmebQ58Bnhtags
usfYCsgiYNj7geDiLZQlIHuVyXX9RMgW+CR/WoauwV6ROrXqZuA1Lkfcb37KJDstXWD3deeaGmqR
Zad5sGe8j+KsoB+FY/ZhLjtswsQ0Oy/if1JxDoovUoNceYn+ZbsDIUyOy0PQU80Ih+JAyCI3DgYR
nKvEmxh+GQyx2LBYY9crJO+GaX13agabcHYzYSeKUmif9178m9R1Wda//dqCdrNu5alTR5eN25uT
NmCwv6jcFlHdQJll+pEDgZwCFFeUCBok207UKND/nnUc+JX/M05CPeztsTGyq+iYw2JqKKxWw2Vi
ZeOAvcoKkISzXwqO6gFiBaB65QgUG5eQkhvrEWI7Koh7on9xJ0FENpCJtfyadwwoyFE32vBR4qOo
n+uMNtTygfGl00WTeiJwKkgWz6mv2qEiPlXbZCoa4sYmN5iX/UK70w8P1lmkhcaoLy3LSEoY4r60
FXuWFKCa4ZpnoHzUUJKWxrLsYAZ/h/OUDmQ1CGVTCE9i2XPFbEvzl7ErMSi+ifsvLZZ/zlFWHidG
5GG2PVVixk5J/v27FMxiytTfAybJd42PpARRvvEPGjHCUckP8RcbSYH5mznps+kiUKN9Yia91Azv
8dAHWT5AEhmJVWfxjbJXmOZZJSAszLeaTRcKjjezDtmXnvA1BrGigXHQCIHS/zMTpjxpoBCNs+w1
6r9pxicgSBeYnnJjUauEQDK6A4T2D5tRXbysD6grSrBnVIXSAYBc+7txxbRQz3+VKBaD3DtniEw4
D87mfj020cAzMlGQ+ULoHVW8SsABb2/eT5g5DTfV6EuwL6rfAqYLjKD9dYZbxtABXd3eplhVc4lk
yZnWOSna0FJz7z2mLw1//GLUJYD4lUvy7TOG+otReoUQyFylEPsfM9F0/4/c3T5M4yUrgMRlXomv
2ryDC3vnk25tGySVyabbKEQ7YFWYEplImI6n2QFYsXPOj4sRzk2WhloJzlH6NmfWyWpoNB/TFt95
uNL4tn+T6ZbvYozJ5ZVm3Fxc9rC29Xer220Jv+9cUDgVwySS43+Lq4n2P0jW6/UYfqzlIF9ikYWU
Q8s3MBS2qxCJhFYl/3hdyq6JWJBVdsBSnnDjR4BLmMf/XIbG3fxsxbKXyIuvUJ1wjyEHvCn/8XqL
iX2kwlYXV92i3sECZmnZ6uDw7tgXJOFNWTR8sqXBKp5JmXxXk2hfKGB2srtgXzC4xBiwwRNYySOf
A81glxcTwC1tIf049/F58E8YtGcJ4+gRATDAdKPGO+sxqVgBVGUE0Hj3N8EkCde3SOUMCPx9hFta
nRxr69/OhWxBhoTzL6E/WUkCaWLQir8hFe0TcT1+E7oo379/EdnJ+sWBDUhK0BIzBDGkR2HKCN12
meDqfQ+ypZoqAkzhk8ltlDC7rjdaAVzjFM8oSBVMpWRHQUua7tYSnS0bDnVUWEAZiAfmJ+f0e3tH
NUzxT6xNH0HT6e3l6Jx+zLEZ7UgvDZ1i0IAmhDsrAWzNH88CjoKs6yadRk1GkfrPofvN4xyyyPTG
u7KvZHFQXhokVLHRv2Fm/6U8/ECQmnug8bYDtxjJ8tL2INQHZHTcd58s29rpB/Xo0h+NXd7cRR7G
iWIwFLDWYHp0Ag8IDolzde/hlpmIQKwVr3FtJL0FaXcgK06w7BnjOsBrph3etYPbx7fHXuuakRrV
OpUW0VqcyPoZl5ItBmeZ2WhQMklLR5utf4lbpbcIveIxeelgFHHU6DrFaIEXuUGmkvikA4hwsxqm
KpTVug/VIM5HMIVGzDZ/8y1nlburocu/ybV6deVFiD4y2GMlrEQvp0fGHZY0YhC5+XUywdYFfzOf
dWhAyPOP3hTX0SD3vNb9dNmu2Nx7KG94VkAXZuWbAB1IhW2dUAexYFyKHxyjIQBNZTD3ZrAUxCu5
xnwXr7cTNj9K/XoJMfGzk1utX7gp1mizoJe7BN6RsqoB2gDxDA2zTPDkCMYwS70n/sLACEa7uyaL
2OCt85G21Z7hIJN6dwCUob95KkmeyN3cbAMBC0qbRjFXhDb8faQI3VWJ4zUMoWRZAJjQqBdRb7i2
iioCRfor4Q7QUYqQY8bTDCXmM6kGY0RH+uTKdgTkxxBcfvW8pjs6udlWn/wY812PkI0dBAKaVF6p
VVwZLFcf1HHQBQ+XXuXG944j9S1oCEohkQHJJhdxLW9jkdIm/OMN2W8FBeKPFyNIP32dYwYdMx8Y
NtuYTfPZMauvMsQQ7ygMrugtsYYlejuX3HUdljwK88unwwnF9SBasZ5Hxjt2WypTzxXGS0U4+jmS
hHFdnMntiVNpDBb3XSOCIP73u4rbUfrJjR1oWZB5B00v45VAMxB8DoGcPLhj7t9D7wienZH/2dNk
XciVMlqDSW5kW9ePvzMVyNI5cAKmexnuOllSpnAG/Vnrf/eea4ODsd3pSAluV6LSntRy4OxZUXy8
yy8AeBglxG3B+OZtBbgVO2olNut6dG03qqEeRdZWlXacZIF2WDCwoUZ/7C//n4q3zjglmKZhfgdt
gXHyVXBLABeQc0JJqKBCoqQe5DBXpFxesNY7v/PQ90hzZAznRelMs9G+FeX++xOOUBQTibqFU9Wg
VENu3bcBnuq30Zhx4E8S5e4tN1QJEzAikC7ppYgy0KZABZVPc73EbL5RimoLJwmfOlvuw1Dhly7Q
xN4J5f7pyzTm9b1iRJjfQ42uIbpSpajehnITAslQFxX9cSD39kiOGYCx3eY5orEDrD7vmie33tWd
4ly5QdZtLXVws16a1BpIVmwcyit6IVjpgMPI7iwhHa4ujP3HJUNrg2SaLqSdIdzlZ/2iLzI27ye9
YWRMDVQPujlk78EqhL5VgAfUhOQ6MD1g0kL+rXejDIvNP7k9NHXabKlMd9rfEUhnRER6EyrntLFk
N721osgnCjq4Zw1d2ZXgFqYdcEPBZBAxU79AlnHJGwOzcxy0BlqAHimnxXVCLJ9ri3f2zgM7Awi5
Jr9EcxvtIN7tOWkCSamIfnb01ddIEEfMmtRCRFs7LG+FIY43nKGQpZbT/lVvHoPv2JKiIUD/0zli
/QIqG45A41NZXw8wW/E2n/5mPzYRLjyCle3FDX2V+wmrqVIlWycf9fHPl4Ynmsbgo6XRv1g7s/GZ
AruSJgEYezO2fldCRytqF97RBYYjiOypXr5Sbe0Ghi4X6ttQ9ELLRAOxASVMwXDs30miw3GJbAo5
2cgrxBetMMTPBFnv7C629LunNjhr7CUL+Ombil0ZZ87ExbJ8zK6HTS4XefFICmcBEbaGwyumqRO2
AcB0Mkv8IW1PUszHlXxGfODUmD6F4iWOQ+jI/wH3qyyoM/2JQv1dh97WyBsJtpk1IQfrTz20tMG+
VTEFWqyB5bOTd/lGDJ9yZTXroxZERgnir/XaPLGqwBSfVyJZg+BmgjHq1A9IFtsXf7Owbn+spWU0
8FMbfJQck9yQ5/MVHpoqjZjug7KUbSYwmSID0+pjSqUcCx9Fd4O1lhYkYrIkwhSHf9Xb8O9KfkEa
Bps/RcOPFx/chdcyyvVt4YZMLvXMcYpm5mjYU7ydKs55ZrhoIotiyZS7voG4IlAhYnmJuEJWeBY0
9JxAxGu1QxYjFdSTlnIDFk3tUnieClr/8l21jWAVPjGPDEz3Rm6pHXUkzEViEfi37DGQAF7hpRWu
VdAkoN/8dVYJnFs/HEMdJF8rqhhKz8nBqOvgn7Pe5xuA4/d8Jm1li2bhfzU4uFH1KviGPJky4M5a
GQ17Kg4JW3HcTJY0n/JKmdwecBMRuRtCRXG/rXUco+xko0WjlWEJPjXajGBAnCCQVHnmD0ClciAR
2IB+vyQpBLl5VBXkVYtpBby44stbmCS72x4nWnh1GvyAUwILkRBa9E3RavDU5+kCvYYNpk7r4STe
+YDsRk4KXPC/BH1xZWoY7mgyEAnH/NBPM1F7vjojEm9vwX9Uv66xfRmI8NeNamDmlKTo83W+3kUO
Y407ritl6h8jhjZC80tYHc1Aamlv46iRB9YM47wqKWKSqoZThSQtb6hBgBApbyn5Y3niMfGMFxTf
FiPYjDMVvQJGruqgo1hASpJFzJ7eX1edrDCZ9NQp3NanLMXPVVVo7e/1Qn3U9Gk9ulATSqpqJVd3
uvK4x0fOwJF0e0tdoVO8O7zwjhufAb8yh1jVjenMRmoGt4reapu/BfUlw0cmLLaz+fgCM6KRw2kg
MMwYyv6gTQJhrK6QlzE8oFyPQxO9kKSbpVTOoWSI8hvDtaDyQlGEBeucT32DKhXUK/gBwTdg5Vvu
zEm8aSQ0YH5r7kTBaDaIry1cleThavaEXptw7zUo6x2/7wswgW6xm/TYVTRSyXd7BZJVKDeATGDl
J/NWrCR8uRReLh8xTsGxuzT+dqifjiD0dmHlfjxGKsmffZK9rtLH3cUYYpeRcfjsRwOoGqkUo0Nz
rwAM/xhcYm9c7x+f/xKItIDOWpwHc7TNLIMmWkifhlwTMUg5vrwgdVu5b1mAdiVkOc0bwbKrIMgI
lOoK4wRJ7n3sWeT4iHZioPQktXfnrlLiWDHPT+WoV0C0LEm3+mxrhqGZcfjVe8QT+EM+WMDULxoX
OsFjGipM9UGtiQUL3NS/TFa0fQD8lSoXvzA9KdWnl425UlzoQvTiQlPxfETlMtdnmb8VlKh7QDfX
Nei7t1gT0ITcIlV3A0yIW9+ltyFiZNa8AyAhNBgG0ZqlIkIescQdSS+nk6P5EQCZ320EGuboqW2w
1OD6UOY3o8GiqFWkApW8evTJBlYV5y++byq5KKpBgVH08cYRz4nvj4a107DHbg13UkAZud+bkMi1
ESHRNKlivKOFHGnUui/LoFPs93vMC7fJ37aNEP4vqzqqf1GSFY2ofG8mAYogJ+lZYcJ/yCK8mH9l
OBPDJ+wFZks8HKkr62/z+M2L+pw3KavBKoW+bf1Gxo3MrizpQCBw4YipmK96A0c/43D4ANRw1heT
lXtWGUez0Et/MqG1iQdwC3xsEzykfxne+PckGU7XeBynqJt4R3Ydoyo/1DzJkmwCVL4F+S7Qhvcm
vKngPPRHYg0hwZLjasDDrNcY9gTvW2N6wJRU3ajUw7vIwdKUTVAlh2O68BARK0ZpSHSMrmKBL4wg
y5m5Crd9dC91cQ4HHmsBS98flOuQAR+vEkLZ61Q9lUdyblux5dw1WzVRq68tmqtQ9m58NfCxFHQJ
awVpaaaAhb+1t/Q2OvJBfskQDg9MiZ9n6Bc2lsjsURJXOXexjkpDQdJ5Jkw/cLhxWkJT0KcdNCKR
5TbBEiWSrSmobvXUeiBqeGPYwPZKgc4xZbMGuwt9r4mZrObkH1cHIt16cy0xRO6hN8EzqW5WOYJe
YTn13lPTnOItC1FbsaEaANre34CmLxAWQyaVU7BtBLJMq19bc5GT0MQ/Dou4MZdJgnS1MlXsgaKI
sClxlHLgQ0YCYc4+/wrUCx29BcPqqP6zjx4JVSpTqnqgHJ/Z8vl5Wk1qCrVBqp1UnitFieVcr3rJ
Y1z7kTLCBA+bnisRkIOh1klYv1wWPoEYi2pVi0RwobTYOkXDMIQqiq1okCeA7OWtlqALBG7OlGkF
8dGf5qTYCS83fnlJ4CjdFtZRVoYPujv1TkHud64htBdlZGznW/45Qb08TgXPWWcri+M2Xu8cQYyb
eRRQoIHV11AQvCpdmH/ovkdWdD8HA62gLx1UywFq+dgDwe9wbq0NNssBqzjjfZheLLntkROtn7PM
ImUZHpkhRhGQL2AG6ba8nKxd+e2y9r1Hf5heNnHdHBY2xMeRZ/V2m9URhJHRiSpy5BHd3GwrxMSn
XXChyR+g02b0JLDNFyufo3omKQD1c4OGuxGVIbJ89J0Lqr/zGOc2b8uyEodpb0Sds9biqPrL7FL8
NlREPGEjRC4VZL7QJlVPzKYRZ24dxJ+OWvbVu2WN58B0w3LJKCg4nOfNqBDEt1zYs3Tqg/UH2vw9
pcI8FBcxhsyHDELhBgOgMaBONh+idKVJ69rBs9G2M6/Zq46xAdrP5X2mVt27Kqi2epqfZ9/P23dB
/RS1bHYUXL8tzTs+fV761fg9Qy3fiI1eseiif6Nng0aj232C4amoThwUaVcdg5lJQLXyhtq8qt31
JHmpMMhzH+mlxM2OopbUwaN4xep9nxACwMvmjV0XgcL0F9BA75B59+fO+yXGkpKYe7NXniG4uS7o
FVkPMvrlZrWXdkcKQ7ozoT5oGKcrfNxCmkShz6PgqzgjCDcs6jbFWO7XSoYN5txfYSgR8ykqGlnk
WjKGyt0D0NwqwVenHr2pxJSm5/VrtsA1gTJztBHR/S/k2jL4rXJ4EXWYlAHJCWN+B1X01WxUFHMW
2tTNVu6Cl2Ujmkk1VGyLFJ+wNu1X3YWty7vX3VXn8/MsR6EoyturhrE4YMG4dCZ+rdNLNZhfC9gI
pkHcJsHwy53xEqDuM+esbK8y0hZ7xdZrWHQAM7EkkpE6W/zpm4BVvvy4NAeOUSizIsRstvZeOzMq
3QqlX10O/hq68H4eH5jekHmPIAaIuaS4Hm2aEzwuI6c026UE3KacAyP31bZIQ+Rhy1DUr+kdwF06
VTpZEO74/EZUv4URWV7grMLD4CFSjqaOgWLcKNv69fYX7bTGKc4vKcsgxEwUUgpOSHB0wUo2MHLL
nKKrrMCqeVPQuF4/3+fz+71ikELiIWPz4TFz1fsXGaYvV+5dtrAmBdbZSrmY80GiJ/cw6hNIHyw9
9GlOL4+OTwtYqRWa1GgwncD598L5a1fNk0GO4UZKyU8RiPNu5M+3r0NyU9aD2ummIUOxRVG2NuDh
uaH75jf74V2bVvy/sSqLfVtXAAEk54Y2TP7b2Si6M1bInXJfAR9Deybu8S/GDeyIamuVpujMNrGm
mxN/YWpWC2UTeUtu7uZ7IrMWt5tM/2p/ZuZIOlE5kRhQFjc5G/j91xktK6RMXMbMDddTj5HcFGeI
jqxqMrfBZgvWr/H4TrWGyJdeo+pI0Aqt987O54rvzF02UmIq39hDEd49kiDEiemIK4ULPZcrkHev
G6uqh5XWbSnHTjXMBAVJdfBSO3JGfCthfduQwPeRJDfl5nOerwjbizyxqAGitH2+nZYaoA3rfy2U
RHhCGJ17ny7WJABc7lmNg1VqdGEb3CRvf2Qr07U+FwsWNfzmJpaYw1S/FNtB4NOgR3NxhKNy7rp5
5aKHJILxYIfHQ8NBAh2Hr1+2Y2JVdlldD93uNby0m8iclxqnGDK+E9bcAqgMAa4Zo1xNnPduZcJ3
L7c7kMJJ8gkmv6+A7phRzXLMS/S3IRCsxyiieQaggh6S9MUCFKVcgu4+9ONQP04BheDAZpbrZbmJ
CzssL07BfGTMQWoVmce4cXHQOpAvTDlgjb04lgpqZN6PMhzA0xH4Fth+Qz4NgTBq4lCxsHz/cJNM
wWU6f/E/1UKLX4UCGT6fpy6i2+02df/ILRhKRtl7RCc+BgzzuVp/Io6VHQuUN5yaYjErXooZBP45
Z5f0jYM2DUdgmsGzr+GTnsCrdyEEiEClyTwKP3wYP3xIUzi2vWM6+onqCP4oaFs0XbY3KhTk24lo
ENd+LNA314KEzz688MjeFv338khDEbN/UcOQDsZkYh7BhRYSfHamTSMw3v4bJpShwjcSLsH4qJUV
c51E/LholFJRHuFKeA3ASSk8tFcEAqOyc0VRp1mcD7qo1EoDMQyS1XBC97GtGvl0LWLd+xFXGnzE
HmzfTHaakY2ewREXwkMJaLM61psuUARM36CSkfGKsvAnhTBsk6mge+FswkY2DPGAQD13MDCpUlgs
fOqskmbRCHW9NNnl/vM6k5FHiJB9o6nQmvDxd77OgqG6wXH080+o+a5djElGYsKHWu8K0ZV9j2K5
kMyBateyE0LGEOopA/k0tTWzQlMkDldBxTm4CRgfYzV1zcd9+fUL4c2/2ZN6h4uaJ4hAhiaRQVIJ
Xe+b0VwkwPVZ1YOdQ+AQaNIvX72WZLCk+KEfiI6x9mNic2ItpFx+l4wTjNoKyaCjGzF16B3yHW0P
Y0cuPejprJeGbt9eNQZ/p24kIJK+ap8A+3aSd/3ZwlLwxS0DH2wlrHzi8gG9XlVgCpT5MYVhkBb/
vz4Lwwjn2sSeOK7C09WJCwiJ1iXmm999mtay0i1PX771coBH0AhHjOwQyOpIwSt6J77DOFdsepq/
gOxrnPSWuqyjCg67TlU20MHYH6SLXiXyKUxs7EMD8732rKCanuYflaWy4Dk4Ec5Zgb0Ivx2w3lie
bc13g66XYRD56iplTZEiO69+GnqwarOvKfVD2XbNwIpU8uSQQ3P0Tlyq7kgQCqXYvc0bB28AC0dP
Co44QO2Y91AYi/Gu/a1rfNAc+T1Z+MxdhnqkV+/T/nqC/oiikIoZQruXD1j7m56WY8cuV2jQ4vyu
FQ5CDcjL7GoVi864sXwpftO7fk9ek9BcqHeKI0Mv80TTTzRYfFlhNz62kN6lqbAojoxE3ss+sTa/
cOvxsFh97mQEganhvoOiVMbrUlEqqfLp667b+JRUJ0IQxcZRm+ud3mS0FkT4HQf0QzkzM+Tb/26Y
4i5e3zcpW5VqBU2hOD5NdKY+x6aUi96151Gyppx9hbmPGYNG5eYItsMLqxdlFG5p72H+Pot7oTIQ
bcd5lRDajPkiBCQT5A+kE+8GIKM4VaUV4CU4zss1rzHuG2gzEqh+traWnBjvZbrnbEaNnjNFmNsf
8M9MxL7UvV7k+fP7k+K2QBAV13dvPeykZM7NeimVQU2F2mSnBDDsDUQvj5Px5sATGUOyH4Li90QY
7AVYWeT6HIVCyFx7oGbmKbG5GIyW5DtIkFPvd8GBg1VNXz1n9cy5FNAUy+bcLOYQJTP/pPWfQaWK
bn45wQ8jos9Y/s/C3yalILzMGPNmDN1gPfSzMkg8xs//JZm5y7lAmWs6tPTSYItVDiVDSSWX9A95
Fi42IbeuaXyz6K0CKfCFA43pFm91U3WQswb9G+G8aDw7GWkRrbUU6lLQLMnS1lyl/pYLFeEdKMpI
fa84VDC008+675iEw4bJDH6+aJJtkQXk1WJvO3vliPtwm0c33i3rfOsHYZIfnU3JjlMGydShCSyV
oqdDFpj75M99DL25g/qmdFDxHgFupJXBYbK8GpPWA3525t/ZuLJQ8jw92TjQWQUg9VHJpQAGYk6t
AZaanM48hxyWGDqqFyD0RyG72dzFBju6aw3E26RmpyWN4Gv27Xk7EIyF5PB3s5+hWk6ijHE/5Xq0
68qcRX6cDBBHD1YED2OaWL27Thjc8UnsGYCu3fxmdtSyRFcGX7LhLdGzy6l9MLcLagV87Lu1eLFz
DmRM4ClANZQaM9J/1OQiweosQAYdzsG2MRFuzqUGTYgMgJdeiNMuMLDfHkGMbqve7xymElMwN39F
2cYwR3B1bqZsnl5tH9pDAYKE7bwtoApUlLeqYNapED/raj7ZzW0Nwkn27yfF1BkKcARinHOkjEa4
B/VikA1Mv7cj5QF5+wpyM4qwmTKUzuyIoJxoTSvuZ6SIr90rgjCCJRET9c1+VsGgiCYKoSPnz1+l
/VHrZgBx2lycVtI1wAYHGbDMHw50CVflR2QoEei5CPA95bE2JjQs8VRgF6/EtWaeozyPqk9XxAlk
VWQf+3tGR5e6M7A9Ft67ZiK/+hmtgMmfkLaWXX0VRYeQGsI1ZarIogf0e0ITEBkBtq6U4PwVQncc
srarCCD2RKrMa4QcMHIMIOA4HbjFizgwJB78Pv2Cy8zbxdocQVkRtVAwQ11fNRIOmVKF0csk36tx
AH1h4BauOTt68F5LeVonGuTAQtFQCN4EGle+0JuMIKZV5fi3vN+VTxIHggYUqr1VGbfdqWzQUX8p
LQY4o8Du3m0Cx6121ijcrdm4LNh8y3WmaIdmh1/2cOBi97iz8q1yRkAba2itlOKizsfAZY8+4uW7
V5USdjcU+SA/s8Bdk6wTXqFsb75fNrlfmQYowI1tdPwtitmB4K9cvfsqSZQYEGFq8DtVMCE7wnq9
RR75LIBZJXN+ENRobLDlpbFAlp7fQVVvJdWyYKUi4Jl4kFiW0MiXetxLRECX1qVvkfzYII8tSxF/
Dd3Ro6A74pg1cAyS1RSongWun3GVEwPTJy3TcUCdAL9hzfAkhHymbmRMh1f0LHBs/0J6Rc5gK1+I
NDlGPhPdazaqH1GX+VRwQpme6zQqaAQZSVNDnLd8AhBbssxZdl/DSZ0886BDwn4Tg8nTfxUuj4Iz
FelgBSorGkWUvSvsYxgNBHq940qEaXAwVSzI3guA1n0p2Ml8U9elwMjgSazS3jDbzhGtcykcpSWA
S0BPqNG29zritDVNzZgZ9wWYzFkkk5J+LLZiIFYgGjAQkobV01tdy88frGpf4LbBghT0SOU8Fcea
GYM4QM5mdGaIVbExZ1unF8oQImu1fuW5lsJZZxvx2Y+laBU+U/4KC4ouaRCScF69mh47JuXhYCiV
/FUmM4LfEqP5mu9RZ0+MqYfC9kAmCLUDBvj6VMKQAIH5JpMLD8Rucc6ZcwuCo8JHT57C1RlyV3XD
3L+qjfU7eB7spe4Hht8Ngv5LGD2e0Z1k4TY1c0YU4HDFwzxOE/a41/3/t1aGBIOn3v1n8Q6nUKtY
WH7epE8qcSoSto0VQlKK+uXh4ajObHdZDuLcYN3fhsl+YQ6kCNhzkLLMDO793V3via4Od4LdMCxc
64uPJxQa4DKEwLDwQjbIe/tJg5AIWrKvmohx0siUNjrzCENdSemaWL+YvPRj01pSO0lTyfwV9qfI
Or92it8A3rK4SOXa2R2M9entabz9E+CXddr1SjszjnTSN2HG8iX3aWr43XTml/EQLfJtByQmWqsi
pOhLcJqrKww0nXC/NDfAq1YX2E+aOb+AKNLWNq8NcISFLc0iHYqjSPXgXyuA4EmjrfPa9XVj7UJK
komaa/lD4hJXtRsWmhfvOb5zf/rhwPJ79H+dd3EvEIJPUaB8uJ05IViQBMIkCrzlOPs1KxMRuCHB
Cbda2uOehIDXbf+RjlPtK2jk66uqIUTMQ4r6dofey+ActU4XkQFPNMPw0z+rYnV5Q4k/ZO9EuAcG
pm4YZjTwx68r4LfX8B/yiAQhRot4rRw/lQNXC+XIGFJ5E5pA6ncHeau0upFS235uwCjiCWtnHBBd
uxKfviuE0TZNebuUqeJySkNn+04NM0Q8imUg1rYuE+GfmBbMlp4xBuWel08z+zRpjiIJFG+1hUm+
k8zL8w+R4nZt4eQew8P8cE7ZN2DhrcvUg+jsV24RchgTmHiPkx0661BNoVuSdAKYDEVJ1natuZGm
mKHYE8xV7ioRm+0c2mDBRn1UCzv9dYERkgFxUvXErB9IdIKHYZqXy1yoxcHBwYdsc7VYsvtDm4db
ILq4whdpE/ZbMnhm54TjLqYGv5RedKgSjAu4/A90+33N+61VnS1LhjZ+E90ViRlXXCvmDRP/bOiq
L0UgjGdzlbHHUiRSDP57ItnBeXYzdTIwhn7TfRn6FGlOp7AynitdkNnUMRLWjRycrDMP/MDXvHJR
dDzSsOL6uqKhVxji7RdlKxkdPl0CZ642R5A9vHjn7XYp1QfpbjSnNpCSeJkRE0itp/ERG2oWhuPz
yFSe7UvPkn7chOCX346S0V/XoFjHwOqq4zBKRF9kCg+9nRjYUuzC5kBhrdT/eHS8sDObZJiKJifC
cTHGqUINrsJcif9/b2OS2pIGuK4Uxxno3ecWt9pgAdUIq3grnBP1tDP6nvSOHLOWAELfScX/QOGd
9Nkqsgi2clpxH6JxrPJGVlR5lzhWpLzqEcjgP7+auxr0ZYMLm3HcOuIBebDsgm7KJ8IzSo3eHmvZ
8zVSAD1/vnowUcj8gV51awk3Eu/oOIjc2FKZEGpEBqRVpxC2OuqvBvMjD7s4Lu6c8Xf44ksm5Ei2
Opwnefb3fW4txq3gkkMjojzvHHQBl+ugHduX7TAxpLvFulZZ2GUFA8zYM9iQBURaR63NQ9tsyo/v
8zvdhSpuxo0Hd4gUIp4gZsBLUXunor8Gh+rfjVBQ5N38Wzl93+ruljM0t2Mab7bGeKfNLGkO292A
4Q8G+Oeryb9lQLTpo48tuw5qeV9fCQL3XYQ54PlDoLXPeAlDdQCulMEV/wBDNJ7nD9mEe823uv1n
vW3boQWq6x7PJW/2EQy5VIta/pxfWuNFKy0fxtO3W+u60LbMJwWvhZ93qncNaswY0rS6UmboZ71I
3bSaM3cDH2QUGcrhDtgXIkFS0mZvm5nzzMN2BMM6COET1iJcUsmM+tKOz9xPc3kUp+6DuJQnN4CK
6XVcPZ58EbHspLWCCj1ELqs8zFxWSGT4J4202wRiQDnWx8+bGbQk34/CDgrFpsJrJUVhl+VGiCO7
tLsQEPsWJ8ShWow0lR9prj8cI7r86YXl7L3MjH0L8Ju5QeYBxI0ESm6FZYJBqEN491WYnTsyiVxf
TAoSiZ1EZBkNu2r002GBTNX1Dc87tOQV5jKmWv3S5UVkn/SfbASRPinhrozJIcLEGq655K52XQaa
XzYtT0cS7U6JDvXPJVUwfhYoclBdoxTjlRK5BtNmQqIc5wVTDmRrKj++g5bxYljQGlOlcv/dVEsD
BWD0L9XqPxzohFbsEsK062FQOQaWho+gorXLPYkyV8y2+lxBAJwNFGF5AHN7aufHl7eLMIkJfkKG
NlASP/rabP6BKZGXxvFkm7xaz0TkswgbRiOt9hOdXS7mP0Xq9pDYMKRrPiyox0V/UsQvTUgXhEYv
cGYcZIfCtnXBF021BDO8fIuCj//0rgvSFX9mSb1TPJIDkq22/i0Br/WDs6qibnZfQBlKu0jI2qSx
nKGyCRk4eAvLCT0za+CkXTtPZJ0zA9TAh1ayko/3OABnVq7MwtIYRsnQq+RYh/qsZTwhovICkFS8
sLyU8VbGXcSeBUuNqnFqPMoFBpU0rgzuRm1GVTI65saf9cFfpDcTqqfKpRRXkTGoPKbKsZ9wvlkU
+OOtffIV46YrkezMqIydVFfFLJXqC5voUAU1+jAbXDmT/lh0t/Pch5FIkr/H8mP5OfQnWYd0Roab
QluVAJ+fhWu4QMyx4ONpJk2R9df1z4eHefsP328pyH3M5Vl/iRJIgHQv+bT4eYefh5n5wZaGO5nw
DILbpuqv5IB5qwnXM5xp93usphsEN33m6iUc4BQ0aHEaB4UAj7A+Kq69xn5d3iDDPrsQaZnPsO+m
Lu7BfDaI4tbjVrLFpBIXa/M5gzGUHnSxqsAaBZ2zd2FwQUQ4fDidYCAP+a47o8cEb3iKLS9UnL7c
kZZ34/JQh86As7MaD09GJBQFgZVIXedW89zXQeJrwLFFt+Um58mij8S5pjO4+qLWzhJOWjUFAcw9
Wa4Ff03pWmgxFo6zR39Pwq8fYGTraop0X5phUuROg2hPuc6mgw4waGu0WL+w58Ipu6LtF3j9pihe
GJ2t6RE+SCtXqa5lVnLzqPSYQCIRYMmeIWh2cY/+k98CzwIK84vfHMOvWdFMSyB8USWtnaRLj0xt
049NjCM+SYWupyB9m2MOqwA3Zt9oIsM/zix3XXX+e/DmEttTZrAtevHbcAbmcpe0bJ07YuKA5pDR
ny1AE0yv65RH1vd5RTiY1eg28FAilyfk2CXBtxCTD6FCH8R05l1790dZ5VuK7iGf1hByKgly64Ar
KSLhMOgUFh2nBtCp1cgVuw/1HW5cYDix1pi6vFQCgFVXNNQYsVPKDsGYqMA8eLlDFkEO25Rxummv
eBlocSdFphToF7GsOPzZG7uoMFKaC5rg2+lxsmJgJx8XwlgtQvwp/+Te+eODWxaszGy3y4j8bfe7
hxYca9ca5+Z5qobDPRBEGuz9sjQyZbbdWwK2SgfKR0PEE2itvVBbi/idJPAMNhxKdsb0uQknGgIi
uiIAf2r81+zz9sAsvOcA0DW6gq3gMoapgtcjrKfRxIGPQeKUq8GthSx7AYwP2KTr3+Yq/mi8pfX/
SwwNy4Jpaw4+0DK5/uYicOiloRpcZLVxZHF+Upmlu+dP76oXdBWW/ip9cESVt8bjnpMJXngz1YVg
uDCEj5PQq/73aCHqIo0f5b1bEYqHPR6lbZQFdjKDvxOBNux3m+6cjnK4yk5jIRIjgn8LWuXf4IT6
DOphla//AXKdVFClrNpgtBch0kLTFOQr59j3eH809PSHriiBBR5015Nw1im9Phd7RWtcSCQGD31T
MDX0ta/qhafYswE7Qy+60zXw6zcKhNoUVaMwDENhN2Mc+sTX0HQSa2my+YJn/VPj9PDW8rH9s+pJ
4gS0Wcv+ChH0IPbmDWf5GZwSEOYqEObJkv6E3moKOXkF8a3HYTnDV7cYrxxVF7hhszfa/pTASo/H
2o+eLrD25XSPefQ3yM6Too+lgV0afBFBMJ36Ken/xRu1dFiRpKXA83BXGOidY0ef+8OLoLfOFce4
bPOy4QOyfk64HSfnD9aXixdDbSirvINZ6TZaQPyT7rKmRSWolRGTF5VYo8hzdJnNDJ0iPpn+vfd0
OgNoxe5QzsnaCN9M+Ms0FrwgsGM9i/WriOe/YKCXKPFS6pwFvzDCcJaENxFYlu3iUmZNB/W8ksaT
Yxu7y6ota1/chpiofiZhKKoT3WCzvLNlwWjsiaKYRX9dOFmGI0gl0ZIOk3Kfs2OaYqouCjyMeI7R
9I8lBXCTFL0Ddwm08mGTUloSNIwSSUyhIfcBkGXucGTyoYGPXXwwQ1MgWDaNJeOyHxLKQE+q+Wmp
GBByae1DMQbCKnQn9SnULSK4VKg5oS8b/Rkg/hTL+ziiNAyo3sQ8iqUlLeoYMyp459bOoheuhFq/
GtAc74P8IzN3tOuRb04DWdpmmFghi09JUsMEv4whX4bleUIml+K5XVyRwyjb+Az+6Kj9FL0iqQ0z
zqogvwV2UhGIB1+HBPbWM+Tijr+oSh4tBlPsERBP4VfVb+lfM5ZQH/r9jyMRcSb2cWnive1IYg0R
Cdk87VHSspG36U0MFYh0Iab87DAorXXyBE8SF5vxU+kSU26/zffKCoSF+cYkPk//gnGoTFclNNBy
R+AvPjOGRNHIUOzEfgjZd4VX/KY7RT1iMcmvzA63SR8waEIRSSZhneB4+ojV0UAKNlpQaCFUoI9e
SHK5UzY5vFO/cKsiUusHXIfu7bfjf+zFaUGdL9dDtYsx26qJeh1YwwiBP1OJ2Xjevz7EcKfymdxi
ZvnKHHnXzNvluS4LjRszOVnFi0+jXwvpUgMarxqeqSho80SfM5EYa3uudVxr1agvFGCD6WhWNdAM
UQ+U9rQpmUnlwWWTXxau7qirerBTR6bGKPiOwHT5PEVIWVWRINUoR+w2s3YPZ2Et1ECmvl5gsB76
FA5+qvMYgLSSwuh8cVhc25Fc1E+vwRm3XHdc9H4yKerepGbjtjcx7xELLD+h4G/lpKFeBOpr3MPy
N4CBcDeVofWJMrp26WLRZgDtgeHTupAEezRyIe+XTkIP6YjHSr+tzJINwOajhqNvOKJvyUQBIvkD
Mx7E4ShqaPw4y/ik5vbQd6oDwK/2RHC6JJfzbc2STRkGvCm3u05J2oCuUyuaVBvUiwqQJlfMgfxU
4Gxzn1WFTzrGB3RoR0ehNB44OM0KBKZbTTmNROmi3QX3ObGOTiwxqQpb5mg9VjWOrXWlW6aQFy9L
d64B1qwJfGm1mFmOIw5vX23Vqrshh7Wrmv4k1GITc9eNMCLgSTXouzDRpwCQ2ZPZ3T26gFwwUy2q
0/GK/43aFoeO64qJbugGJDvz33YVFb+SS89ireWXvOy8icueR77I+m9wLMOqrKIPQ98iwZPZ0i/1
YW5sEWHRcrW4IiWgjG4+vbx6SL7UrfXlADJk6aUEu63cg2rSoNR77wjRYAXntWeYQx5Ht/zMKQZg
1eNAVsOXGnWr23vLzgdtPbp1BeN9EH4ZvwKWxiq4Vzowksm/pB2z4ZC0xX0kjP7pmJjDS0C2UL1o
SqUvEQLb9FkXmo105uJHixe/zrf2FhlZXGKhkBz5R+4Ndnqq+RcmFXGPYIeuU0pD2hsdLvTYGsTt
3K5hSHIvcMclm3R63eWnejIa9VKsc/XSk3zbU3eZ8E8R+qnnOFbCnmZTPkWX9ktD5D3gNhXa9xMf
9Xw0Oi6gG0LYFQJbatSzOuC5EuU7uqrYk1KAoBTuBFYyrsYKocxsTnNuE6LGWzTopFrABjsllTNn
OP+tnDgWskf6HTtAJhHzguAQjZnMEtB7AJl4XZMTTmHUoY1W7kVf8G33utoqj5JgDkyu0Pfm4NWd
oAabNiTqa5nvdDTKVEDQE+R9SxS2GqoF8p2Ey2e2OEq7qJKnznm/4iRBYi4T99aJAxISwAsnba8z
lgSOJhZJvggndPh0TXmUaqwm4oxMQMQ2L1xDaKRuLrB8iFNkLLseBXvMpxXzGw6G1fUJsZL4xn4P
Wdz9ngzNModo1FJaVtT0ubQ1178GljG3zhWmR2LQrKi/KyBZXVI/XBqiWCoyJjvl44ddYimCvI04
Cd0youU1Pyu+BQl4oecObzVlXjXrWvNK65J8LW5VTwAruAfpkEkfflXTMgD2bMnHDesrVVyUqtdC
c9LZb72sCV3+0gIVQipj5xge7BYYc9ROmVhZEQx3bl3XogqXgqMWY1rqonQd9JzoJ1gZhkf48aW7
ABlBlH/+oOhcOb0rFFy8XkDgsw5QyCS/vZYWiwLzZjMGX0z5nPUPTXRZovw3HDUvWM+aHquYaBcs
B70JLtqd1R+rxAPdhryvwsFdhhWjT9q36dkX4V9knWTZ4MLPhsnb8zLu92SbyYTbE3k755DQ8pom
SSFAoJTL+9l8EPGmi8pAmiltBe8xtHCQSfMzfUUusAm+r2P6/865SpLMic9C/q08AbC5B2KPCPEE
iGBZnhR8Ggb+40ry+BoAi3tp6M40o4261bTfrCYsaBt24zPD63/oESBK2IZ1lkwDbMd2hGOXx6IO
Qt4FTIOc5EEejDLu2AqICf7CeET+saX43t+HF6HZoAhC6P32Os+Lj3OID/9my6HxqFcMDdSk2vyL
lc1Ogtl6cZqNVTq8bpUegwc/Flm2xZF4cf9/57gTMPvAidH8l5Np62SSmaEToxXe4FPyT8yrEWQk
SBA+XI/pe+lMryqoYw+2oezS2PD+fUCtzie7Uf+dGKpQeHuGTsWn2vKnbP6cDjn8ZRVeAp6FT7ox
dbngCMIhrNauJSGdTMgURzk+dygwykL+jHJ/53itDQCLQSK03NPsc/2NIZ7fDM4IN5OwK4ha8U1u
/XgtAP4wyJiUOZIgyn8Q49jGGhiJsaUdz5jF9RtWWdPlwVY7b59wJWTMtcMS/hieyLCoIk+QPk4d
g9kMH5+j76jGzo1kxIr0LxYIbftpf+L1UBzgUqjiVXxnCVMiIdageU1UUYRcPhK+yjJMUhNMUniH
J5yNoYMVoG2CLS9klTrvKUM/EqyiB1DPNZShlYTarODP8+mKba2ukKRmGt+04/DkngOMwmBGzxKA
W/Bm0Zzoz/oZPPdsTgGl0vVyZKfxbUVAs7NXppYOMKECUhyrWkD6Zd+jiqxVqI0a4PbO6cAnYaoj
h2mGYHkKcdHLmHo1H/yYfSyoquznYVW86AvKUGErNJ310oqeJDGv+/62EtVTccpv4Ra1mtzqg+qA
46sF5Ds1ljw+HD7Ss/0oxZnRIZoLDo12jjTjcY8ZTsK5bZFDmkjObBBMyuNpx7jdA43rJ+WSBX4A
/iT9E/N85pmJptkD8Ni5pqLQiudd+4dfFnL+VdyiyEp4qDBvCSRq7RQkw9F1+t9aonob6lyW+wE0
ld9qKtd6Hn7WGV9azE2DxDwJBI5eKIjfV74z0xeespMiqPNyBp0J1UVAR9A0yn5i+CG8/PHaU9S2
WxxbRHltBr3PRPrDmhKLGk2CSJhFIGvrBDkSuwMWj0YALZZpdD4sYunve55PcCCPBcKtOFaANFoE
lTYvHO1/3C7zXMaCho2cu8QJ36b4PxFex5pXAcRCm+lcyCYnYpRRZUdVP0i6HZYLbQf0I5wAMyUa
J9qgtF70Cn+tUsW8pq08DwZGoc3F2xDQHmYFN+wrEOOzcoVeM9e0wVbycsdHfaxSj/i5YGjrMfiY
sKFqy/cLwvT88oOy9u1ZDtyZOOqc6nT1KyTuWjkDboolq2MVJs0NtIEdya2SOTqoe5lhXJYTd/6z
IfM61Ij4AcqQY9R4GFp9ZTVYgSa298GvEa/L1BFesYM/cnrejI3ju04fk+qA/ifPyWoWl4rJTOim
SOeMME0EvpVpDuYIlZMOvFmyTG/nuNMPf7GnqL1YIUUyHBPCT9KbwUgI+n6/UDEykLaeXPtbGIkm
4A985XX5S0nmoed3p+liF8zoavBSPgMyxmrDaBmQGtrfuncET5nq37vFSLBYcLLYpVL225uhdN1i
v3N5YFDjrPtl4dgPBfBU8y8Bl0EKCpRtKcv1TM+nFdYzEPRiSs0iIz5+U5dn62se16QTn3UcsZ7V
wPHzIx44Bx0H9TDan6W0nvTCwAD9cdMZCVMwEXlv1PV4jxd4Md6xNBLATbsRR97kV5ibRTJ1nGWp
e8vMBlKu3+YXiugOH87XAyRRmFfQX9MOmd5RRkmMdsoWiDIPRC37QnO7Yjl6duYj4Q5cwV1k0htf
T5EPyIUsC5S8o5OW25Lmmt8/KQ2ruOovVZqjtyURjZwVupTJKDYD87vKpBxVppR/Q/HxFqDj1gLd
CFp1OT22fdVZ3bn72yuKu0qkzZWr/cHuHXs6CEMchfi6HKT/0gDzE6Og0xpF5vGamWwWNqlpVaVF
XfK/0seDPrq9oPOZRT0yswQwGdgVUWl9Ho3fXaNYCre1vP5BBvv3zky2iN57TSUCGdns07Tpw74X
5+EINNJrI60GvDXGZeHj02Io3stKluh2cD3icIJDd0T5gsqgdX7g4JcK7ePq55/1O+aKNft0cHkZ
QGV6A0w+NOyLMiXRldboRhg31LBeX83zHMGtR19kFp7k+ZGIim1R6zscWDvX5QxtiwaImI5+eHd0
N/gVk8VlhhqCPyIAqM2T/tcN/x1LyLy2fJkxCDkR8cIBTzTKo+3RHg6Okz/XZPABxcQHbTRG8IeN
HyGhCGVSNleIFGUUANdsmsdaDW1TtQ5SeWuZkqK1afan2BDox2TJJ0ObTgqI85mTWbEGX4ugHGvB
Esw1W08FCjfvPCn2ApgECzSXSGgbOyyjYbrddzhTD2JHXq3gyYCYolFyKQPcjdVfFAl+B4aTkOU0
v1+k574jNt9+XO5zEei6wjpTdwBkc0LqRiruUnWWJXeFuHWcGxKQZfUXUbhNCTl6VHvygluhELZf
bRj+W63RmmG8GH+sYOvX4yXNpvzRsz+Xt7xl1ZT/Y2V28obW969sX0+Se11Oec0BGtk2Rp7IXOx3
Z1yg3vxcfCOUp8bcVwnCYj+2lWnHuNRmzibqxupIb6UlLV2xD7BFVI/hiLMUx9RwhtUN0iWeTdy8
7xSk6RCQc5NGtLH5v67ArxJuDZnfap9B5kj7V3J7V/6xc95myFEBjQ9LXVBvNamPXjdu3NRk4vt9
KswsgHXOMN6xQo9nSRJt9SlwSZS/KVA93bvT/xj0B56yLY7LFDeQLCnymcDtSLrnHB2sWSp9uAxd
8iShe8kV1iYUvWSd1Sr6PFXKBVt+BKFxpzmrlbYaSwDF/sB7MtahkX4HX2XVyqJwKiWK9kzgLhpm
0nnnxhMCSyy8pptMleHblLRuLIfmeOmy8ijdFN5yS+08El3tJCmWdjP8CrThjsBkANMNdwENXSCp
IuMcq/PedJXkw/27hlBJvjxwfV/6EW53hOCDU7FxPFnfaOZ9zCiMfCZm9SZY7p0rMDgO0C51gVbn
v4HGD6tBPSCiabZxpx7LhshRXgjnpb53qXUU1dFGbF73LeV0xtLs8VvAVOkxHD8WZ7WfWPt27M61
YLZ7648IEe1dxiRArWyw4Emsy7W87gX5asTYhJ/UNnAXJBUsSjdYuqSsZWp+MOmQbJoDa7lpbAxm
BbL7oiBR1pl26zZdZAJuwx90aJ5qhK4MZe76Mxp1j0McZc5NT8q4kPXXLPOJOy3XIl+3CfoEiuug
1InFiu7O6QEaEtdAVJPHjcrlQzWVlqSYCWz8GyFdDSpAqsUiGnL2CIhQdnlGmD3SBD3qAyAnUuPT
RaIqTx+K3/rWlWO6nvZ0sM20eN05mEdkOsorCUl4Ic7fQ+XdqJDCNK8Rlpt/N9ZRcEDe3+cFcwdv
5V1MQouNtAJqWUs7YsQ6ZmdZ6jt007mbS1WTfCPylTyPRJiGcO6FLTqwlzziES8lE3od1/lV3ywD
soQKcCBdeOPGm6Nbw1q+pipkx6bFTUeA6oZHdLcJLmArHdl3Q1yRVNvW8In1EcPeP/bzWdZkYeFn
Xd9DsBdXzGCDlSWVHkZ+cheidBcsba+ZWXXn90HH8W7AqCmeCkbYBB8srjSSrZVtdlxIjehZHAWC
2Ax7UprfFVe6K2Z0p4ky+wn0Tc0YZvHCLgsLDIvHXYZmVw94JCOvcNy4WwxsubmbPMa9RaqH2bVf
1o67PfdFVfPqGKGVsxJ51RALSG9ITMoej2H1BKngojCLvsTfb2YE85rvuhczn/B1zGo/hSTj+mAa
n9BWHl/shuRHw8oSHUw0C+PDnqKrr5YZX4bd7U/yIVDp0l7U+aHFE/TsKwn/4B+TjIZ1tOcZ/YwN
p9nBiH5zVx8lQ0JkZ0idzulTVDZ816ckdRUOs0yk3k2lApF3uzVxMeXownrgUil88r+of0i3qDcJ
sC6gwyQWIwiT3o+zent7kYZU80o8d93TPSHf6CYzem7H/JoZU6Zn44+BdkVQ/hweeH1eFgWCC0QQ
3U572K+W7e7FzQCwq2udsI+x2/vB3+7WYeKKuhXea5NaC5zQ5QHRzOCohGjfhmbRBwzbSzfxHgMO
8iTk6sLRykKwhODGbUE52GvLB0XEE1NIXNi2ajf2aCCkpmNq5L/dvlq//v9Cfq2mD2/Z7WfYf5A2
dT+s+1a/yuXf3m2QxTpN7MoGn5W9EP9J98frbR7k1pQJDbYUuI2RmObWj8Vli0mXF9+yUJRtpTNV
9NxkSPAsyCdRo9a2t/VBPLYRt160LcfDeB258D3b1AGHXwRqxabJuAn1llgO+z3UszVwHbgbnX66
ysH2uKD3nZDy1dwIY7tjT3DobCfq+XwVBVggY2AHImMNs/OTxhGKqtVWhwnB7MMaRhQnABHoX7jT
ilQT8nBnZ8OUY9CZ0oafrT/c1WAIGnnMR+woIQecfq3asXm+vTBzfo2Eh6I/UUqHx/PVgACO7il6
lb5GGFAd8f3v9jUbRcsZ1+YtKYEuWnrO80jxDTzrAl+z6CDgkUb5e35Rw+BNFZcP3j37BVJqzKa+
BlhaIT+eZmWZ1LwsfEy6gha8ooIgAG9vn5CEZ2u8XY1JTbestWgVfnjS5Ga73lepG83+UiVKm39G
ZoO5fJMfLn9Rqkvh2Bko73eX/xvI5GTj9Lu1mEvvruORrmRo/pd5fk0xJQJFxOC+4KrLI3D5bI7M
FBdQW81X4otas879GKEAnteggL06eqnVSMWQc480WjgvZoaZadIxa+FJbYr5l2Z0cwq4IOmf9N3S
m7pJzQwryOD9gTfwd5k5RsE9I5up7iVnt2SHL7iu3mDx47TMr8/Ng9nB4sFRDZiXzoS0Q9cD9qJ7
Oe2/QE6Js2PSV+PuSHm9cE2Tt4R7rM/gNSqjS5YrLiTPGRJRKn3O54sgLtshHIaneAQ0OyQxqxpK
3vANH81kLCZ4E5ChevF2r1NBwzPCaNs5GY/oHLn3yWedGWF+VSofKk3Gh4PyqWQjryNV6D7Uv1z1
bMnU0UEaQzDRzGRABpdAN7jX2qtwXxxF/riPVnO/JFhGDwB/LqJXo8D1f3ANNCeCwr0Okj4Z8dZz
sdKaAtJbOs8hJPwFCJqkgWek9oFZkE+OYkx9fYcoDeoKTv5+ELzZVUX9FQfTZqCdn0BygNFWPzQs
ToPYgpjvulZH/w7U3x2sGSEr7e0e6izpsdLHoH7EyXKi6ckYWifxJ8fEK38uSSCgfzexce7Z1EEd
MNa05FXPcrw9mysFxn/q9ew2wk6X3yCqf9sBTz4xS4h9GO7XBseJhqW8n1Ks6gsyHIUjFfQjXtKn
FcbcMh961S4cbALwKPGnwDRY5UhWNnAoHWp3aOLEr8oK6aNz4yo0Q965Wk/xlpPwXJ1xamlWram9
ScEZ5P75jQ06bBa7RkqUG3lfls1W062w2Cw3LvCBgJB9P3B5k6v9GcQKlw8EUBuj8REO5iaTGq5c
UtoG9RHA7wN+TkGz8gmp3Q2SYP0JuFrHSuELWpAeLl9wOKErido3cgUGB3YOGmv3/b9qdlvXmqnl
w41EHiCGrHFTJ3sazT25tZORSwidGeU3fEik1Nm2+JaRZNsVE7lbDxVa1qNQwfwTURvpqGB2RoPA
aWgkWOlkU/hmQ6CxEwKmNfRpItalJlXwiNOEOc8FxvjBw3MG4V0JzQfktUb1k+nRWad5p/ZiZ3jU
ie3rudOUdooHA3Ko7UPiehm71bCRk9kJN26ioD3JPTMeYgiLNkXoPiohn3CA4CbGUBusUx4RydFw
vfPu+Bq6CkFVk8QEMswY/taNh1xnAdEFgljCEwyemWoP7QLFwWqGZvrQ9+UR8tyJUOKf6mKjQCfJ
/He9Frrs5LKMkdDFkjcFwEueZtN5mVH69MSXEVtnnke+4cidGV+zTz0ZWxZO+kc4jY6vRZcPC/ke
mfE8Zpj+z0N1k6T+D1bKWfol0kfmv5DbnHFyYqKa+aer9sTkZV51IopZowZSSbExpu5APh4Sy80D
oV3H9bvfyT/h35SjiqhcpfyeRNxEd3UYvVWMEsiHdnJ2sJ4Aaq605Ln17y91kD2QGRLop4FA8nog
5ZaNIZ/gfk4+dWtGWuAcZO1cG4Gnzzb6lGdcmW46KgF2DL5kirzlwNBhJ/XW2I4fS5/o+3/vb7eI
ECJQ0eFWI6CLhjog5yIjo9gppz461a4QCr+333CwFPonwSwERD26YFyRmekN0AkkDhFleOGGii6S
nztNqe8PSVvWAT4bkjw48XrtqXx1yrM3+4AyKSRMENUvHZ1XDZ6SMHlk7a+JaaKp5OO5C4nEvsnl
m+Zn53nn/E2GLPQRGJLCBsNh6pzn9ZTZclwma4G+A4onrvpYkOicPaVo5zzzljtwHqbsyWJquyb6
zM6pbCCOJF0gRf/TVT1LVElkFhRuhEPF9qJ2+vT0EpvuJtE+0D+JgLReWZbfxfpGAMY3UHZk6EHS
GAWiVGT77okUMbsVyAwdRiEMGKfUdsjgFSt7XQOz3eszVI1a07/p4tNE5LsgT/io4NK+6SdQaDna
oLNRgtxPDq0WFSJjD7Fm1JPQK5gOdpM5z1+bo9zpzy52TRmc1vxeFZl3HtzlnH137o4Ah3aWV3nG
I0DS3r9JQs/7CVVXHJLhKvEmBTovYQIXnClAwCyk5fxqCnDTrOBAbXrAFz8UHx54F7bm1e6DoE5M
k/G1tChoxmt6dPRZUiZ3D2oBeOMAlk+HiNLG9+pVLxdsSvkRMvMDfYHmVjnvPt1p3NgLWu5YqmL5
W8sfeKzgIcQw9me8cYj1NT6Gf/0kZgr2BQFM4AnBbFMHFwpjI1S+tg1hGmgHl1tzuFjD2dlk1hz8
J8drr313nTM9bbCWUDQMU69DE7EKVGGDdVM9Wv4M4+Jb09feur4YhIWdlIQaYUMggP+6HVvR48Xs
AWCJHWA8egIeqq00Vw2j6VzxzRZWVEleC+epSg4qYwhlCiggt6sGRqM0SrFeTW2eXtylUVWylIpq
IXsEbU4VkrfVOM5Bf2oBb5dbnxuq2X96FfzDDHReXJ9tBiZiOsDdDu90OYTIKY5/pdxYSCpJphuE
WAGFEtLdPfbZvPhaN79rSRDVUzN4War4nTPjzmvzkDLUgH5ixIbHBerOZmfsD2j9dPnGQeDXTBPn
bkvP6UHylJ4tgux/HQhbsqoJqtdtkknb05p7Bq6UFYAazi7irud4kWaqD99CwSy0XAoTaITiMsXD
ze1pJ9dn1vVG4w0Vx31pIcxT+2g08TmxVCCWwzIetVAgJtfMSzzupKXicIfrBqjSAnhpubvRxu8f
bJfHi2WT7N/uALzZLFyCeJT4a6rJGImwmgu1eVn6YanGWt2WjJmB96iuAiEpAz81ojln/HXmgwVU
vN9v4F2hIQ7kkDPSpHCG4kFUegLBGKITyt0jrO4+TM7K1Vk3M1a/IZ4pekU2R7jr55rAMRERfRG6
JOJDZF05w3lDxAJhyMpyVzyGcwDGFf3QD1XvR5Pw9dgWbnE0Nii0JUaAWFgjABLqMkOB3HlZbVjF
X8T36DuiAF9Wugc9t/Y2vtivG0INcWnPxoyswb1WpshT7c4JeWmTf79W9B9GqRZFFHAaqCghOfWi
y4mZcPc73ilnHDnYbjYSw5dxry7gb53/OP23jtpSkjh+hEPCgpMVFVkfiuPBZ3IJYqp2kMo15gYY
kaQNCFk5fJeEhXjkE349lRHuS2FXQ2eam63xuMODmxiS71VnXhk8rMesCaJf1Zsb+Jsbn0r+3ZVk
57JhPqI5vfC67+5h/K1jSW2bXXca+1jEUnCXHaEzGHRLO8GuDhM52+2zKr8iPn1dJ63Fab/t4yjO
n7xDwbNOogx450e9e93Bbcos38aPk1MOR3M20HV7FMENaOD25lHaqc66RaaaNm+1gZ93nVNFRcgl
QcjzP0KADRfGPOA+2klYsvk7GQkyKFlmhnEp+nZGToO1irw3B8nnEP6KPVFQFPfC5RtP+6M5Xjuj
xCn7iieXmMq7IShpVTOksA8/lcB3i9shaxFVIpsjfX6xGtF8qdE1mtV8tGPe8cimoFJEmdCfqWW+
CWdGAmseyVVU8BK8DKfAbvHvU98J04At8iW88heUldoB4f3HInqssWoIs5+xz+HXvAdK7ViMWdHP
SZDS8UQ9/m6d0Y5vWp4qPtC/3scGPlCGnxJx5qPyE6XQGIGyT2aotXc7tdYdRb4TfyQd3lRlb9lg
AgXXp70QcFAu3Abm8jhnJTh3T2dHSju1ZqaXn+aY7k7JpCk6khEw/dqcZ7lRY8VXvLuWase+xqO3
0Hh7x5kdD71ZALnylXdQYopLkQ9jM/tWGBRTchve9JfBWNz5KCFDWoArwWF9e//j3RyFFHrFELa8
MZz5YU4fO9qNVX57GQ/VfYeBjawXOyRNR7bFM/sFH1i9XPgjhwR4/sgUbPNEw4O8VPgae1WGCpJs
nlr9Tvzq+iV3X/+u/ZfmPGy/S0IpxJLHV8RH4U1mKx9FgJXVA/lO28fvuaHpOnXyRhu6gyf+f+k0
JL5CFaQ2aCFFcd1O/qLNeWDRCmT/7Ebif7jUaT2ck9c7+kSDx9r4+uzI4uVe5xYuHPo4JGYCaNUN
M7uGtHbGh24Dy4MvAYTq+dHvKoejrw+4pEV8EKznD7ZPc92DA+8KhPxIeEqaXW0W5/ZEZ4CrpLQH
+fr4FWT1b2UyLG8VrmoozeUg+2ueG/BF9EI7h3xJlCi3BrvXJyCI7QTgkO+aMJFllEJLWSWvvjIZ
TqTQQg8HYsKiKIX4fFEftXHWef6HrmgljKxh0IR2UWrx2PJuSe8zsdNQlDitzfFNJXqExYhVSBR9
2ZQyb4XmKd4qA1CQz11SgzlkE8SfHnpb39+2ED7+u6X1CtrssTM7NnrUuJy8u2G5P3aswlLWhoGf
V/ObS1zQAwyDv5P+9DIsYwRogoOi6i+ivVXosgGAx3PHrl4zw+5NlUhxUfqR1/iiojpbfa1soRdh
BpORtlZh8CR69QkJbUd5Q1rC+wQ3JaAV429MoxNsTrMtbAlMlGCOkGdX8osNATWKAYoE2OA44aYg
EWaWXuLGmC2x2jZXoRmEU7xggRJv4TOd72y+k5ULTeQZuWZAmQfplfuGPXbOzu7Bm5y8k5mzFY6w
5WsH8WaY6osDYltCn+7t0NHjk2u6EVy8MTO+j7s/Hwgt02Dl0o0NhV2wmrlNYdOxBdEATi1tDI/L
/rXrAnkAwTNPk2QiJGxjtJzbUbIY/Rk3+7mOp0xD3E+C1Ll4chvItUd4WTrvs8O1BCrSZp8KNxlN
Dm2gOZpz9sjOJ/MbFN5NHBCU5L41JJqefdfX767JBeUpRIZabnkAwW3SUusiJQT7hyij9B6oUFF0
B5S39kzTtPhyTOcjqj5KhXcAF+NaRPh5TOfbHNfXe0bv+K8X7qUjlOR4SV6oEz0L0yvbO2P/Xhq6
Jc1NfKPe577lQlEBRg2oB+rBldj3UuYrK1Wzeu4+VdUFdyDS+l2T1X5sgJoWbZjSa57ekufsnrBA
lD1dSkRvDb4FrEOV7HLMG4+GF08ZkDYfQ9H/KlNX4IKtFJT6jmdEat/4JQJLubxeJfwAe3EpESNZ
eJTzhgUsg3Glaqws7zvtHx6Irhr4nsSCTpz3VsKEYnCPQ3jmvyLWsItJt6ju9e0LY0CbGtPl48cJ
VA79kj9uxDynYcdVxpyw74x5Gh+lmS5SSaAeO0BzM7vNp84Wi2qKQh53csaqmpg28XPu0fqOanvG
Id305zBgnoVAEtO6p1ZodDXkd9xfnx4ekgMFhVzkyqwRXA4B2p4BTEGMU4Or1dmwvDjYOTboxdjn
xtPXGwpzL3FzLuKbe1Dtx1Vztu2FPJW25riDeN5TsVre6l8qo4spHDh/z+V1dPz/VyiE3hQ3NhCj
HC0vDOcxHBYHiaaxjzc+bC5Va5yN/GQGm9qWqMD3z1RWkOC1Qr6UpT7RkSqjxg26CrWjLKpedRIJ
GpnwK8akR+tcAzuPHyecwhH37yAngauP77zNkvtFtLRlI6OCg8J0d1SgeykXw3qau9wvm778PWqN
xFrXhwI/QZiHzGYzvmPZ3jv7mcDHv6FPCkxfgigKz3KrqqKOpOQ4/1TgPjs97V7jvXZJk4PePOCO
op4yQbO/JTUavzcfnAakEeJZgTDZgib+ytPRb7iO4/2bBOAizcgtR0OnjXI+LxiRCob5naE+gEMs
IiPSq4ZLiMeMFbuwH9Jhb0Su57aQavSWaKPh5EP898KQcdrKNlHED2bEYLCpavwy1aG6PlWP70Qo
51SAWxp6vwqvoRZmHg9sxu1NF/zZJFeTB4lFNvI1Vk40ilJNtn8xdTIKK/Wx3Ty32yNyx0iOY/ia
CQ7FUTHNc4bRHIUHt1VYxVp2uv/hPqRCxVdnS06ocRq7ZtkccOXznEko3Zx3UOfq6a6o7F9Sje6s
g/Zpo25FVMXlmLNd+uwXPkqCxmKZPgZp1TY2ODmomHkyYlgUiOEX2dYXuHqRrQjwIn336467t93Q
VmflHQ1MTosDdaR0mAKzTe1eJvPjv9euSj2Qm+PYVOfs35Ilp1lyvg9VOFd9dTKIknIo8GCAQW+V
ozHGUTzgSvtkpgXG+VztTmWnK0Zlv1rH3b4xh1V4XxBFlGPsF/VXuEeH1yT5MuOsIu644PYPPJCX
lSiTYEVYaZqWr7IQIZRP4LX+uzIscKwbvJAcAk8HvKHsS9IdZ7FEnpCsm6wpKoiPdq3u4pMTZCji
CTfGdCzotmtvODabjFALulLCr282Yfa8olL4LMxfx8LaTEkpiBXkixEeGCOZn1x8as1pAmLEJI6p
y8JUeexqpgIGm8DDYOD92gzopn08CSJUwjPm8vqGUaPH9l/V0zQgRdeZ3n95AYXfm5Cby0F/P8pJ
vcQf0vZNsX7YUzuCP0ei36m+j/BwrGmxG9NFSJzjMl8Rgo1ZqahUMJfYc8cfUOfj+1CCbViYNbGb
VhuFM9CQIvHtK98v23Audch++ZW5LAdGGSJl8rEVnCvjUnUh/TGgRtD3Wl0+FxMtqzO3ezFpXJPg
uSE5rmbptaeXMCdcRPTVHoK4TjpEO7eSNNheX3DkhI2USHY4wqTeP/T7avmCMg0xDL1rDavmoN7S
h7PhI5YOCHITadE8hX9QX7AlW/8+kCesT6ZpfEv4EDtYOhHxlie624xv9pmuSvMDhO8qHhAYPk2W
LhSUD9VUS6l78s2aIFTWiSrSK25oVCfdrh7bdpxFDayxQ+6SmirBw0vX+mKSwxH4b8sGb6MkavT/
3sxouTQKS/ae4BABFMZ09bSby8hGw9Lt+UCMIkODGWg8OjQiiXugqcLoH0oFtzbCVKmRcRr/yNrh
yZxVvyJBuTshL7KQygdY1adlCS6KTeDTeOxLuMXpDpnfVQ+ELT3yANLW91o7OY133fSakxoEzKaM
h+hGpt56vqgX+D11FJDUmU5vDfJ+wY8W2O3Zc1gmTZ9Rt2nAkEpxjsWkbCBbea7Ebak2NLyvX2A6
wFq+lt+DwM+nHZzpGKDALsUWcXNjo8TY7pRw3f1XXTqJ3q7zK/zqO6Fa6GLNukgn3Fit18aK7Tkj
eC1g7w6Xi1pMvLkpM3oZNrhYJmHFyMkVONnqj5OXBxeixzon81QSdA5CoTMgYnhoRVQhtZEKsrcD
JUKvP9sDY6h6CUhJM8yv6tk8q0GdnH72ExhwFCRc1V1a+5C3/+NxCKaYsrZiHaql8ju5Uyq5+nyH
G+iKXm/+2HigAsr8iCOoGxR05JgMdYpuCPHzDIhP7kKIKVnJb3lMovX7rheOkp8RJR9TdOIYvN94
QTLMuCLtSyvZaaOBz/LaBRetQGCjK2XN4b2jZitqjVl6hxpMwAZy9rKhB8eASe9SorT79r3Fufta
mC6crVjaNjnkbacWKWo+LWD0HVa9Sl3SHZTVE+j4+6qsvufZ+ii3dWpAvdCPQZlJTfvWHWpoE8Td
9+rjwwLoNE6NaU8U+BXHXhPKEJal9PPcKX7k4UNeZMBdy+nNgrwR5DA2pPSqhfUPAruw+oNLunsE
1kRkR9/Gq0li3pNtwgEOxzhb7yLH8aCOl7UQj8TMDQW8GNS1QwBrjDyhW97Wz3IPhAD2eEk+E541
CRFvsukXf7KOa41fV/xZ5W4p2Af/s2neTIthcWaMBP9CJtLedngaEInd8FDo0stNv4qrLsOrMuGW
Dqqkwp97dWGyllPvIdSv0tpClhWsUOHQyZWv++fUsSPgvjVhiP8CzJWzIHFxU9tAPPDPbMrDm5F5
4hU6jdwOveVqmrs38JSfeZ4r+DVICJgHMzuXsLcAXtCO8WcmAM+yB9ZYf5aNGgXTllqlwmyEuMsR
8YzZ5iOlcMp76h8FTj9Eg9ubGhfy+JUZQQWdF0dLozbNr851kqyVM9JK1mCGlCq6fdK8vrqblstD
BLoNw3eZ3hVdBzaHRHhnbKuic4mUncnH6HPVytRHJBGUqtb2YI162B6PTabxGXlMmDNmu16nlHvq
Jx1hQuCS1oKPhz/kP/eJX8mjaAgczrrlyQLgqrBQM/KMmDUmdrZHe/V2xEaGdgtqyVBFm55oEC7T
c8EWdfHxLCzWTDOGGHUG9KxhJ6QzI6e3XiHIy6SkQUJcJzEDhx+bQzM2TDIsRLCK7RgDkJfaWtJG
cenj7ptofdEbTPxLAFBT2eBIEvbw8vCtq/xe1Om785hZ/Wc8WDqejaIZCNPsFDrLyEdQxRI0+t+3
nLqfrlndw7SHPVs7CFLP4xB6qC8ELpH34a0cjA3IdCzt+qnyUbYeZoB2XkWPFxta02fH+0LVUMG7
B7lK6f53Y83pnjeSpVaAqDySgPkaqJ5vag48ree/fzclqw2LVnTvHnSunVSCtu0VgrPipwOBfRIb
g1PYiSb16sJbJHlJyKdagrmszxUSKT/+JvsmVRxkfUehwt5QbbbDkXGE56Mb09hIn04b9SZsvVfk
LlUKHNuJZNtcGeWhIgo8xJGun+BAK3mFk/SwScqOso3JY0rl2GkteZL01lgqSCGiFZyLFw/Hyzdg
e5sLzy5raw+t6DDDZwWEK7/MZ/OuwiadkDbMTd3x6fcQQC5rZKyFoQ/cPoVlgFsxp9saRexChRjn
BRV38U3tRW1GrdPSJKxB6HnicWtE4Ah3oRGBlZwBLYy6S+S7S/fLSTMra4UQklgAA30wF+ShaZfG
3VSs8/7pzTiTF0YIZitUIbZNxeoFnpBioe28DYHIZfmijSq25NSIvNcnbLftNnAw53OdVrujCpwy
S2L/9tJQVI5mr/f6JjKrXBUxYza7QAl2Yq7jyFFJOzNDuRMZffhgVYo0xd1BccfIuP1JRfh7aDy3
AG9+TiTUMro4t91N/1ndqbCR59cyR7+O+yA7ZpR8fGKMeUC3YBH6128Pof8tlGKkx5PNjl00PkdX
GvDarGbjGocQC+8676L/j0AoYULx+w8k9DMHE8NWM9vXFE2mTuJLRUDWgnE2J5Pp/r7msmUnxVa0
UpZQsG1a6mNor0Ty/f9GRPxVM++RJr6mnMu0VXXluU5/EW/ou4wvTRJsZ0Fcld5QpIVvix9PCnhI
hodI3ziX945j5CF0dPz+ukPdI2EYN/4LBjuZQZXGgvu2jY49AZPtN/hhXM+Fz+IYZjPrhp9gJ1nq
VNksNyKzNwN4JGk59I6BYLzk+eHBVO80HIqRip2SJBAHOFKEKRpsnagb5+VEEULK52NZWtD/P1CU
387tpHXxdCQLadyiFb9OUHpN7GYQ7ou4WtjeAMNuIsIqq4XDJi5DOsCZyx4E9DbjrfGcG2zFomk/
I71FbgTCTUGKpbgkwL6LPY0bj7bLbvT1SbT3cOfe36LJ/oXNsq3MGZMH/SlgNFjJdHvQrFMkdEKR
jLfDd6mIo+qSQmO3u3C8WEaqiZzWbr3fuz9UQ+BVUl0+bvt/7cgG1/R2SmsYeApC9jtyMbQjUI6g
pqIkCgzuXdOmFpXi2QNVIycqZvbCTMK3NOQJlEAr71ILnWLTwnZYqTAQUDELGoD7UpV0Ydr+pmtZ
d3VgMmcUdlrSYLN0kv5tGH2ZujLHJd7t//aqOdpXLMd576xnwDR6Cxz6gSULaj4mO54f/wHN+0r7
3+2ym5xAauBF41vf7xreK0+i7hJc2qhVICKQZFaVP1GYQyFK/+Do+7ehPce87RlYZoq/vpRhXa5D
nXmrslB9JblDYLtzhAkmN7dBXgEc8agx8wBCRW84+R+TAs9LjWSFEpFdIqwFdpefX/ALGLoThQUO
DLEjJxkfe8FwpurK/RAarodT4JUt8LU0i+Yq4J4FHbVDSX7466uTlxKHfI6hx2Gjs7ZC5htDHbIn
hLDEj5JIoFUfJyGifbBc10SXyV9TG7C0ZV8PWdSLY6bOxL7RfyvwyRn8bgh+h7C1fAzMiu5sw8r8
ECGjXVsxzpG5t4yJSu/f8Jk4qsryLX7J9Vzz9ZDUzWVVPxVYobW38f3pu2o3F3HFrQaKLLLqNSYP
xMm1hIiwMp2blw9dXywLaZHyIIGQ35c59oIRTMZzOHfg4twrxRvNcW3FJFYQZ0FGT0yMzkORJZun
a8dukdLgI7Fbt/eIg+/1LsGEpQswm4MXjWQ2mGQqdnhSiqs9VOhJGkdWVAk8vnkxo6YC0WvUGDcn
t2Bbcq5tJXCUkrl8Ieqz8aIvbo60tUiiCAZTFgRvZauS01NmoyGM9ku4Ixg2cwU03B/eVE+c6L2h
dcGiUXYW7TmLuVu4GNTUQaddy9EO2xgNQkazhxagZWs5R221CsnUjZISVQw69ntBrX8DnBF6uEqe
J5+Rv+mdEuBhhmTUxVM0zcGE1/bA+zVjJPZjO8vqkTZay8BMiBgZfUT8NOx1aW8IFBDDrcqH7gjc
lFyHdsxdYN6LzBcRp5NozeYOp80IJHorF4adqWrsbZlrSstjWbon8hIGZx2nLprRv093Rnm+6Qub
aG50xjLZaiw9o6pUTuFQyX+z2nzfOHUIAS+ecVxC68vuNq1DGK6F6D2v9+yo6Wqurvf5K112cx9Z
mxaRB2uNWF65ClbycNShew5ixa/x8k+UWSmzzu8LXjBV2jrDWImRaVtxn5cFnRjqYWoHozdS32sx
e7GAbjs48wWf9Yv70tjZXf8qYPeLZg39qK2U1Iv/vT/1uplGw/09zmJnwUpxZph+KI4A5B3vgtey
oyMddsfPFF7vUuIuYAgybkMpByUjFjUvLl3W+deGCYwMFtatpnhbpNomqyVnXfiGYtBGnSansCfB
1ZH2y/zvCxTYJL4Yg+P9iVWqcgFFFy1+0VXgkkvPA/SPos5GySjJqJH3kfLfvkxPcUPAVDgHDiCE
9gaUaXFPd/ipH9rFKZHLKXVzWYr/uQ53XTQZSFrxph4n+jcqKqgEwSrV8RuWvrIuxYfcWOmCfjhI
5tcmLRYWXvaPCon6/j3q4vLahIreTmEDYTCJI3ZmP6fWLSwfV16cDkZ2H1YeBp6A46iDC98Mk+qX
0T0bN9bOasM9F/MlfKeOryaQV0BGD+026YTtCqTRSEUAVqg9VjKs2pPX/cT3W4TFSxoQNmd1N22k
EVJpJqnSJ78t2cuIVIceaFn3im8xKzAKRCKhyqb9IGTzMDaaoACtgwa0l8619DhIHyaTCew+UU85
LdXsNfvZTVxhhl7b6WnlkvwYDXZCZw6Hs3I0CQqxLCnjakJpT0O3hUwWFLJGnZcAPdv7fVkdwxNJ
pJB0npBtcq9jSI9d1PodIuMbvyAnCZkgoy2HrFWX2tSfKPCK20lRM9Zacj/HQwB3qIZVuUqoe6ip
msd83RerIC/ZLIix/PWnM/7evcZxL0/u9a2EBTgWre7sJffKvjHBcFxvmQ2M4xnS8ZFWn9kYFNh9
N1UIkxY+X393ZxIeRCD6Cg9nOBY6oq7mpsuxX+peSiKhr12JLclDxDQ7vSSf2xpOcEVPOiHiwXup
rzlt8UElcsAde+P1L8km3Wvq71BZTr6MQqGdv8YXrMOkqr7/dODJ2527ulfflQ+eU0JbkYIa85Sd
ytvd3WybXdEhJtVspEQO/91colOwfEumjb28xERTzEsF2XRBHwDbPQ6euE4fzqWDceF2i8/UnZoQ
mONboZ2ZuJ5xrGOUwabD21bLp0cSDaWQvXwE6Qxj3kS0qTHchG/quhiSxkxPIOKQOecC4iuwoOFc
wgYgbdalRpZ3aqd6BcgvOA/AlM7qes+Gb1Q1n0QcW2jFYh+PNszndijI4MuSkGRFrhbroj1d1iyH
nNfnLgS5ix9g3yyLqUxqVL27tu4vpcU68n958LkpZ9WddIJwca2aahHWEXrCR15h4GCdA18LrT2J
qyKV0ZnKGLz2KzM6ZWeo+Ir9Rr+evIYB70LCDwRRhNQ4C+bLpNXAyCLp9Kp1mNu0jRtUdVGb6ebJ
gRiIkE7PoI9Ap4xluNkWyI/OnoemgjIze5J8yme+OC6cM36KNHwjIaQQNng0plS/xDA80sqnjjqN
odZx8EtHXc0qJya3oAAT81su5/Zq16Oru2pjX+Ime3w2RxGjOyWfv061+6BqqrF74SycyhCrhgh/
DkxEHKNBF0BZVlf8odYG6UUZiB84x8Qxzr5/PxjtqtzObvdg6B9MmAs6dhYSHCOzrkCf3UWKD7CE
uRfGSRknhnEeZvE0uqtN8VqKZg9Ze6iRDyPaCQcZUbFEXvzrSfUSf+2sHESm29+SjCQe/uMfpIj4
Z7K95FcLjy2OJIQfjm+1NpQlWRc2fCVyQ2P37Y6ANpIOdF2ZcrIJjas1hwsq52A/sUQMBlb4qKnY
vdxzMeB1mZgz+FF381uO93muf2KCBWa1b24wMo7fMnMxnIpDZ0chqT6jMYog/N0KmqjYK+aUOXmK
A8DLSZyLePKe8Oh+GaTqoFSGin7ZxXxwEltZo0AEIdIn9ZIhtSs9xYVzmzy+jzsy87XFovATONvZ
lLOg7hW7i/VWsmjl2EdXHCHghk6rOHMrRqO/WdQmlhFZnS/om+aj9AJESZXuibs2F8h0TSLNHfSP
n8cXj/zzVeoaOemB4As6xcvx9yYF/BYAq9GoTIhasy0PdXkVyAu0g9T0OovmvyQVz52CRzoectx6
3jxasWnrQ70fvkOJei4C3VMFQMruEp04qIDfOThbacFiM6NhBb6nv073pu1H+7hkRlUgJlpsszuH
idIs4DOHWHse7f6i/yT68oX/oib/dhc/Xr/eQRR/9RWRPEldRLAu3PH/HTgruCMwPxO+C8Zke1KD
veYIoMzGiainjEryUVnEgg21zxLDxmJJFKycyNLkI1rxKniGd015zSU+LMrBvO2iEwdFKihbvvpl
vM0G1Wd62/fjgd76J3Bf9tpzjijlnhAJ1sk0xjUr7ocwJHFsPakKFVO4o1Uqm9KXfpphiugPc4EM
lEp5BZrLcQtIja6Ow/dg2rMd4KmlqctPqN7PiwPpyJp/mFV1J1eekuTIM7b5kU+p9AqsrcezL7eC
M1W8vBx9cErAn2YKiHEDLdRlgTYVjtKkvDNNSDhRFMnIi580F/VTlGyzxxABODu8iiUtXR1r2Mzk
eUqnKWdkY8ICqMbPLxCLWi920tpLlbPtQ5BjQTcavVGFZUHYI3FfKMqTaVVqgwyzU2ldnTIcYAd2
1kcMl9d0DPsEOB7SucL59dqwzHzRcjsNtxTBsJ4o6UMUvrnsWR4hf3LNJxetKN26l5QKXsuEnOmE
Abdbgb29rYDlQyeWsVOHkEyUaPjdBtaXFZKz1t3QDr8kA9lcrWLdoP4DGYSWrWF8dyLPraOuzQyu
4oBRXd6KmwhH+1Dw7QP29ZgfnR2ISv4SoMI716ILt78INdK+jHeCK2fxPC49QZj7LrTUKxxwID4g
ytFFBFA7N1YMyl+TeXNbcrzXGeY33fh7BBV7ZzxdjmXOTx+v0TcQB3V3mky/z/66qsOhPevapwKO
9CS4AK+wqUUMwlr5kNJGH3QlhYxF6tt6kIK6cL3omGjdIZEmPVzmMd/AX+lYtyk4DfI5PiHPzlBf
Ib9N8yaw1EgJeUl6JgrqGHdfncViuf6+6b3nVX7bsiyEYVnpSNXkXbY6jV6/eNc3lLLxO4HDWwpY
CiLIPpeHwkq52E+GgC0tfTc450YrVqclGpErGktqSEykVokwV72CDNXUM7ZMhPRZ15q+nJk7j/Kv
Fjh7PlZbp6E/yo/RzBVCUiGFnbIIjcggJBI7VPZFFs76SZeAmUbLdMhi8qz2mhFhAI5FlDSvJ0/y
pUIEyCGYYBUT5jZ4C2zir/0tJV3ystM7hGL0DpIrKoIBiw8tF+QNf8PSV5ibG9vRuvKSpz8swlAO
w+KEPhsqp59Y5tCAz+0hHk7s8/jBLERQ9t6z0IA1iaXbWI6i40+v/UqvrriJOqIgkWW9tcHSRT+D
HOay56DwVp0Ylv906KGaZr8mqQTQLb0JND9QUUefq2UA5+K8RPzNMWuCrq5I6aMI7SpxwkRrQ0qG
FYtWVa1/QBkrYHo4KmgnM6yLhfvUpGGM6h5wK0kbVgXMAoYOhRg1264D4DN7LF4NZFVlOddBKRiQ
5tYK5bSlfZpqurSwXqoKNyCU+izYVrd4t3D1+cTb9eJICM9aphLnmkhbgBPkFrLuMKe6vOcCrrXy
8gjJrvB+/eh8BeJqkRCE/JdCfaoo5Q4VdAviK2QYazw8t50f3jLD7/Kf0rrIUoqSIalT7btoO16O
BSgit9/3Xkab5XdEUZujNRO+RQXQsj5MIxye4XSgqJrYv1DAh+O0FVGMYzfQUBFtI4iFzzVhfD14
kdQxQi2hdFapQxXBD3Gy6OVryYjG595PV4jNkHhxxUgyvo7TzdkDEYuLIc1TXz167oEfBVnphZcc
qbzPDI591uk4DAPsNEsFGixvbGpbmWgADnvs1A/pSq8iqLHTLBtf+B7x1VzJywd0bCy0BXQqrDaC
tDWfSu9+x4bes5oN9xQGAB7/A365KFQF1tBb8EcqgF1EJ0zahAh9ZrhqZmg5L1vjIYKo8Mnoa++K
pZCJJ0yGild0GOcRWNzX/v5XhxAke2SCYMT2nN2LT+kwDV4COk2JfjMJyirOc8veRV5lxgyUK1zp
mxgjZ1HWHt8M5T/YEuuw/WVV7WQy0qNFYE9ajgs41xszBfGiEfhYpDq6AykGzkn+kY/m9qJzXpTs
mkIdWHMeBkGpFAWHjTObw8MsS+xf2gqNfBxYOohhJkXUXQcSqROcD4EQqmJvrSLCq80BP5wbTlkF
z4qsqfjILuDxrgfcQebpRI6zZDt1SzFiNpX7UDrAayjcSb26Gm5O3F55Jyu4XLEgoOFQf4M9RA50
B/AR1d0Yd8onVS1y7tz0gv/TXr0SiKBHrU8JWZHRqzBKx5/9O5X738UCGB7zG/sg9Ypj7wGoA7Jr
/7Sq8sP6QdqibjUHHQO47YwnJbykRzlUo0lhWQ8D1g6zWDu9qOi3JTfy9y/5qoamt+dTCtfXGAxS
h+zqgSoBilk6nsJv231LJ2uTBut+LFDjuU/BLUOtXE2Q5CC6mtRzYdIkeBUgU+CtLsz+UqbWzrTY
ugPsQuvoX5ugB8B6tINrivt2ZQR4qTY0NXt0M9Hi/ku8+apaCGRCYfi7sRZ0zW11Km/ZftejIlaN
rlOE5U0b9z5U+Z1cx5bgxMhY7Yzi9uXRCBh8mTDpxj1/txQJjMPfD9erYL99TKA1IgPpaCHs7b+8
MkJO0i9sGZ+xPPJV2oKPcyE/OnUXu1kEyGHTZ2CL72ZnmWUUBBosPYpiYeHx0OdyBcTS4xL4rvbR
QddpR882TGBPnLi/o6FcAUODmsr6bBkwQL/+dYtbnjUxpF3SSSeAcFvcZZkxgNtvAx+dcDPMQTAl
1otb/a5uSOi7LFtaMYXSm5bZrtZEDnbGTY4/9u93P+hokhzOmRaZEjapUerwTxTUN7MwhlvGdeVf
BPZ3ARdPZFOPPuzjTDk9NewX7meLmX27s6aEcMYnXFGc36FrVbQfKD0iLr66n76spHiE24M5g/aR
mhlU+gAk53aAKupy7U3TUfj0zSW7ANGRpbr2e6piqKVWm6C0PTkDSZbzMvHtQz05KgLbGjdUcNWc
kw3o1Xm8HYJxiJ//1qP/c6YEvkdSvkSQ1z68FvnhJvaJfeqbcR82ju2ZBsHcFvrCqBaD2DQRM9S7
YrlHRggHKZxmyV1sKWnRPdvsPJLwZJeMldt7l+eLgurGq9RVL7FIg6Y09SRrTsI2Cph5o03YKAkX
o99M48sgpO76RfYv6r/l4omvaG4mmAGC1+JyxyoEUOmQDmOo+AHFO2NbSdBWJhspzED6btIMUUXJ
iwyjdrkV7ZtXeHyEQyzDW/2bQDFsa7KC3TW7XbdxD5E1Ub7mdkK9FlG6qY+dpR5lC+W2sUwpszja
Eo20ewzmsZrWAuJQ1GS1QTQY7RDT53K8X+5chfDIlq2axe8fa2JuHUHtjGbg61sUYGYjMHe60jPM
ktTGYh989U0tifNzCbesMCjErLd1Pcs3HQoCD0ETJ2PBSsWMr41BJO/I2UGC4RXvARLp+7wgknLs
EUMJJ/9ht3UBmn4gMztjj02lThefe1wG6xr3TX64FVb0lyuBWj8GKfvQN9QUX/1HiM72Qu1gM6LJ
U+ARSpEb/Qu+TvlkTBdI0qVRd2QvfLRW5AOltRSyNlRXaPgGHmJJ/poSOVjcReb7zagU03KEqNx2
CYHBWChvaMG7cX05mMgYLuXCnyY13MdZ3gDUz2L6F7NUkkxYfz4l+1Ayfaf2ZYKQl4fTmO0lhZAH
LGnsgZ0RJLNXqUCqp3erBwmp6g2xd2RlmkECNJRmXMKNNGpX1MWfSNyzSd//1t37cqkizwUvwdfY
YUsuo4nnT+m2f2Ge1jxhiQQcDqcvbWVa8of+bA1Czhj3Ek0xkjFKT6jBVR/ESWQdRIvtgbZFdfj+
xzQg0V3cabTgd+Y7SS79W2Ra3YREP2LTjYR4+bzJgVmKq8SHOsIpDZhzoNVn/Kk2/oC+bZMMLYL2
B1+ezaLifs6rWzdB2cobLEsFucuC7cGewXoSEJsM36LN0Ezl+Gb5P2AUhx3kApIdDaFRD1nIb4Lg
TrGRLOzy/PCCVaR0PCbmn/q0hZPGb+Yp3PGZzRf0Mgeqstrgq6oRi7dXcP1/qEES6TBOOrrtPwM6
+RTwvIpVERRRafXYVqtpLZEbrIP+ACqOExtZjGcDltj6FLpIQx3Z04PUaWLjZyOL+E14KFLOcAMV
MJ9So2v9CCKDDU13vCThQ0kH5+8Ag1+V6KxVEHirxWdzWKflv1rijUT3U48ZHusrKfFJvGhN6xWH
X7fmdA13zbwaYqpDtlj9KveiyB8Rj53Qy3Y6TMASoAPOpYX/VK+QhVJ11MlwCIrdWfO/AfIf/UiQ
cwy2BbiN3It44Gspbxfszl5QjFw1HEuK4rQ8V2DAoIg7mG4zMc21VOmMoW4tGVKzSH937dB5bRqp
zhMJRJu4qW74Y8Y3lxO7NEzJr7moBMos1zTZw02BxrZqlbFCUD6sD4s0OBPi5mJw/eNAnhXfii6t
92l3yPiaH0kqveVA3tRbXcXaPkqBZGpdpbPLyCXDSxvl0z0BRWc27LXZYXay8dRXBbanxMxLIRwA
pSYMuhY5c9avBNG2ukzjZ1NvNlB+DKVkj9q8TgYJ5GKclu1cfpUHC3OfCUFs0cLtdFJZJ9ZNE3/x
EIe2TUsNSRbAZ5EyzWWNwa2n3CNr3XGb73fldpss12RbftSTLGdhy07k82FlgAgA+EYofmP8iJF5
tDcY5sYp6cj8uNJ3G/1EhDyffFy2cF3sV5UlwByvrt4W7LCfxGiBdpMy97o+8Vk6Jxy3gGQdNP5E
stIw/5APE34x+1ghv2Iy03PxDLX5gkdg+UXsKk2M8Sf7EDP3KTZS07+8c+3OPFW1MRMbxxOg0T1M
irXkZOzNq4d6fO6sDH3CUlVfR9AwhaSvbmWgtXV7iP38+3bPNMLaazR1kTLYAdaT0rCaWpm2Iil8
yCmEJRCc9aoWLn5m+/Ipdah8oqnZvRbz70EIgleoq/DkiapDf+fZLS9/cSwWQGUTpxsxKizuRDAc
ic6GVW/vIMJ1pcWNwjmQzBC5ZdN4Uq9gFNMRTKYLDjFSPMlpBFXR3PVkjgKKnzlTzGLxSF7g8ic1
eEoz8JX4mt85K7j7FGTyG952QQm0Na58ejnd1MXR6DdalGEY6BM0AEBe1TdVu4r4mFJxRRvMAtqn
Qu0pKdphm6KW58RAERE9Fybkc3H3m/EmqjmpKNtaxZjIQaRMxI9tHc+yh6ySNN6PlVc4OsH5oI16
sLNCg4t8oIe83d5BzOw7uhaXwH9TlFdh47imqVdegIRI+VCsdq4mAwrIBeWfybSj6s42aSZZwxhr
i1zqwzEXj0XQq4sHslU7d5PPdBOTZ2cghoSQFOGo4PFQUXA3S6f49U1XsvjRvgfoGs1bygIfJ4Iz
fQu832MxqzmVeL1fDS4npNfzbH7jCkzUVnlYIeXkYXVs9EEyb9dd1QbvTqTjwAOdJ65ZKc9TPqmE
2BTTkrd8naTeuUiA7Mm04W4+T+kdrVvHhVKS10om9HidhKwUpLYzmGXwZ+sj5MG0L+ZEF0vabBjo
lkseUzqMUd2Pueau5YtUqBbICiHs+vE/+3B2cbPekK5TjdwLhT6JGhQWGZBbGr8dyBtHCEJhWphD
yo7+ttDGPDOWMLZWbkkO1+341r2XTQrN0rUMjqMrs6EZ7GBY2o+5QPmnmpZ85U1scsKlRuewoxau
AouMVzjrAo9FO7E779yMyiyls0w4P9kZxiyffrmuCTOvr5OfvVh0gM05avg6MzNgGFbxOdm5T4oW
m2gto7JxKOxDTUtN7BXbKwtXauaXJgAD4fCt0iWf/+uUZRR0EUbIrt3hxHRskFzDS7Lhj5iwfn9d
0QADHfYAzi0ppvxdjAx93WExEbPZGDduQQ+EuyWhwFYR1ASd5aQm14n759bXlMrRSPAdMDPSFKOL
/qGQ0+R+WNND95OYUoHVly9kzIl7tjAaKUNMZEMOy9u0r5lrGxQkOKFvolWfRY88s4ZCYSfcyqlO
v/o9q+zNfvPOSbFgZATf0eZwXk0bbLwJwVT8i8HtJ+QwE5oSwPyCw5eOOQRL06LkTGU7GcOoGk86
FNNvzuhyfM3bth81sE3S+etbE4jCjpyMgHvE37gvrNqdKWH1NWNhIVkFZPTJkadk6tbZPiBoPAoo
ogObpS6fjq2ol85mDOQmTjkXYSRM9ThMeLBKyfs114yZHV1h+YxBotJj17CGZdT1TF4YGQnIHpri
UL04FzCg2VrzzgaFFQYKSCkYAh3gz0s0LHixCOJj1oclfPGPRRE6xHK5hRB9flATmMJuHdQo5Qsr
CDQ8wo5dqhaavv8hjbss93Nd4RMZppH0ejk/Drx99IFg1gQ3Z1lNnLCw5svUjwgsnwfiToe9cOt8
4W8c/TFhesDr5N1kvaC4TxtIXYa4erIhZX+oY0ZbmPzH5wkBg4tMBfdD8NERLQLkYe6yjrcnXgGt
X0hvdPUt1Q+AtW9fC/dpKFWjevhmNd5Hr/zZmRROwwt2MYgqAq72KQbjFBWNRMUp47A5BXtT9qpU
4w/uhFI8SCDQ9r8tGJqLjdMnDa03gC0C+PhOrKqvVfsS/pypEamoJpAEf13Z84Llw5wkXb9OgNFW
IwYh1TUKcKYfzfJ8xDRrSvRje0C4O2j2NptbFk8WXSXikMZ339fwlyDzEBTDx2fEYVtRX+uZ+WSZ
WVCpwUuHxX38lucVff/aXkpLAVygKjbp1ldV8RVkhiUFezcT3EU0WOLFLqrI8KT5DMtdG3TPrV7v
OU063jVz4uZaB34OwY4fLnln17urfYITpTB1jrzaR0jgH6UlMI05aNglSeOnDVfLGlxh0abV6oAx
iS7Jc7HaL/ZBHYHdvNLQLY/hiYH126mCmllAKmqtL16K4tF3lDPqOBVTWnrYLHvdtLzgWWzfZhmN
ne1cxF/FliBUbzPcAYX4gLWWqkkTSeuxqxvYEY4O9hbfLEmzE3XSFR6u52wPMJQylGmEGujTJTDx
qW8G0kBQlKpmpy7fV6dfbmy8vCGEHfu8ou9DbVt8SN6dHpLeJTu+5D6yz61cmZSIHZi896aBDTaS
+OxEQEot87FU4ZMpUXSpcc1EVHYHJm9PnWBnNcunTYmRRn9XifbLcoBubWsAvNYQc/PmxM02QBoO
BiUQWEUKLpto4DMsJyY1ExWtOz1nS69R5f4IRMsROrW151zVkMSuLCIiw2UcBliSL++gAUg3mXgE
56/moVitPu8NHb9ZQyldsK8zEB80ThDpFUfSkV36abtL0KS8mLnScR0zPhxUxRbMQinf+xQSwO/R
PeMudariaOfM3FEpjoOuIuPMMawWvCqpTvI5l596YIXn7VbAO+5Fuzmqe0CC3e6fhB1P/wrDj+Pe
0yraYF1ARbNtB+oZW+xcQRLEu29ULHiBC9ek3Z/61Dq+15KcCVSOt04ObbbAW8W26EqjoflwT8DI
j1n5ysCluI9xl71aY8aWRUt2xHLv/7xAIhnwnxueh4GIC9DAKwZG4sH++V6f3uhsq/0Cf09Yr1El
GGgmBNTJgghbPrpOijdzXDecOwCKKC3k4O3USvm5xQDycxNBtOvYrIMyx5MMUO0UOjiqitPDWK+o
zAU2eTcxVDPVVmWqJI6vMqlkRTUhiheUsYRErZXX2el7jpWvBn0cVoThwbJ8TQ8FZvVRYi3sblBw
QWfEF7gwItwTF+vb0wMQ5NX9JKgmXQ5wftNQL5Aa6LFBpS/xEvxwTWXjAQR/6C6fMyX5T7RdsAMR
o3KbtwFTCCn2U0dRSZ0LdVUlPmzo2iMbil7NBBf+b2VFPPRH48D6lpQp4BYaA8XsDv8GSQ/ZMoLn
67AJ3hEpq3qRD9GDYx4wiIFLgcraTGNOxmLRubgUoM3pFnHzyXTU4Ie2AGF/JIt+3Go9Bz4THuGH
jQbNZL9hTdeN7wM0eGXpWbw9kthTsKXC8x82jfZw8ZJRUJbjibS8CwFNZIklV//Z6GgtkX0xTI4/
1xrXYZ0+Ye1MvKXTVB/CIgcghmtEJAJ4OjEYJvULJgHp2gj2BRiH06EhhxTU4/yHA+zej91dJB1l
94gt/aB3voGAjrIIYXTBFM+lQN3eOTlylpDbohZaUWo+y3O6dLjPK1qnqSEEesW8JhEtiSHzeX0p
SqGfrL9V0thbAoJtl30tbwNFau6BUqjYNZDRaMbM8Qyn9R07ht0MWUVIlCo6RPVI67vMktFqgAsM
jLW6dOLtwiYuM4Tk6H5dJGvxnGB0dctVzR4/HZHe1beBPcjyWo6iQlenI4OKkMv7B5jIII8L/a7P
ZSzPLok1A7prNR6hQYnN5eXRtDToZRVcPsgOORipeAekuo1SPkP34G+ri8yxLJfGqzCcz/rTI5br
bmPrAh6wxSwwz7h784ALbDVSfYZQz1Sui3aPV6WX3SVMBwkkyNQV1OxknI49zc09M1ObpL8dE6Ft
RKPMM6/aPNO8pEuux+3oHfzu5GyfmcWff0QmnE1fmwkbQWjTO1KuaCJs2SOC16gqNmplepDKVBQF
ivIKsXxCi9JETwcqwPDFaDxxYOsRR5Kf8z7+zbpVTm8xscVRZRNGbcYIqaqoOnc/9qKqQYifhY8O
+pfUhuYKrbFw8ipDRm7IgqD5H3icydnikuBGS0sO8pM7e3kStNmPSH44le2w1vXP5HjVD3Nq41sV
MyItj9nvz7NUFNCxe3kl8a0FbpvAoquq9g/Xf6taDaJgDwzLaXpw05rdkVk8/U3YJZ8kpmPkfeQu
8TsLLeBVWvGE9+61gcdcuuvuPGp9g2U0+TqLrueml5bdk4H1OklCtLY+jxadNFO18RLuKZAlQMR6
3wGb0PJrSltnrzxoKTEyIKjSC7xmnrsSyp7fIH81ggjjIhV0aeADBjc340dYnannsR/KSNRpQM7R
kkDshILG1xmcXw9gCYtK/dM+CHdAAB2Y1cjT1jKgGxGGgtzVKVGyvP2xjrKErxETVzKYwWKXNiwN
VzWcW4eeELVtRrL+Eb4tF/fUvb5zjwzZkFSUtBG5KlqCTyj/m0Rzd6xsmNJ+w1bPlmIRw9r+jSsW
3d/dVrZjcV5j/4Q8PDWgj8TakYIRkMVkSpQLdqyhVS+/bkNjdxIWAc1hRxq4acJrJbuPvAJdxURv
CWF3U0CuVUyedG9pDQsMPhKXzH2ckao8SMY9r6mmJ7k21qvoZkRXp9wFGtbFVp9p+JDOAccN6Lvd
zCi3eIICRopiYpdg3jNUunno1u14ORVLJ8lnLuz/PD6GISB/kY48TTq+/PZzq9aGoHboOC+s1YUS
NG1IQKUriW5MKhnnPMLrFvJSm+UWT18HVrOx8nRefnOBeNXMcAAewnCgxvRk1gNgdN94N4yAX7um
4HeiMVON7h5AZ2h8ZtVI+dniT7zTVVXB5sHtQ+WJZAe7gLAdIk0AOnbYSOAZl9WWiwarHXGcs2qN
m0DkzoRsMgWwxVK39JWBSSDAKqj3wd4CoPgm23/qvuw6SAcqvrq0RFKaRkbGqZ8t30EPjKiHfcjm
2zJgllIbElLkOTwcM2Il7ublU1jek4qV/SlC7oFbdRqlIW1Gq2B1t/Nj8tNcWxHqSFBHr5Dbul82
O/AVkFHVHhxch05uDopFNFKj52SCEiwnQ0lO6o1p8AlgOImexWRZezBD4XA9OC556SVKh/aREJbQ
WOxTLilyV56Xgl6RapVJWWdMVaucDkYExDh9DEsNEDpGZ31hJtUxZtSagIAQmfDs2Ub4NEcEOkcQ
QWuUgr0kvcgpuIV1AFm1qByaS+b5+6EsSzwrnBlikvvkAh+NdFahCICAHGLfbNkdcm8zj4hdWG6u
8k+6bWgReyGSrK1xa4ZuhtQ2NuXsfk4K7bfN1NzbWRy08bCe2YQROgvCPcWV7sLVLHOfaL115h+w
67ngbBjSZz07qJQ2B+GuKZq+qaZR9TD76JuoubG2AN90tO5mw1YCDgDsmbM4kRUFPcuZgg2vqFKL
7EBYj8jISY2r/FDcBL2bYb0YVK8aVuCbTbPfy8TLgpCeKWAJrn+W6sa7Tb8VHcCtC5bIqcGu31ew
oCpN7bvRetRPNwz2t43cvo3Jm3EIRJC8tKzl387FwrZLvvB8mXxeLJbptv6mLNjQvLwgM+FsetXs
cs09jrz3QnSlJCVzks8Vrddp0u13Fyq9KZAUBEE1UKDxecRBCmE3t6x3glA+0YGPQTnTw6MO1Il1
MdtpayuFZ4e/tHrBoMO+hWmfXSMUr5p5j/M+v9eK9d7abkMsLUEJga/wTcvZ2teu02dIiOerEaU0
ZwhrDWunyP7QM0pmMFwu2s1j3BsoUn1Uqa6vga+7mEPiVp94NxifO/RsZoU4+jFDg8FOfbh2hcCZ
d0uAEVZfJoaZ8yj0oWznugHs5dZgkNsmjlt5Zsm5coMKnR1OZqsvrPw0vTyOTJkRrheHx5qVoHld
M4ddqTEqdgYrrZOQ3YVPdmyIi8pLt3xaKhaH17S6CO3UVIawN9SflumKLz9FJn16HCIqqeH/yUyx
v2ORbs2MWYLPwAceN4uwUz8Ep2JfW659gD6GPkrwfomjhIcMMQqU0aSVcUhpgrFMnBeTjT8z3643
q9+JsT9azxx1RFA+SZq74w8IP2QaeTjFLX+fa11dI0PfNx+k33k2dEBd0dCii4hGIkiWklFReoPd
v6pHg19vjvVJudWCdiMTE/tj2GekVI/J0kDKH6QBEXc2Q/1eWRatYpqnayPXvEbWXqnxGxovIa1a
+cJbxVWKB+A1Q2VWL5cS7A7t5EHwAJXh9QNzaIvSajXZu28OvR/+FNnQ6yCBKyPqwZdLyWrb+JME
8Pt6/y6X3B3IpY8QndlGZjOzblEZGeHoJyTRgrC7funNnAiRD5DGdmcYvLzjHeQGBXExomMoj16E
cKOhZr1LYG9DXOCz4/1UhRaQRqLhWCeYxWu8XjKKt213a3JRU+yBOYpeRbjVR3PO/ixqFCfws5rZ
Ii79UDdZ5XBFXviCs6zRBHlCrssbmf4bsjZ8x1otO4Yz8JBxLMnuGJ/pHGesJamKDKcayGn4m0RU
wLAblyB4vlyrfJG6FKNU3DNGpXl4zj57V4ExiU5NEyVthOdSp43Ulq8VziVMNbohLXExeEi3O5qj
FbQOYWrRUiQM+NN915vKaqvaF3/SA86PvdBmX8X4MqCeSy8rtPs75Uq2yMYLs37CQGI3pk5YXUEv
sD4olmaMyYIVNi+5H+Z0T/JYrRTANqnb1ICMujFOgGcuArbdvtDKyLCM4Bx3AMZga0Y442CqP2aj
mXV/dndrFYnu6KJkR8wEmp1OAQ6gx8un6NnbtVdMPxjMCE8RdvPLoqSY9SOmg9qQwKH9O2YMnQFr
sFM2hzD4J4J4WmSjrSUfJxTq/KB5td2v2kMpXXAnvjIkg3qwmfCfbHHegg6XViRHXEHTnyg7PyDj
SWKFiLPfZU4J2fjptIRzhqRLXfFL3OM+kc9+1uVmN1a5Ks1wwmO43qv/p+jlllGTgqQjsN9Npwck
UFzxUdFsj62hI2g5v9DEOQ9oJi6UhXY+f5WcVkEwNM/r/MNRiWHMdud839xcyuyLd8c6Bj31pUo2
X4aqEJmvTc0K0Y57HKE9rwicKcIV6/qSHEEex6vU5SEQ8SimY0VBxaBdacyKw+CbqdA2lvmIT2qz
AIDXpWC5DTXH7iTlQARBHmk9GUM0KriKP6o1F5PzDdMnM+03hWP5ToGGhnJaxC75G6yBoYtNDVzs
tCSF62L/w8LrbXYVp0Ta5hcVAdNSq/KC98sA7xqiFxMX8cV4TvDkRl33/DACMeJA2Wi6RRbduHU3
gOa4kTQO8kVaIqDmGVO8gWD3JDMOlC6q85eoRj4RxS9rLh7wT3pTTC+X37Tx4jj5TOYRqMLndmBb
IMAvaUE/tp0r2efjopbduyO6unxtdftD4rcBm1sGq0Oyed4TDXtm5R8rqeOuZ+exhrpkJ0iXmbBl
PMqc1sMZREDLr42IFUCkRn6PdoKOSCVXf3Vf0IpgijJYQ9iACNf62exZW0tM4zVDfohdyyM0JKMW
Eayg+zAjn26+/A3syHYq/uMUTsVuacX5YOGriVZ43F9r6ZOI0l743ettJiYJpZ0fO+7JxUyjIzF9
Dikvpnd7e6gxMjyzUab+GBapPbr3YXDtfTbOAAE3nKF+whOCWpGE8A7l7OjiaZuCiObaBQ8SB3z0
idktKmogAcyCle4uR7fk/VuSQ2gU2Yw9MtN6vu2t0W5jzEKUOm2H83EkUBbsxWGQ9RAcy+APJHmQ
sSM9+eI9LqW/XJXb9uXlZWaI5t1NXQ8Bz6U+z+NtHnxcImdtb11BO/PFQGOqVY0UzDZOe1CGdhbg
awMfckyjqeog8kbzxWGzuF1qK7LjxH3YQMPuMUVHHBoSMmQ5vPAw1z4J3qG0LXRXYvxUJRc/7xUS
s8S2G37Ggea5Q0eoLJWcobLMl2eHCufcHmSUu6Cn824ufrbbZqDWv0gdxuJAiMg0c2vV3CfafUN+
udWbCcmR0uIk3Mn+ArtyeJqdWtj1VNOFqzE5FwHyr+b+c2OfkD3nBBcL6BJRUea9NNCtsXcfwbA7
tzHX/kNWt9G7O/aATY8lxNg7ksHN7atMhCpEGsi0YlsybUTC4kz67dHVv8L5pkEM6xUNEOpf4iAh
sd2LRsRLdomk5fk3eEc5hGywzn5ernvjVQlIrnI45jBtIADUL3urODlZz/iHaFvYmTSMfUFixJjz
cUhh0c56UQ1IWq0jWUUf1kG5k2FUyYa5oJMHVvp8jx0jP2Lscw/MwBYmY26FazAsWizHC6QlmYbi
tPi7IgKnb+6XDL6nbawtEob69wZ8Z2iW6lDsye847Zq0SsJi2FGqS3MCxhg+hEeAmvGkgwnFRTR8
RZx6Snd0Y+Y0Ixuc4nte6HknuoKrdhCSjRnsakgyApT0MmG4zL9xiK3tTUIzRZ+RwcKfkPJBUIi2
Y7o7ymP905kUACT66vewlUTS2VjW+Q6OHHuboLg7RT1sdsFKdJXQDytcS9DW93bfZe5Qoq+pBZLq
2yvbdl10/fVy/+eQiT7NyRpBahROZuuaDnqbTXH2+F9iQAh7rBkYxRpjZmbrplkUmj2ouqLOUEsm
Uj5o0Xu+mbYudOrURoba1PlT3bwO6D1/XH/t+OYiRgvLJ2abFNTmldXApRsDtt4v9a4Q30H/V2JV
2d1D76uP9+xK8USUnxSSJPySmoNzidbjcgeR4gFTn90BZeLLscPBFZvlJ3sI/wV06oChgVCHJmtJ
f3DEC0hGm2ItS/krrJ0o5B9ObS0YI/lUFH3YXHC32PQP7LdwE7Ngjr4YR8A5Kn1JabmP1DHYCJUD
VuFbEslwFxAasmibE0Ucyxzr+WdSZZiIH/P5m8/AxbpH1P/iBTCcvrDqF+caTxQOiorJBwORpAZ7
mtAM4cBJgBWZ6IVkEXds9FawQ90Ok7k8qLZFPVi6rb0u/XUPJJuKvFO15yBY13tzjGQZY/1YT+ws
U5HV9qhYbjDoGUgq8GXXYa6gaqY8ILbzGjbQXR0m1xYU3LzWycl9/7Nce3tKndvdZ0zyvjHBHU+P
KsQnkZYrUYuWKmskBOqqJ6ZH0pPzxbNVNjf7b+qEbSK3435NVuNfKoq7FtIccSzfTDF8BXVlgTdO
fb7Bjclxj8n9XkwvvRFUQHC/B5GXbn8UyNPq+2vYFwqkhSEbitt7+dzHRIb73Po5ZTTpyltSydmB
EuFQsuHGDqmXaJwT/HmhuNokSrOy+2v96/VeKdgeHqXKmkniYQBLCaLUXkAGzICCM8sJhxxGSr9R
roNurg2v3tcJnC3mBNK5a/iTCNR1lovjTIr0JuYJMaewbngpe7KW18AwIwua5eWWVEDAf0WZiwhH
JP0MLMylZvuTyZbq6LuuWkjU1r8p4wMshS1EcRy1b0DOskLghKI2yZv2+fck60DHUC5WUbZM6ILo
KB0hkVIamPONiBl+9Z6nqw+0sR2K7GZdy/VBY68DXfNt4PsRKTClBuZl8kvh05Cn9JywIYdtQCih
y00zcQ+MFhqqEcEzTPyyka6/ih9n5xY1JWWryO23Y8iNzyp3r8M5DdZ7tDPgTJ8eeLXKahVO7rL1
aSlnY00LqAlawRJ/GYqVj0pkffcKwyB+HSpdXK7P1au4v4s236UvVcreXNibZcD3uwMCoemKyxpj
9AlV624+UlQVQ8jYNCdSYW6B6u/QuU6JeSTb50pFKAov+9+E5PZYDj5RblHfB4z3Pcat185BWpig
m72PF/aObKFRQ2WvsMvl9ogl0b/blaqxvO24fBJrob/tCJoLjqG1ItNFqyf+gsmbyV4X8OYcLvE+
xuOkG0ZHgnjKv+iOn6JkRYQd5oRsdF6/LPanHF1ocouiJVXJlocTeKYeU+NOtn9+TEnar+2lkzHO
EGSW/l9VuzvOds0bDZLneAXiLzZ3PJkTVs4ZVw/ArJiwYVj7sA2tzXoT4ggy2YM9NkETI2O+RTGW
eZHylQPN2h4Oxa1091J96+mBdN/ODnCcTTjkI4K7AwWkWUeAo6oPVMc9Lt5pGLQz0ArVcqXBzP8Y
3StOifV7yKGZ3ewguBEIv+M++cC1yw3umruwoYlTV5J9QL7BQNyWCRAjWs0QUEhGM2JezE5E07uI
obVBLU7DbVhfzZHycbJ2+Z6OfPvMxRwazObxt2JmbZVa+ZJ7VhCPNGXYXLy+3i2d0wqf+DzCbdmg
ezBTJ5jpK8lZ+KFwtJC71Z1TL1ksV+qifBPgE9BbTYzc5Ap53MIth9txx01q7o2w5DjjReelsF57
LA8O7YpELQTTnH9mmLO6UmgWhuz5o6JKNZIIxiH/zbb0LxkLYJbhQPbBNlpHjST1ymxTrC2PoW8n
Q2pssuET2UQW6PFWzm2mPB2CA9sYkJWFxMzBEXMCneZSLcI0Mpng3C9Dho13QmmKkEHX6FJZc+xG
z1+J+zSubBNf1zeFoPeYKmvwnYrqLqgJ55/fZlA0Fk4Y01oWvjZyD5ye4c/RqtE7xDUeviGdv+fB
PCvd/9mPnhfvP2YhndlLGvJKBzldkkEU0I+paJAC4yjt/b4KSdp9MXA3lAmqb/ZE5bNlnXX5iZCD
NrB4DieC/duAHJ6DLKarKtGXFd2ftEB8qKTt7DOockbCbgJ0Ok8KAdL74zOGx4qeSC9pxgoN8aT5
rp82SIJ0u6HulSrokYbPua2N+kLS3NfB3vuSrwy2p3/BfVGo8w4SKCl8xeac0qPj5Fn0iZ9SWaCu
/7Rc9smUwnK2FSvdSukBkQH4efsf99x/Sf69mLf6ErC+2OezfVAyQRqIECDFFrhrc4mMG9BTXfL1
ncvJkSCVFJ5IYsNEuGspWSRe5bs804W6a6KCm4IIAd5Eb5kYJo1v0N0DaPD8tuEOtKfIxc6IqEBl
4cISmcNJNP5YU9+82sKLuiZwwB+gg/1WOPyyJhXso0gxM+61f2rNQclIkyhdtp9RDEMNJiop7vcS
MzDXYak/Fs3kUB7fS4evqd3DbsRkNLujWhpXPi5kLpBEIWHRGQ4ev2DxNPZZaM6WwbOLJECWCvg3
ydCWhQ2nBrkvBZoPCqDFDRZvEnw2Ns7UthIGJiLcf11T2of1krnyKHMrhaH7xEt9/sO0mnDDu0mM
WFbl6FPZt2QeezCMpSJ5DVm5tDL6ldsix4sP0SVpTJBCCB2o5mSzQm2vqsNQM1cXYT59y2roylSS
vh26VRQ4Gd5v+TpD8Qq0DVoE9oEEh2lNWKzbIyc3Q0GTPITy73c3M5uU5ProU6Q3HfYi9+fMnfyd
GbhW3w37rDBzbTL04LVkTvw39a635BAfbl2zaKv+qMtIO9nsrPOWnZrmDRah2izzbl8ONpGlyejw
coLcqkMS4iaID7hb4RCGCbF3ZMR7TCDHu5Gx6wsk9YtPLMqQsv6Gn0UnN7BoEH6nCCsQAhj/inq+
m+3a5SZN416uTicrbpTEv5nbleWWmSQ97lO3HVQNJfaexjmLP+jxFz74pzM1W8UqoKa6SzC1s5QR
PTslm89rI8kGOlAykNThs7Rkd30+RyIn1naM6jeKelleRFI4ngMwi4ohv9bqUk+nJZ4DJblNKu9U
TkQGBkNXC7NbFQiM8NbhLkf2GdTHSE4QBvUrAReTK+1N9a8r60yTyuwQ1Do1JcRLRJEKsM2jL90k
wpKypKz9yeNgDFRfrQVwZzvEN4FKfbIwdVNU49gE7TEZYDBZZPGu2aVtgW8B46uldd/Go4McYQO2
K81S83flxmeso3Ic9e1kx+tIf2L5ZrnumPXLl4bR4CzKRQtqgnaHm32dZH9t3Pqp3we39Srz30l8
LFI7DSyiCBp7ILULFAFiwfPEJpoXtVo6Ctq82HgSuQpiPs20RpRmyV+ey+1ocL1BzYXA/h+Yws3/
HnheJ42lQDS7bQnJoC4yPol8Hon6Y0gUN/ANH84jPYdQ08fIwLyzlCiSbHjRCl5v5dgB5v8pxF2z
Lxw0aXxPMCN9vHBmvX+XPsYr4GaSLbreKCZT5Sx5cTMaIgfh7/T+wh2+u8rJP7QfnbVfm/XAvvGX
MboW4Xy7ckN2696CgIRPnC54I9cbEMSCqB4LM8UH7Q3iJbib0AhUYsMNEdO7/w9jED2Y0aHLa4E4
zCAAvJJroaO02A2gSVO5bhOnZeaoHfNnys2pcJHzoZTeQi5fujJVImeIfw1qvim9gVc5Pw0iswUf
Z4rW60l1tzxfSToEEGyc7U9NkPkZjh5sgHaOxivdV1vQh6H2jt6a8bQXi1p21neNLBf4kIDo7OQp
Q1o0a62Rn7QyocazWaGdl5sRzZNPimfb8y2ujDAfSsOzI5XPpFZYU3CwVOf6I75IWKUtASCqGMIw
X6hMt0Gx3S0kO4g0hRPIluxpRCNq6eUKt0o0BnmTDd8k/adKvOSGRILuC95Jzo5KgbjMxovpfsL1
G5wlwAeCMcUwk34o4L0brP9UPufLt4sQbjShvF9uKsz/FUwigqWJsK6LwMW+R+uSLNw/7CP+jofs
Or2GKYemJRzivDUcsLKECh5djq3WpslAXO6Fx/3k2/d4vhX/7ciVM4A9RCaJoLuQ40FXWX9rZ6Ry
eR61X+fUtvTGjc4AiBKkTIWY/zkZYeqELGmGo1S1T8PthaS5Nrw3yVQrOZNoqXgBxtmsRbjXwRHT
1eQTVIS4OC/qEsorves1qxzPtnjoLKN0QqgJjMjpXQXOfGWEoozlgYfzzYMw7nle4p9fj80G/yjp
qZnfpcErHjOzuztCBZ3kCWV2IMtPKFXnbvJXuCEJiIdsRPqxP28eCPXpQPUqxbsvzpt05VmBXh0w
bgqp+QHE5APAMRI0Q/HraKwneOQxEFtszs5zYbynz2gc5Pg810X68wp8HBHx5FQUjdJFz919U3Ki
N9IjHwc+9+Nc8wRwlvC8C6ootq/nk95K+2oEqWumuwepYSWNRuh3UdFlMhV1kL2WTo6RZr1xDTUA
7gaO3gLweRFQh66ifwhAx83GE45LnAy65ll0OBgEpiKQa2A8NxHbHIoASs4d+unS9+QRwosbZWHG
Z3TmvZdGCLzxfwa4zxNCGQJ+BZJ3v/YpuPbuiwx3a/H8RPlUZEyL9qTmpLc872aNWKYVexlsx/5O
fQiZ+PTjTSQV0cci7433TSOCL01t8A2sBaAjCepxkfruJi+chVve76B4lq+ipacB9sGInxS4CDkc
lGyJ01EmtqCK2eyhnDoQgkhf5yqu7nCw/F42s5lzPDxUmVVfD0WTorIGmYOkGl2iPUcjm5cU8Fk8
QXwlvkRLsYQ2XC79USyoHmg0Jvdlq0w6fBLM/llc3TGC7Tpv3RMinr7ip31pHLEYPyTXV1iQLT7P
8jii3WkmbZmf/tTKawtyZvntO3WzO+qrxktBUt+78iMMkXVo+XSM+DNR9khATuOBtCAfDEr0E5ck
Wu2DcO3I7NblilPGweB+aOrr3srhDugwdaUa3ps61WF6DP1lQpE8d1l5nngnL/eHUwNFeVQY0KQK
m9LQE0Ji+JgsGca0mAkWkg/OZYuhNqcTa/kpUGuB0ASylqo7T49/WR/N0MA370dOYQQMDAjcykdN
nxHtos1XRDLnDi2MLdCI/MCjJqVmc+CIyuL88sAP/zq7cbe511If5vT0S0s0iSDYUZy6dCMR26sN
IvkODf+jAWSED58xrrqeLNMKTj40eMMkUBHg6VTNJcqQ/Y10rfuQnp4SM4lUtmCvW/GrTulUioVm
bZyWTzvIQuAclzl70o7vDUE1MGMbsrBe1uNWp95FwATVFFgY7Lu+2NLP6HTH57grIaWaAICCkb18
6Knp4nEwb/fT6yZb6XvU4sHOPKMQUEaWI1poeCH5ecEfJDRxJOjLbWBGQIGRD9o818SzM7C3s4S8
j7gvZiIBU62MnjQBiY2sZ+LXfzMZJTtYflw6E5j8okklllhJ5Az18v8SCEW8UgetwPPDAhBjnGqz
bFEbOJF7ZOEXp3hEXxMgh1k3GvcW/VZX547zucaT3kMhJyXNs0rP9zm37wEdx3UUZcRLFkgmMkxp
0lLJvgYwHx2uTKB3vO3cFdY02yegmMSrRh09UJuatH8PcjxOCmMGVFUR/axk8blSuWeUC3FqBDEZ
rxTo+GSG0EFO6K0J+jc3S26XuhN7aIfUiaFe3B37FbQSOpZ62/uLHw7v++9mw2CX/3JgR+vQPqVT
RWsZctwVyeaeIqbyFy1dzbN/IIBgbsl46+UO22bMwqBz7H93Opwcd6OwiNDTnEuk9bHHqSkru2mQ
ln2V1DY4vhKKq7isqAWT+kh/AdwABHEkXSJXnZd+S4MCIpcLz4htz3BKq4MWnvaQJDdV6P4S5OZa
PKT3S6KPnljyoKvSC7hm4gVPsCclLxfvfol4u3xMWmUohMjtudYQvC/hC+jWmNocIboaWxVKqG9i
S4+AvHz0JNNGeRFmgD+8aeWp1IK3p08YTWYoTvyH9MSI5TqjBKw7fvR1yERXxRlpAcNytdgqU9Mt
uhxy3YTcAzMB+daAfbD8uovI9i6rP+ELGTrjrqZUZSB0zCHH9XyNUGmMLXTeiQyI8vDEogCUBSjt
de4Kn2No9cDd+lttyHL8tDZ4/UrjZTgFOuz20n+vmQHIBeyfO18mVnBXnWIfME7C+VDO+07Qn389
w/AbWBe3Skk9VI1vpgcDfSXGny25Gecg8ZWuLaiFuXtd6gGaxRTGhm+wpUEGjjjcZUmevcdu7lPi
DPBjWthlnJWfO+TWNfdQs7wr+/h2KV6jcZgzwOAumRlv7G0cX40Cr9akLR/Su+4DC+qLpp7anSpJ
XLjnB0845y1cHic6zlasthMM6LLGhB8O/Bpe0mDD6gpFODImE+wImmuzXZRxt1KgIxuV/nilrycc
W9Sl6i953BfKvagMT3YtTw0wPfegOMJvvv48aQuIZJQ5glwHIZPmqmT75RkbMR9v0GbC16J8haLX
aAbGq5B/i30rLMPv9LmxxVOxOgMQr1Z5BirHwN03s44K14CPrOYeS3hi3EoLrM9BxXJ4/eMxTcH+
4yLSc+lgblIVQx+SBCkG023/RFDUjwkHRUBkCdICz+RiLe6OpX6zdaZuTtROQY8CIRc+WmAq5HWk
zYgsIolkuBo1Ksx9/IsCTBivIf+KTM4aSEzrNoQqAdonmOUCNASoFh5PUeFO2E1AKEpZfA+q1YcD
K1cp8x5V8oONy/+yFsbab6FhwL1sfL8yotArQoygzEyQ414IK94IEgQj0Ro2EHDGp53n7hLHVILb
JbqDeGe6jNJFoA3XKWrRpmfSduW8h4s5bqoRclJs22+esS7BykGgOJ+0M9hPcaYXa0ntgPzaXjCV
PAG6myswMiRDdc9URJpwsfcnAEmy40QW5t/idvTcQ6VWqjId0cULj/B7dlfwJfqa0O5d9Qg96T0w
2NesEztCMBQY3IwfLq/uiTW+UEkH4FS4+fo7mz2Qk9HmGYxDi4SYba+Is+tijTLPbncm3pEFg2i+
bnh4hC4wfDigv7FjLoEabeWECg4ezbRCP6WmZVK91AsZnhFtgnPArqDdXNSD5SBr3Bo7dU7TifhO
uDl87FXNjdfT9IbNQAdOVMNalXWU/5FgmGRdT8cErFBQtNpRIRp9djlWMAkJ6ZprOY9BvRvQHUhD
VTVXvLjU/9OVTTpXmcEQSP7QjYqut10vYpTzN8MaO74du9pdJxTZenZGPektFAiTuWgXmg2UYbC6
MvhOODbNaVztqAH6GgKz3h+BqGNunHtIS/j8OeQwsfXio6QDKXV2RnGOmFgFDesIi+y2cHXfZD+n
eIq60Dljr2VaBTJ8wKEiKEkRZvVIL4d+fuJRUPVvt8UNR0W3oQMw+wBlczTbLNGCETKCLel/J8OF
BGNMhIArYaSo1uvMz4hDhGyqgVk5lqGBwSlJRWJkkhV6j29ZeKTSR4UmFjvxLeIq+Rkjs6IypBog
V1lHDFR/C5VMII/ep1UpCcllJRiZEAMvfjW8rgNtm1QegqQcRPrit3PgaHR72pt3lcY3g3oeykZw
jw5CmTdXuf93MnjduUwccGxKJXCtprEqHe3UlO8oM+1dJatUpuNrMFSzmSWdJ/Bdc4TqDmq3lOGV
G2wH3VWssEUmgwjr3xpt2ECcXacf9Yi2cbpQtEdu1Fm5nfpnfwYUtlFhDxcg/C0khtAqzR5jVCQX
4ESg5CibbO7m45ibmZUpZHEvTrl2RB5lSKuLABUdCBEE6y8+/PBP0wZApGkZZDMmNjzSvTANmGZi
2Xwimxi8gD7SN1vp/W/zXKokSf5SGaXYplh+ha45DUGw7G2avFAq+MUWP3PN0JvhhXWm3bdo5F/c
rptahxR3gI3VakuoFnnO9j56GYma5PfT/y0BcilAoNnQIuLL0idbNE+U30KA00VrHLx7xCr9iY/6
yXE5nol5rN2OdmppYogJ/cKsen9amgmHwLivn75A3CqQCV+/ssK5vHPj4y7rvY9ekhfhbRLEm9ZO
sDq3dxVGfib+zIsnnOrjeWtyEe1yTk/k8IFpzq7RNqCxHTUXUjjCrlrIKGIZtRo3CfA0JgjWjqZy
QAHGhxcpWo9jjStVWXmGCUOGv+RL+4ov4YO3BC8J9Q2b19wEPqDbNf2I3KXdBj3I/vyg2k+3wpNe
qzklvewOjYHaZiFkmeAdDjohryeSnW2FBK0BNElSZEVl9AsXeiGYQdYw1BYml3Y5FJyLzM7/uLCV
y29/pHkjgvcvs4tXTH6XnNymmh+wydQ8so8U5+4DqQV8WGcMkYNCxeG5k77VIidMQOr78KoIBZJb
rBmu5e67YjDNHvnE0V50w4T3pCF9F22pULokEgItUpJzrSv8knkfvwD7Ji/f0Y0E6o4ZX1DSlvbm
WLWc1oPZXQ5qhcCw9guhql6Erfu5oH4DWw3X1fycBLfbaJEGb5hnLyKwlxnENulSIOBRW4FbLUWo
bba/F7TtIpTjWVg+n8u2N0lY0OTGBTtaeeOToD0g3j4HAN6FIAZ2MxE7lxBUGgGzvsA3mRZ2iAnx
i+jdcsvE5VGEU5g7RDUoZ8GshMZttnyTKQir4ZpC4OUT2fwRtHBgkfJWhWSYPfIVOcY4j6PItCG1
gIHWBeKFT1O73GhKoIAQjAslpr9fKM8uHqTCH13TgLK+sZ+IoQf/175yFDNqKhpdnxULOKUPnTgH
VS7MdTWrc6137Yg8dVWgyEPP7j6LQWmsqO1dC5dg335bpOGKpkNQ9BDDapdUZls8K4p6Uhs5qQS0
NVUr4EQOHlcvpcgCMdFkNBowHR0UlsfpnSQYtViFjc5/8gBvV0B0J2pR3m6BqFo48o1l+mxerN3D
M78i4ZDtm+zEAk65wSNMZjl5iPP1SPLJl196COl2JOQdwru8oHFxiupre/83O0LZ7jThsrRJFcyA
V8HMY5tzfg0jscK/QiBKT5mgnEeebSvdJZcBuA6CDmPbhRBIkfEj78l1lMiuo+OHO1wjJ31uduvu
iGj+AvAe4C3mUEUYRSZX6FB2nhVMu7dhgTDmkuWZXq6Pt3r62J9zG2yFs7Ixfy/lVUeBXAngme9V
ZAcAR9IjEhuzAR4WZryMsHltG6gfoLFOmHNpICEdwbaaqqqy+qljYXmA44lfCepXJxZAHXGD6ItI
U5bBEZ+3WU6d6S1O3t9WQ7ZqrCS/1b9Z3fIqTlkTDPkPpL29frRee3ME0GObbYOARJ6bEgQpqr+i
+veD6djgfuq3SHfh4jID2DDyYnomJCUv4NrrNG50yC3cuJTLkFZVGpUHnnlM/0R/yX/An5lVKS+3
RXNzZ6wVMffSThkR9UqAtYJ8JWKPAa440+hnOFlYCeETwD2cub1QsvYBsJZRC3rsCinGFY5iWjp1
tMNeHayOZuezyqD7sDlHC5uCK+krsWPrdSdohTr/AjwmGv3YyMO5TJ6i+VjWTS/eFWuTihtHuna7
ENDUpet/qD/DQ/XdOiuSxuLiugAz3k6rPZP2BU8rWU/snw7k3O2Z0PvS4SHK4mIMfJc+BRL8f7kO
fD6nJrqXj75YMmHGKtNsPmmKiheEr3rnatiuEOLZFJlq7wkXCkJ9gN0pZ5Q8JQHSxDDBH3xzIaZx
BPc71j7xdGbBQgWUdgECOQG35dbhUTjFspprKDMzPqeYT0CQhMWPqnq6wezudJyWDgses0MtGT4s
KSYGGPSPQSLcsBYWrbPBL7BnHIYmpFH6P/kdT8HrBopEsZZNbmUeiNVtySo+ZeTdbZdZxJTCa0Cj
ZzWKoWeiTtOWQGLgd6GrMXeksndJ5dmtQcSBycvuZnWPC470jMvDF2qJnNrdS6+0YYo7P4x+PRx9
bDuVMtZl42btUNMMu1EdMAtzYM6OQT1WKdtbAyO2kDOTqV7vvHocPRqAcOJ9PWOx8KDbwgZG7YsT
gg9534hhsExsA3HES6XWxUAzKJyhFMGPfT6qBOCL/ieCBl46fKAjLD8hB+2ZdxykHqvmWJDUoQA0
ITtXpUm3YL0cYFBjdGYAck2+HfFpLDnobR/d3ecgFWltOJ/qr31W9MMup5ePzsVnor9qCgKSlc62
2BzsRVRoT/8exc42omgq0Y4TkRfCE9E1RmmEMk6Cz8FcgCfCBKceQyJfd7A6KJft+nzybbPPh7L4
NdtIoM5ODSiWaTAa5Hc5gRZ++Fr6A5A9KIFVapHa2flcfcLvZXh3T8+oYHyAwl/ifvyu7rpyr3L3
ELSkJZzX8/KTuSgEj1f6KTepOtyycy7i5jlF88JmqFwwWI/QDUZ8Ok0GvGXfn0iV6qrHOlaxzMqG
lzasTocKxqcLqGNod6d7ARn5W9QsbP4ZWXwFcpj3h27mTGHw3fQ92NM9ivDTZ9DHQvL0DPCUMuum
BMpWCOhrxeD8ERHAmgVZLszb082fSFVQREVQfouJKKYni6+DX07SaR36YxuBR9CNZyPMRSl+ypwl
FoWnBKdf3qGbp5j9tKX7mDS4c2ExVa3rAa/ZokCpwOrXWcxbBjawKeQ3iO77tBuvlqUrDRIvBFQE
WbqkjbWBI2fzvKQkTQyK4vdj8eATaSRR6UnqsFSJjwwDcDJsEATEuRSU1yMfHkSU1uJZyqkXvpCd
kyPK38iRZMWaIhgeAvGeg3jZl0PrYIxKDn7cPu0cNqmAxRGBotUfn99Dv2pSp3vVXOUcHP+F1ECx
n6jfIijmi2uv48xJX0nh/fhVgmviCS7FdyeOvy0Mn+I8bNOjIc8Y4zLci5PI7k/j7PPgrtNyiIos
dW7YHiXMEtOyFHLLNP06rBRvvRzoFxIZPtJV5qKcujRUJEaKsLzNaHgd9B9uf5Q9SJABmusdgv/o
KnyqnqaeDH4XRTcKb0ZbaYkMOIcxGO4o7gTmQtCm7JIEXJkseg/DWAP/Tt+9olCl71COaJavuqNI
bXxCVrf4Awei9xKEQy/YymyrAi4uUVd6WG8YpyryoIit+wR0OM+UBK5RY4IhhTfKO25uLhtNlb8r
lTymjYmK6Vd+QAbg5z4GnnB4rus/1bW9q1RqvaxdYergoLbI2/gbsmKLrFrRYvV+l03KYX59lVhZ
con9HYhG06m7cDfOw7z6j42TnS/Enb3mpF6IHSEIS8Hdnn5w6kiLx8M3H0lgNOeNIpuqJDaI1Eht
hrHWYgvm3hrHvgMysZwCSykNHpKBud67RPueA6dfhI1K6n9Y8MZfJiImNlJXWAp4uWd0ni2ad5mq
SU6VZpTwPp3ZDGxpyXO+1b3PjvUqwSVaFk9L8wIdoVCUqcmXpKq8v0KQoFeyuTOOwzrEv+NaapNS
rwx4DcLgebB3J8forOHRBQgEdUKiYPKogxcwydNKRERLELsXOE4TDxOp5wJFdNTfATpilkBtdV2K
i+J1PvAXIPHqLxc2aqqx/jeow2vBR8j/udxoLBR1d4Zelkpw8dSLI5J++0OgfkqyG+RlBuKWkE5c
0OyhyaaqN6Nt4QDr566Q9/4z0aqMBBRrknut4KGQ7WqtPJAPKpezw/jVcinNSDpm4EVLEvs3bTa9
aqFhsGmQyedSgBHfF0EuKVzbuG3J7gFuvqlnWSInoH1vql5+kPlfaIhc2L26kgIjSnAXSDq5Tr5P
QJyu9C/+9GzpAxcXC1hzl7yqBK6axH7JfjluTgMwhXwM6OKpUp8HJitz+OTk+9beIJz26iSFJ8DQ
B4KAn8j/VGbm1QTpBAdyo5KsTGPo1x80CXxW4V1tuEmr6U80yCe8aQGGTMXx0wZ6r6SIXSs3hUCC
T/HmVF+JKw7e6/SYgd/rTPh/vWFewfz2Lvg/UGnPhyIBzyE7lgG89LGErmd1+ASgXQvW0RJRyJ3y
7D/TgaoTV+YzJHNnK6EvXxzOdLI/zucJ7tyYvPhuoiph/6GR3Vpdsaw4sACmsRl+Eqak+XdA7df3
3aa4ysZWJ394d2zUfwBL7Pa4tQxoMkfX8741hkqmEaxTRKuvA7iWPzMMlv3UtkWDWT7GiZLXHxvA
09R2dfFU1+0DQCDgUseWD+/t6jwWmxOoyCHrFT6J1z3fXEHVzzSA5yTzv6D6uZYY+uh6mbHEy0zr
iCPwrIPBnx15Ht0eT4ABiSFCnSIS1e4H7b34LRYvQ3VeDtw/8HctRueNTMI5+nKJF12KRUbcIm3K
lRVue/AkNBT5KQLG4PwpT3Ou9CBKr9D9FMTldFlQTsD0UuEWVCjBFmxNZbzUnDkK+pkOK0ccPpov
0NOBO2pBEbH1GMqjBTuh3Gn6voVTa/hYay88cyc8mEsmLxEt2BISS3Ry3kW3sblH5asCkgQms/fS
e/+uDxE73OCsUMP3WtsBH2QQZP4aRX0KFwF9s0dwr0wEeqdLnXsLaRHy8ERoPGfedErbU22qUwOu
trHbeQv0pjoYSTyqIDYh7/csg8IMFYBYys5ll2ZF1/QWPUXsNG2r6sVEaPDr/WibErjBiPJ/PzH7
pJmn+apZKtMhoLQTMXbN6jWjXuXadmOn1mVTlD0tR4Oaom5lFTEVvfZcj7ANZHhWeHYXSdo9Z7ub
DFbEE/t2U5j433XgP1fBODToTBC28X1Ezf5N/O7pzrBfDtgJTQaBhSJLLa0xVZU86Rv/oB5VOk4I
E50E38oiNBRYhD38OIKRxg2M0kcCilob338S/hAlz1kKm0sKE9AkpQs6PROqzGMDXdlFVPGwJy99
/uwThy0Ybkr24HCdh7dLwVo9pG9bP4VVnms5ttelM9kWppcOO+mIX2/9hzq2IIaTdfvXGmFdNgd9
m3uspDKibooWwVvwvOgImXXA9y+XtawgkWAoLvvaI3dpqAe0xNKfkp+RjpAMtOcaXqmIJxE84OXP
aYh/iGXHqWRpvTZmjXtBDgr31RE6f/67knZUebEYvelmycwOKjUBz10Va1emIHVUWaVQL5G90kSy
7NBH+gS6l3eZLzjl2HHmdUCzOJ6DzRoC5WecfZOhJZOm0AUXQsjL9N7vWUpj+Fn81nnl6A1C+5o0
U8iluvr2hdq8xZ0xipAmekUtww0ni3ZFf6nD73FrCAYXCJLcG3QTgfsSi3nj6TG+VCCp0aLFDf2+
U7qp21McZNBT6wR2D5WNcYTuY0n8YKPd8+npFmHksh5kGKp3D01V5JuKEa1qefDa8WELj/dPnx4G
deJZGFmvWARXy7nmGbHKZ1ZP7wU+IVqZ001V5bU6m05FCHxxdngW2oNLizICsCZ959oSn8Wy828Q
Dcd5tX2dY5CeujQlmyW4iPz8U5ebRaH/Xwzs4Gg3HgvZzd1VXUZBe5mN6soRiBCpLlQEjIg+IjgI
wS1rz1hA7E2FYcVVSoFtkwgInjlt59JhTGQdApdTGHxsG3f0KdWfVkR07LrcJjuDuUq90TCGwvMi
E0px68coYRCfjBxnz67qJypmaWthfWMQxsp6MA6KX5FRECKMgdAcKXxZtQy6LKqzWVXaQf5u9Cck
7kZCe2LltANGyn8agtr35GGQmVXbFRJ/n4UGrS43sjrd7rSFA47kbnHKrr7QbqsnJqc88qivC1aS
AgJCjnyXBtuwtGMn3YekFohc7J7fCM1FPz+1i5D686H1fzgL58xtSltv10K6OOF4YYp8Rb3aznqC
1Osw32cVWMPfQFGHBqqyDrwgNlFRLY48SToJfphKpKyOGMsoFTupusnJFUO9dpAYxBR0w2Wjpbhi
L8uv/dUVPKPmsdDfajW56gy/5eWbHQ7CPbJ2m7RzTgmdAePsj/ullWCESPia1+j4H37g7Xr58TJd
qNldbmGjXTsdskC5YjKPfLsmwyosp0VxnENcU7M7jViBZ/LkOBbmkRSXeznrqdJfHIknL/DmeLBN
DoEH5ADR1duISj/0/bStznYs5nrHli7zMo4N0bF7U9YazUzS8x0UFlXlF/CuR2GYEnjm5MMA1gjj
kAD1Ld11f35D1snv/wdg/4gVUaN+VJ591pKZEYCHINWLn8PDZbmPR5UHD51ulrMGfPw1fyZrciDq
/jgcPL5v9pt4ibBu7QlKTVxpL2gYyfBlph0rwyALr2RfCnPlgOsgcTPXf5JXtimKOMDeNS16gUAn
dVSyvupF8W5AYSfDjJJY22X3EUliWnD6alkGGb1rgJ/m2m3JahMw3CrE5wtD35/XhEe2jtqsWonQ
+KcKeG9987m/C70gRJpcvexpLAjgFoYGA2zXz7l+MVIL6mb8AWkdD3QzSaMc1FCxmLC8zieqZCoL
n40dp553/n7EsMbHakgz/1Bo160taQwVIDnEKcCWEj1F7SsZ6kD9G0O0MBrziqhU4UvugVHi9OLn
h2WIhH0CmCLYlVXazw9iUA/gQpoF+jpv0A3H5nAfQWhsq6SZjM69UjQ111GGyq8O1xCj1BpSY2Ti
G7/KY1mCv/x+WBsqs78kp/ASPQ7TN0xWZlCDI6ySbN6FdeIWMDW3VSFkP5PDszkR4wuP1TagW2m0
3uyKBU/JzG0fUKzmEMjxQxmfdL9rolZxP000lNJq/oH1GH4cUA1sV3Xi8CaS267Czcwb8ML6JpSI
vDzjnAnDA7CJTIv6xdr9uOlu1a/KRVNRjwUhAA9KS67pGzekvZK+O54iGikxMHHMILBdNlKF9lFw
KE5gOsv8V0BdaNVj18BvJN577YwXVF6OQxPHQKxI5L//06pnjS/ZWCPmHIFStObTKv2v7sO4meLH
thKHS+1Oi15pLmPrxSyn8KKQZfSEpmp8WZkDknQf06ZlhR8JWnATlQACcaHMK/mtHyIxAk1AEHOW
MIKr1K3/g9RERDpUAs8x8pZnqHNhcFqSFlQ2AoKer12sb/QKJd+cjzL+NXTwqtiv8sgMgT50y2Ih
5dOJ6h7KuIdgo5np+bkapzTau9qwYLvL+EsPbt/WZA6eJ8WwaIsIDCUO4NwoNwZYwb3HGoVX5XfN
DyPzNpVvHWLMYzUj8U4zJJmgSiRwxg/jM+JTLK6c6D1HGzAJVGTbmKCb72ikszXXinAxWAv67j5X
UMtaotazZsbbzKJkWadVFgaqllvCbkKdQY/Ct4p7FtJ4IFFwcOGJyowigY01XaQ62bV/tJDnpx8Z
awlM/viS5uo1VVa5rmB+su7t6E5C/RmzYMpsoGbiMq5LNvge7770fxXk6WmQXsNd2elyR+nGs5j+
nFcVXceEpDPNJVtGVtXSnOzSwgZQYzGETjJp6WuLN4mleGsfRH633vP0g5CYbI9+qfidNJ61km+0
BzvH5WtYfQ8Wg+OX70sMQBUGbCgOCDVezWYU4wP7Z2UOSJi7pLYSQQo7wgXt9c7iYjWJRVWfbVtj
alVPgKA+NafGR3iNPrkCwHJEAAKWIww3tlr/8zrVcZOQhFqgp0Bp3btqSi9dG/HI22wb+twlWRgV
cYHbfYfouVdcFE1Ho1qz/xsyoNQSqRXcJmNJcLcosN5DkC0HshoSe4DNQki9TMBJVgZ8Q1TCnzM3
Jdx2XjFbbx18uTbFBoxoqFerhzDRJcNbI8UO86E1IYjaoDhJ7PkoAIisz/38Jc9MIk2qaIdiloiw
W00WQOWDxXBXVrY4/tJsLF5g3GAeDzliGh0xyPo2SjTm//C4Fx3ORHa+1Lz9RBlKVqZXxDgHUB+P
YxSA04XbXqiiWFJaLEuhj0ts3lbh4QDK3HK7D28eB7hfu+23yFU9snHNWdTvGLkXQkrdOz0ThuLY
pvytrNiqbNsoMX4Z+aySZPOpZjcT6Z5WZ85f11KXuSRZcz47nThO4l2RWkvczvMmJDGZUAXnYrnb
monU0VDpCGnqavRrAZJNQaHCbyRBRQb0F8wPkYwofvC1/SualGCFP+RkaqKogxDjYuAf9ZLHaXri
6Bz2FPNJQXaWnuqnQfRd4cDalyhxcUGWU5sUnZe/z4AK1bu0rvlarns19L0nCFTChFfTdVRMP5Vl
8AxGawx9fB56Wmj4tQljCLQ5kT3CMVP19G2K9T0JQLtK5B+u1LDAgxopTj0QBbB8GScLYy4+96oh
+fjXpqGr3nwqZBh9hDJ71gcaxsgUXMi120hEDF4fd5tzw3JLX59EGQeJMZZVzOvjiam5RqRaQtIw
+FSgNlJatAxaWfdpCT/fAKf4Le/UZarCHGF93RUxhIP81RhMVBd3bxk/+b/ElwVot05JvBd+Ehak
k84MOj/eJaCPP+AWsngPpSJGQmbxBUqOa9wytZyOp6TJKeSbFoxucHx82d4VdtVCHLSqMHSx3wpT
XgTC2gWCKrRy1MgGxVJUwq7n8RjK6/AQuI9l+T6DPA+awz0jb8N0QEQayyyINj2MHWTa4oSDDs0O
CfeAoQoaAl328zeLOWMUimi/5agOdExgsZBdXDsU5BMk16qYJPtx5aPu+f4eug2djI30/dkr+yZR
81IGuPNiFagdgYSxKCuZ1gmX8tikujI4nyoafbruXcSlQjSvTTEzZssPKNy1hZsXs3BdKbmijAZe
2sFQibjw795589E0Zf9vJwRFf+DA2tciLte6wLoMRGVvFxmO3vXTSu6GhN1j5M4H+EamcBKvDHYl
bMPWWIMlXJ47A814yCExjxqfZiXnif59x6BXYCu87zsKfjymU7ZtrkZaySau+qja4OEyMxg2kqdn
OZ450tLlOovts7a01d4cP8sG/dnwsB9XLxPpA/4QFRvLUnIS7OxSR3bKjG/01fj9taxZeZycGMip
yvp6iNpZa7tbRQ85MQHep7h5By61w/+DtVbxAX9RN1axF/7PQKDKIBHGgO7s9hhoNkB9+659ED5N
jw288gWTSamwr+FkwpezZ/Wec8jLEhpr4h80lYmLGdf+Wjz145RREMZYttrb+6gGF86EsR8ua9Fq
WNgY5M//OhfTMHPU1o5MpJysiGVx3oX6tD0bP5Bxrzr1IuYG6wfJHZpXWwrbr6Sy+stPI+D0E+YL
Ng6RrKa/dUmWqfAH1F5b5i/vmLM9S+9BZlR9ak9OAPhEJqWGF9Oz+rQs05MHE5sy69bjDYEmyTYz
xHadtn9jInQENZZuqKKB4D6ngpN3n2UDC19Ks/EO9cBT+znt5ZVDF4oRxICtbIyEUzbNq/4Wxid4
/cT7ztKmUHVklpQ+Rz75ylHLWM5voOnTVFnKfo8j5iQ7td0xHLrkLFPg33RiauZPTH6e+2hutF0r
XpqlPkoymNPzWNzHR5k0SjfSjCji4uZ+5/yn5rEM053o/7lVmZ1qcedfsug0CShNW9LAowH1TPYn
mPN+N2LLTI2S4m8wj2aVMtUVgsy9x+p9fR5Vq8IasvouWfPeIfA+GkLQoHdhVeF5/2iBv3Y4Lhi9
sPd88F5NAHib9XdspfXo3RjsGroyqhZ0FA/xoH6E4hHVq/aRMJF8tT9e6tmP8aoWDuyDHwDFqN26
3UUjWt58EpTij2dyvC5U/jqkgcCEdPMtqY0/N/5Qp2MXhly4L+FBSxgGOg/nsZb7GegpS1FaEPOi
9bPt8uDXpI0pgxXoECYr2z0jZ+JZxM2Yn2qdGvn6Dc+20MBbKIFUqnxsFtz7a6/O+cduihQl4hFb
iHMQtCbdNvhZklzdmj19K738B9PNmFNKkS5/GNrKmb1xHpXm7VwWPDkzXnYFM0hvEMagfiODufg5
u+ZGMgsybK5kHZUiIh5kh8Klm66qPKfznoXdoGdqWTXmXH+EQGAyNPAB2Ua6fQ+QtgPA6XfhEWtl
UNG9OLbH30YleSGE3V65lWO0IoO7aOHu4wV+hyJQ2+mEWdRXj+4/ItSGlu8q3tJOwOQjlP4+T9bK
0aOTltucAXBeo19NVPgYsR/+RDP/IZ/xfsIIfNvMxiWCvEZcGYQfItoh93UwHLkusg+eEzWjci0f
kIPVvq426S3vETGgaFs+/q03tTqrJi+qcetu8z1G32oEDB5m4II9wCGEQ1Jjj3881J436MCKU5Gj
pTOKe0UkgzxbcXGr5NTEb7h8c5NqJOWiyQ0S9wCIzqIDaO06HSyH6oRcc2xzxsnUAUSC3RaYjM9c
mrOAnLH4ISehKuGEJm4ohj/NIoAeav53SdbY3LGbCK9h2hwwpTr312xMBr4SGIhlQB7481H6cJtz
5TGuFBLQPUaOkoXibyPIqY1I4K186et8o6HuJTUVBawrcWgM2mBuzkZsjqD2GqYiaUl42fJ5J8eF
neLkiDAnt4aEbzcdxa4dJqkoCRdsw3JViFKAoFZyZthiqEj9+CJjWcZl9ZbtfapQNy/v9bpnacx0
NrU2JEbv1JjYFtL18axOq3x9M1V+/4RQvbjlDNRwKzO6xmW3y3tAnq2KcirkQ/DBK4lxqVfqvfW7
r0KuqQyoUey+MR/3QEnJ2ZsDjzEqrzajfbehSyxeIQ6SUBJK5nnyGcp5Q0BbZ1rq4Lzwg8ZlsuVf
dZwh61co+4h0IrFJV8fUr8R7nThloDyqSvmN8N37comxiPCARUhinwKRzvsOdQ1f6k4an0m4Y+28
aYijRVFECrhHGrZBb6ZCmHPxkYm3v/F+9XcOSJXLYsbwCtfELOdP3Z82c7/rfPogd7FrBR+I0R6z
utUn8oyxToQ5sqSdDN3p2WtTeY6SbkgKXQ9j4p1hUg7E+LCUsqOGW+VtqQH/LSag2ftEst1LdJDV
HW1JocZE1vmGkuXP0Zr48J7Q1/iD6KPlRGgbRu1H4sELWrALkdb9CqTq1N+7ufZH72NJjJMkg1P7
GUojEAAyApMQ7AO0gSHZrPQxjV4SplRBt32vZe7pKOhj4nzylrbuSejC9XA5ywsMYQcOmG+l9rEb
5wnNw4nXvHOLbsrj0c4vcw08Gdte3OdESEZj2U/dilIqUXXs8maCimwfE45rGa6wwu54ddeTSJtT
5GWuSZcpzgflnxVzWP+I4PRKOXIu7b3+3QCUEvMBJS8pLN5CEEmonPcnGIncaziHMBECZ+1tuk86
KelF9J8YmucCy7DrbKsZ5QfATTDFltoQuM6i8D0FTANvq7I4rlujhcwp69guyjX3DCnD5P711TmZ
utTS3rAnhCuceGK+eGvL1n8jtcbCDnXpAWhSl7kzATMpPJizhDoZ+8sxOFhpgnDTUxD4aB2cjxZj
GAE9aq6QG3s+4pu750vQ58Br90LjMDSy4liKGq33wQ0llYoTy2mi3EFCPyZJJd8SkOfcZ+NnP0id
l67qqAWUUW3z8vH4fXdtUwvSxxu2SB2vaHsC4tKojWvSQlp5hmJ0zrk/TpNpoFRsG5VoSB/Qjz/6
LKguA5nkIKfHp6uiDlB6I+wX+Q6DJrlEVfPLKhlKT1J7OXYPNDQTsSEXUOtX9jh4WzBH2kMIXD0C
SIx51BN5QqcODX3GER52VAHSsoLugM2WCPB9Oa018cirbO7bmLLDWJpY0trFeaGC32o/YwcnWu+m
CaOt022b6ckgsrMIKfX0K1h9OmOWX+A1VgIuVLrfZ24QeuwJDlLmv0Kt67X41e8hUN7/oI/N9dZB
E4KX4EhkZ+p0hDoElosC8X5kaFvlhA74aN+M7MJ5B2yrchbA5XBVGHLJh2PT6wxCOGOPwsBIxPZ4
wR5gwikGb5QVazCTeduivd3khnEqVQ1y6hsS5VYn0Ug/DGnprK5Q0aWpmOq046ONPdndDTpIJZik
usOM7MV7aCJPaPBdqOOuPRODPUa3h1N2g7w7gAurjBUavCW6ULxzlIrOCFZjku92HaOo6JqeN0Iv
Nha0KXYFoKnP31if7BjFN1E7GBUyPdXB2dVzKNKYqWveuDiI3t8Mfv/pAJhoMKKyAlht8Ui5SuHi
YzhkbelPt43qjXyULtZ1um2Fij1RIudvAawMFnRzRtcw1DNjalD8bXDvxId6meV+48d4lskw7NUR
Tdh6NK52A72CHOgsxSMlQOSJJe7pn9obvN3JaczJ3qCg//hTCepZDjoubd4SmiFBlvxjwnR5NtPh
ul57InV7dlIXCrKqUK9ve7/Fwo9sGoBScqUXQhKMr/iuEI5Jvh2tZ+NvSO72DDQeAl08OjfvrTj/
8bDJCMsX0vSVZ1E0ejFrKFYoJEafnFLg/vN4W4/0ttRf6nH85w1BoB1JkXgMUPU0YpSRo11+iTgG
r711S7vs3uD4KVYQhcJ+FT7jZ22qrFHxjXBQ5XtXebg+YczmzgoUngIyRl+Dw6+gFo/KweOrqsLN
CQZm29cy0vqDaF3sNvQt8VJ98s/4eB1dVd9vXzVE1TZQw+WvNz8cmIEVqELeP54t6KK7G+taUkK5
3kH7Bd8asQlbfIPWpxt/MNLqSoFCmjOx9a/2124AipuamfAURgEx9R4WdDbNOxUhuD6umRFUGdR/
Ed05OcNBVAOFwDom93uH24stsJISWTARBA1PT53/1GZB5DOXZZlSaDZkr4nlKYUP91Gluj3+EIh2
tzoZVcZmXJZstTaWSMZKtTVqrnAcnbSGiqXfRryHvl5MfjCblgqWOoLst3MYR+C+G2BVNWxo5Y4C
+RN+ObmngLHVWaUv9JZ0ZC+JKADC/COB2dELBvncopYE9SY+2mZf21VmfY77F6AxB9mUZvKL1DLu
ZQ8Vxo6m/Koovmk++ljOd5Bh14ZJ6VqrLCTjWPiSjuhY92OeaqUDReVqsbVx270srLBPAnVsqqwF
GIljcoK52oafU+VMc6kVx9Slxsgs7aJc0UV0qpmP46dM/i9ahDN7pVl3b1dFtkt6QOyMB8HiX30Z
q+5AfGIqQzLZAAEoDGFEfowrv2R/Fvf2Nt/cj5R91CrvqrA14YYAdvIkdlYb5A2fduCh0lIJpWh6
tIktviWMYmfeIiy9DFDNSd/FcXcIqhGz+wXmUOgVwkLMGEI472V8xD/jE5FRRlSZNDY4VjQBuqMr
pS3Fsu3E9CInbYutDqrKROdSiqOdIzXEMHHbhfCP0SF9yh5Rlj2bFYkuQovgq9qWDYjqZQuY7AFp
j+jkQooTiKklpqyb7746bvgtbjMvJeBOki2dSkr9TQW0mcqei6zsAB3Igo9Wr7nL9VoVLp7/A8DE
grXxCuLXdR4cRKiEjO6KvP67seirp8BrDUwHGiYxroGf7fdsPRcNPppnwqDBeAujAGYcmZnBTCqd
CEIbM+7EJcFt1xuuHryjOEdxhwH62pYlIKtjKmAT88pTaQUOeqfeF/l7W+s7g8yLRcDzNEe7A9XR
t4In6o6ZHnrUNSCULke3+JTNBueekA0V5zwK1WLg5SSnsQ9oyn5mKbX9QVUdHEtSPNKUtt7h93Z5
Cu8rewG3I4EjBwknBbYvsL9M6a1/kMGCetxrmLkJasO8ICLkj9j1M+1QRY7KTZuv5iqZdZFrdf5G
UHNff+h4mKDCoYKK7gQ93n3zIvum9Q7XAR2E9Y2N7kHWkCkmc/6krUytPJKAFfRyWlUWQ2Z7Vaw1
v4I6TqtijpgrWFuB6J3HYWBjMjNNb1sOdQyyGLA8AqNmoYFonmbN0YYdoFOZop/09bZPO3YTJqnw
jTAAiAOqp1T3Ff4xYEEKLIpTLj0raTKMAgHWPs+GmIaHacPJPBLmsphAa7bjfdVeXQu74w9yNZ0J
LvMnoSxyT5A6kbYOdIm8KrrLXqe3S7Pj8/WuF0w9Rdh+6TxsXeRS+r8uV+lMC6+MjVtHLrmV6P2z
OtWIr7+sZhUOUPVJk5snZkvXurQAVQmQ6R9bFyb5gI/r+TY7zflUsIWZbp8u8eBYaEkW5L1JExe3
eQ5C5H05caYkKB7uw4e9+sz0vGzc/JQ+1E9GtBemedetVrdSCppG8gaxTMz2xS4wVPbd9IItpyod
/1qrJ2YbB4vtKlJPJirCNlJv5KasnvCoyc6s4uU5+fZiKkV9kj2gG6ic6nyvHW0E+anq5NYUvxdy
IIMAOvc4Dv7ZFmwSOq3MEnJd0wFpsyFVUDV7MXqHjSTYe4K+Uqv5WwNqHCfs5m3H32wySEOJ5U0s
icSS5BmXYO1DrFplXMVyOae9fMJinfUfzDRKPWCvr3Hdvumol1oA2ZXHgLgJQzIf62I7cZb47VE0
Tfr9zCzvktcyWRneuprFMKNdP5ZAYBhK/jrv+jO6TsN+yTkmciAicVKI23dDpKZE2zLcNoI1lon6
eAXASNjHW0smnuPgpOWv4804rUuIJbCoGS4ltz+X0P3+yo1Pdo0z/WSwBDGheKaRu15rNKOJfDOc
YKSpnOAMKlWhBHo/L6kVvG+t9g5gJG2Dcx6rv3JTlhtrX9rx7qrquDwYtSbvvypO0DCBm2y6GhBm
3+JHSvv9fIQF+HrarDN7nENP9O3Mkax5+DA/2e69aXdc0PlUbq7SUQ8++cQs9TqxxTFJYXccE0g4
cMqrA271im0F5pk1hYkPzDpnAruG5XUpcWcbSDFtnUXAbvlUolyjv+zei53hv7tdr8G3yj04Ibvo
TcsnkCtdRtMq1m1/nr77Js/QrzjxZBWgOrnspEfRHSPcG2frtAKcZkN4AhZDLYGZfMDWvL0nwziK
B0P7o6iZGK0SOR+nEZ0DJit1ZuuhUn8gZgROQwZdhdyKsJybk1Ssh2zGseYej1h8TRSC8SmZYck5
aZthRnHGl3q1Qt+pE6/SU6DXERis0eVNaKPiLUw0fDTCat6DlkwD4+RGg3TaYciR5wJ5xYpxkqZF
f/DA4/crO2N4UGLA9FYIcE+DzSVWwT+CJ8wFi+hq7Kzpoe1i2bPSF251fkyH5bRsRz1zmD4LolKS
Tu2ht04UPbfpFhsHLMy4RCWqZkN7cO6u+q7EAOGWkPltR2PV0r+U/Uu6sSGMuzP0+qgVnBvdgAy8
fSsSvMdBYnjNTUZ2ffbGP+loUEHS4vpoYuAXc0ZpjhegfXWAOaWOXKXwLN7cwrBSHKMu8VqF9JsO
qtx2QOhzm2Nr911SVfOinIGy4OfZjTLr3E/bOuA6yb1ZLGo/rbaQZPVKZkiDZUCWeabLNn/oG9eT
yf4tODm0UReUaCB09w1tSFT8Xg+h1LPCcx064EG1/zUE2jvQaLig3wePYiASfnMxxykWovxaXd2A
YU0bg62DKZdmCRFawjgNW8RRufP0AtJOllE3/YeFtBvXOKcBDPTzeBVhrG35U/U53SMmOK0YvZaF
xguSR4DiK1UVtWN+fe5V4uWjM+IZPJc3J2JSnaynTUh4UnidsI4JdUD+aSRKcgbfZzODuhi1AhpR
e0n7InVexYLQgKNhdAZi+ZExmlD/rf/txjFlQa8+uTE5YduYS3JzMqbUPVONTotIIt2Nv9Vsks2l
WtzI/2q1Kt5WRRV5xPZORGt3+TcRZPQ6c4xe7MmvOQJKvP6+1oO/kBON7PB523cyEqgCxt9OoKIO
Txc1NZXfMJvO5IlSvqK+CBUECCJOJAjm+UvVTYxGV0+gV6+gr+xR5pCIb3l6ztrzr57pHn7yaMGF
8/4tVt59xw80iGPdWK16JQAh9i3Vibn9aJoHtW8+tCr97x81qrtR5NfvYj9zYCU3Rmtrw/Hl5nYI
cacos/7qp61KiKFelTPIxmQCQFCj8K53SLjTsqgh8lw/47ho0OskmoeAYRUB3YhCz87a6rOqG45v
O9zAVc8PEtxsMwkY8s12kdVRmSE4cnhfVuIzl/YxxyhG+ttfAUW2yVNjWsuTrxLoPgR5PYsteNYu
sTCx6Tb6PMGFWcnLg9Rtj8em8YXRXLzyoDf4wzwHqm7KO8D8ZBjW+ZOq4OGN3Z6+ye+AedXn5Qxw
mq4Op3Pk5jI/1IkBtepFgxBbufeGNfPsF8gMs/1vxlU+gQfQprf/dSKGpfEkx0kpSBTIkzBzoXuP
0EviIYUKRrpat6NOUOh9HPUOiPc+0p88/Q1zCSz15qXNldI+z1Nz1hF4+hYXCS64aj9SLtazHHXG
cQSq9OyZRYI1wuhbJgntSDjgoqA3LjtDO1NUfJm+ESCtyoNEPD7S+LMAj/XblIRYsHJVItjVNZgg
MjxYTtz6caof8f4+xBHFKybklzNbTosaJhadp9AmobXOoTBL1iNWadq1V0mXDk9MvrOY/FEWLD/f
oTOadi7qbmsNMOWlZ9Vn7wjepMqPxIfD4+BHTfgkzfzr7kecejYM47FA3gfxMPDiwWlbR9LmpHSO
uo8+FiaO3enA03z2X1YpJVjrucZbVCqzFeBrImxkATF/jpgOyn7xOA+Da9ahJXbStaTY6K4UdXbc
Xh/1hGmSVL7NtC9WCjejdPpjEY+UUdn4vXq5TAZniPq3UPKHXNLFTbDpV1fFsTm1aMOWmETjMrcn
KfJmf/vuUEuVVaTd9wvBd19NzGz8/A+NaFL8NEPNxTUUsTeQaGsRX6TO179+q02t687p1/UOYI1d
tZvNW4yhzO+YSMs+yWTr39UMfz+kdZhCWBf8ZKS+Tfwx27qZfN8zwleIn+VC9hTnI+Q2UjbB/l11
mk71QZOmuWDaEmkaw2sn7whpgG18aTUEPLvsCiS6HYstq1Ol01iODvct+Q3T0jJxjo1SH6f0Fwi5
oXpdpOpsTdYCtfXzSNuZDaIctbgnc7eHff6Z4XgN4IKoaSUFcEi4mwtQLPNl/SNpum0aa0YCliLQ
60nm04bsjRbG77ZK7Ka1UrG7OXk1YT9PTWHb2RJj03UoBZXmzHik/Nhrj5AzfXqHd3f5XSVCkUZ8
lSptzf6qG86G6FFUNE1PePzqo76T5NkdSduCOLiu+RzJsZ9DHI4tVTX+NWZPf7zoZgpXkCX1bbDs
AkEQtQsY+0vAP1HHUa9p2JlQ5VootAQFD6Y16tHNrZo2UPm2IOWNFD8vSR2iiCcUO8IwcycHc7SC
28lzAqLtkN87SRO3iti2ikZ3U9KzVfXzgqA+04Q838g56fZ4M0znRCKsvQpoeP/9TleODwQJ/Oao
n32eguwlyvuyGYCeRr9lpgO0i2nDtNGqTkXk4PPxYeCl93z+9rtPNqtVfr49LOk2Z/NGZP1XaIE1
3hEq5LzgexflcgSlpqP04AGJ7vVWwKsj3bjoHd16hTuHuAiaCeBwddkGU4E07bi+ysFnpsoCDU0U
1z7+JRT2PVc+efLKfhsWcInIWum6nhHVqxVXe9ZEruYeuvvJ6moV0Ga7NQM5n/5rdUewsTs0x914
AFTbwV9crF3Z3H3R6601QvMast9X8iw5r29LJp5SAFRYaaNpMSPMqHymogDiOte5IlRq6kDct0Zd
N+Q/VfEya1nxJF4xcI73XZfa446dd1cwxkSk8hpc42/noXqEbprDyxXgCLq5vW7H6hR7Zp1ASjit
CYyLaosEodYuRwJm4Iou7ZZGJZ/bVexjnhcRd59iu/erAaQ78oRkV/gn9vSCNbXdeIZTBMIAvr3v
/Rji5Jjl6zgez3uA6lBfnae0Yld1I6kPo2sVH/fnRtlNE7M2mDdvWiHNwk0UM8Q5UsxoEohyTyfm
+fv0J0DWwwqPl35yAEe6aWTjlFw3Wd9ruZz3z5ZWQ9Flv0AUBcBX27ZkKxmIw362ONi1f8gBxvwl
GhIcG9+yMb6QiKjvjdxzVlbjYHU9z65AF0ix2XBhGRHTmEe7vaW+75/JtkVVbF3+yPp7Wb9XkrQR
VEyMoMAGztML7KMmZ5UExBqu6rRAXNt6iKRQpK3cTQhJm3sl50FnF9ogTim61lU1XCE4ioV7Gm7s
EDXEQMNv7k5Oo5rsm/BIxs8tDJWcagoMle9VG4c/CwRbv1jbJvCrgIfKq7rTzuKhKEckXTcsgtwD
Tg90kjWzAYTxPrypAZb0Vt+WzztJUPwp/Pq4dsfoVYq6nqM0K2k58KvW05RrEoAQazFw2psAOqZC
Cijayg0Ly2UcxGNtJa25KKoeGMOOE/8dLX3YAiDL8QihtvkgZluxOTEtMhYY9dtzT8eKBhz/k//U
d//Rl9uRNzWFuNMHeS0WIK+BoTLF4jGPTefjIfAYTLaPqsWcBOtGsGKNUXwnbiFQTH7zpEEGVRTF
UH1/4szi7f0ezodGBH6VgDaABTg7ikiWYtvNpDMUOs4iTM3URMgnam5N5jiE0FyQLp3jAPFclyQ/
HfHU2hkGJfvkTsNxZJ1msRRt5XxjWBmmcP04uKT5eZW4mQSV8Xtn13mQM4RSzygxR3zkQCsV7t+m
pWaUpVgHtyfEgf/yG4gW/0ELGS+ce0yR5qiLcr8Xc70Son7LexnQRrhVX9DnzQYZvFvdyNaMdYnx
3REokdazx0le2SoMb6AdrELrEzJxDW+1q+zwo1E1/uVHxDmIrhejqUnAvssG/Ns8L7cG/P8bpbji
2tNI4/l8RRxp9LSDWskeMozFfcgSkvxzQBWgG7oga/Rd+3mvJWhDr2u51sqtzBwVfEdC+dCXkMbw
Viq9T5756WYAHuBMdp1+zKWsfQQBj/rNJmf0s+GQgg+S84eUzUXpnqyxOLBoJELtsYH4Ko+dsEj3
QByWHaiOyl+uzK0a+ru/WayUPFdsNlUA8KBkIRsnxmfBm2Dir+Wa3UrHF1zNgIUWHJOsgL1GJDeE
q7YmAs8jiRHct3+lmjyUwXNYVa8QxxPMmSW5bMFslaTnyh/NTLlJUA559MAL4vaAagEP0Tzc8j3X
q95o3Y8gqg/pMB7FN140Tad5mOMqWk1M2uLqJfYoATkznyTJxksIRTXQ+gNnV/F0CovBAnl0iRZx
r0aC1PXcjg5ESHxADSEEHWZx/GoTYdTo6VyoBf4TxGMr4lpi1rT5aACUNrw/Buf91Q5iQCA5lVmE
sdSDSlLErOMYnDIncSQfsaKsiujOgDRL8bDLrLyX4B1Hr0q2CPpemRAaeeQusGdXG/eY3D+dMeXo
0M+CsrQhBdFI3dTS9y2KPRdL0Zwh4qBtNtD/gS1M8jJQPFpjVR53ev9lYSgv36ZaFjkuTCs6iwTG
zfAcqrIzkDp/fwJDdvHTGFX2WFYHbFmL7lgW2IVNFkG6DYG8WAnH2Fq4NveHOE9fd+8f+kp/yC8H
or02UAJlh04e5ihqM+5TnQsxoverLU2ZHm1hVT1uwjkpnPnz+g2XGSGHXcxOk5ERjTDlNJk0LOjw
PCV2i7cH21U1NtWr0U2Cjnfq79d7zf6IOK/KsTkxNQg1BpOFGUTHhRFo7vNDfXN9FzrafnG3XuFU
13WKLs3wMYZp+hBue2wS+5l4g5odp/emxf6iwR0XCSFeuqu36Rzn4Lwsw6klyOoFI97/YJxAMZnp
b7QthsOneHuoPC2NldxPCfjFoaNslFtVnYME7AFalYDjb1KBvxieebYm01/kKBx5yG86bHkpCEG9
O1j6uChF/CR+Gu+xqKmWKWJXhV14f1t+fAjlhVTkSO605OfxvTnFb2QbwboJXvXVEYM0PkubO06I
m15PlIYhVN5wOncvG7l6W4lXQ8OfsSFE18owkGmDKdM2dmowsFc/Fzy0AMs5lz3mfNNl73X5Oz0F
W907z2O5FlWgNIGjRkFPVOzEzcQH/yaZ7RUuLVu1ECOGVsLVq7D3B6mt4rATgox8ElAoLndlwC+i
spcXaEphcLlBH2B7B5WttM8v6EsiY6JQbb197dsUV2EDfxouQ9U/mqKYxU4zcfb0TFbnNSQkmnfl
RwtXh/67j18fiWZUQ7pUrHjx/FmcVMoLxjBDkLQBoUq9lw0wpGAwrQiy/OvCkn42X6PSniDn3MOR
xUqrEkMovR60THLQZnc3dZ6ErjkyN8DpDhImflkeIVGLA3t94Nvj2OR6UDgH1F6RP0lZ9/m6FQsw
pLLMMZ2my7s5OLzgq8g0GtEzfz+YSi+mdUlELLnmr1XG6uXTK4c5S0KJzJviGFp0wrtpjdtGBPzo
S58tkYNBkoGrJPclFJ9vPr8Q5DWT5yn0y/UebvldHGiWUlpLQn01EWa3rFfuOiqS9IlEvpgLH1w/
gR5V7dc1Mrt/oYTn8cZ/GBBL7nJ3hBf6ZkxQf/s18jCaHw34XzVqqaFwnjQinjSbwAhzb40zOnYp
p4K4zP2baCEL8mLBP7XU3J1nDGfcm5JDAJo/TPnqA3olpwx1XM/kGJagusq0CCz4T7wPKJSLJ9vV
WGipt5ovvV5U3auUM562vJteaZ4cFVQUXFU9r3DNy7fqjzBUPddVMzT/v63XeMWAttSIc71hWRSe
RjpcXjxBjUF9rkYFVgkJRHF5crR3/2LIflQIlcvQDQRFcjTsLVTWVKlppy4mQKvukkiNCft1AcG9
nxc7YNjHtcq94sSMJAvRm7zwm1YXRMlgFM4sHQkorlrsqamW9m4jP7w+9iFAO7QCSpsV0f2UZJNi
1sJ2mCHXAoyL1vZmbkq01hlBasfw/M1r1s8JzZnR9YmaEylSi6zhpIaXTQXZgBycW6vNWp8kiIkm
9JdWmSLQLUGdHw+nYqU1zLgBK47k+6svRI+k/S1dzDrDYOnt1O6090o29RM+2ygCbBWAqHHLpKsc
4utvBnduCezsbxU7zaZ5wbl42HYiuQVw5BOhkyVhgI8sMEPqrk7qQYD45os2Nxxa2ml62xoUFe69
e62TyVnXdLgxbAFycmYYhiLUmRb6fRLgLiBnNRIjJVU6qa1x2ree3Itqm0SzBpX7kZakU/wJBEfI
kmvTxAqNAmJHaQgQJHv5N327bqd7FAZdeOLK4ekRAtVhwAMJRpk2mjx/uYeZESSAl1QJezPbs0h6
0EZ4rd1qPIcO08PURwKGJPUNR/fS3/426x2qlCNLecUk9nQ5wbPeBJS3kacJZGdnmtNyTC+MzurD
7WFwRHArsK7coc5v62gvCZieTpj7mMCsn1ytD4A9s0QaDoiefX+xd0wxay45mWWFfnS100KUcXyg
mEy/yqfkcoI3VlwpGVdwYpncwHCLxb+WdqAMmH4O8UJ7EiJb/okzFCBbNnExSRd1i8jJsC4q3AoY
vdg/BkyIQuzxEcwDHTOaScEwXk+oAwJLFDH+hDxGv4UQzzqkBi2KT8eiH5G1DLI/CRCbvMSSN5WF
MpJxn/xHpnCoFFH64ijJKcpZlq67/smUyYeG0rpSKrKvFhqbS9b2woIkelcd77KhcK10/y/3akhE
5NHi2rqa+mxxOBJ3ixu8ivRgN4Iv3YCmKxM0ApUk1marxneoDxF4RMh1sbKE8MnyTBTG5sN4aKUQ
INTGGAotkdz45SggoPk5Irh9O2OpIEqZipl/jkaeD/nDdSyzBIE6QKkmPr8sl2/lZl55O6aAbfeV
BFK7c/9+KqNDn/y+X1ZzzVqv0ji8ti3SY7zqkGJS0qLW0FnFKfPoX8ghPptMzIcolLuMy8QOOPx2
Zb05fD5Wx0dSHEgfecY7wPNEtq1I8CnBWJQSWJJWOo+irRbkQqmVbaz750Xwn6VAzplVzPoG4gDy
eq9IwkOgOO3yJLN+OB9XYWE6+glrSnP5rdg+JBlxUezkSJ7jsvr1njXklATueyrpm81t7CnZdgNp
mD0rN/zufVlyL0GjTfJmkuDADDFpR6HWOL25PWj5aDljbncPuzaUZ0zrVOCFi4O4DY/q9Udq+4c/
Peh5PKcgRMHx0Kp2XDzGImt0p4KG3oVZlwBvaPqBcwmBmrY2u42f28HltbPoQCiPI81mjqRUE5Ql
dd7feHsB/pqDOuBm0E5NJ9vLwSM82YpQLpkO6SZltMymp8w2DSv+fUVqn4Lvakzhd7CXxx8NhdE0
7SuqFrGzIv/WvIvJJ3P8dEgga7gHuE327KNc/xaEcMAwCXdyK/J6fNJV22HSw9GvvRHqjkVuZfh2
Q47+M8+o9TSQvoyYW41FASfZ/6Dc8Vb1zNqkltQdY7y23H9wUGzixe/4jkyiI9/BGxftMhXrlwdb
dPmoRM+bxx5UGxbaOhi7vajnFTkcZ9d2TYo/y8UETOGKDpxw2GliRb6XMDezTBBSRZaRwtJkA/qS
6lj9FbTfckwNiIQYAuLKdOnmBN8GZer+i9NqHe3Ah1bHVleepn396gZMX7mRAWe0hvLNHI62xQb4
FcmZoN6dEy9LDZkkx86cr7kuHtmywc2Xc92LEor0//aTNbPicUbhq0kWN8UsiRkArvQtUo8WUg94
zcYlP5wOyo49hCuhUychtCD1/mZa8Y7/wYKZC09OwfVmfqp3KNdfhYwOSpXqKrWTPNShz1ZprHoS
Xg9IVgwICXUfPVJQlpl0CXT6AXki+gEijA13SaZ/CORfk/f1h/WOEKxbEXCW+Y7Q8HA32r3NnYmX
FweK83NoUIhATgnQ4Vec9lyobC4Zzi3llfC2iPkLFGhj+zE3fPGIRqUkeHte2/0LUDZ57jIdMbf7
DUHIOQivHoMDHaj5KI0r+v/0S0gn15cBRmcyNMJQdYCNLXLbOe9W6oo3N9XiE3sWgN2O6XKlkn8C
MrJrngBxQGmpNJf+WmVtq8ytgjosNFoqM8VqQvnwMx1UHXvIWem/Qi9PXmbeKXpN18b2w9b4wBAf
SbsJ13eoDxaapNVlaOttn+RLhPlttXC5QIerVbpOZWcm851whWzuxAplMhG3Q4Qc1kjw1NHvMwMH
aHNZE3w5d16DFuxv5mfVMN4fOm4j0PdjmzWYq72gvh3lUv0T43KDPXHTC+K6/agLASS9oAB4EBAl
0nDv9+gzsqINigIA8Th5xizGVEMghM8r2mDV+cIiJJDxLpXAhdjnHKXNDNbinFVgNvAxnYcEcfNi
jVdxnIVAJan4uVqi1gcNN5rVErAkvO6JZCNL0OAM+5IsnSpA09TwwmYC/6FJynFfF5CYJrZuMGHE
XMGMjxhg6p/Uih9JjP1FRK0loBtaLWTQuyPcYapwnIj+9DCDiWz5BfH+cGyk9upUwhS9Y/KTfROZ
AGvcC5K5EKlagT/bP2IMdUAzeK6ES56D59rVx35JAcWftVDUlGBpTNLwpQEul5nuwieg6gsYbLjO
p+5bMFaSU6Dppmm1RLP1MXW1RUpZUT2d0dnRJ6WrrV5VOMdvaHCTgjUlEWSi8ugJWaMKzEPqdpH2
27+/rltJuNJilCdmF0h5WPBVjT6iVU/I6qghJfAPom7v5iOMQDo6SALWU3IZp0CtsFfnH/7WSdlU
6g4Gn5V9o6tL9I1WSVHTaQ8r30SWyI+OH2M8RFXU26tOLIt9J0IAqp3Pktnx3oPQ+7vHmt+0oYxS
nHDMeW6IWYE7kF35khcGDUajx7P1AbOJ3VaYEcwsL0zkAfyWVD7tOE9QTVvzQh7rOB+kvrfIpafa
p3oaIU1djvSo/oU89ZMf7V6tEFQ7lbql8QlM2x8zc9ATGEpUIB5U5+WfqNJUO0wTPNp2f7UZuPiT
WEcC2l3Z+XGrBvyndI/0eDVAiptN+YRT/7ztw+uQe7kdhi6GrELsV6D8o290idatANyKBmDXQBNV
k08vkKUVtfaQIqznobO2CdXRXy8XcF6TAauW6ByvvuPx0bg52ed67PuBI/SvgZtMLrp8S+nHWLyn
bWTJmznl20o85amf6KOVGd5watCS4g2+onEEWSUKDmEd0AXT6lZ06Vhrms5m55qJztOHHiCEhjE2
PEd4n5GUVMj/W0CRNVp9Yb3fbnmCma0EaT9yU81F14LcEYLAZTDo1QNb+7Ter9FG1+BxcvZ7koDA
lhTP4HJhqs2oFcx1SXee+84uAfz5MeTK+Vj1PMMQ8/cncqTL+Yt1gNrYie+5JnfVrRYHOuK2uyPu
Uh8a0UwDhJUGoEVHpBGgEmfyjWNcb8zc0yfCtm5HXH6viavBPz50znQswJSgfXKg9G1mx2caAGzI
VPXpktMTnS17xzt8jnzUWBe6T7ipNCN9VUld0E2h48qKJiBtaAASlamMNpzUszFM3B/8WGc1JaZD
2D5Qivxp3ZwKZBkdxHXOPLx1iIx3lUT4oIw4xbfGFp+64Q5PzM+C8TzVt0c+mdIoEnaz452jvOBS
FVoog8x+Or4usP74SMZ8pF5+KsVT37GDKW/2WJTodtD1nkWvR8WdUWFiuIif2yXJgDcBqzd2uA4C
hU6BzwI4/29renLz1UDlSJaksmNvoiHXP3fn6GwsG3UK+2OXeNYUXwhFvtZtt4QTkWuot5t8Ur5f
BqPgmz9BhqBE6eYmCOIcbLK2Qb3nNCGB5UPESvKGc3vz2MHS7EwrjTP2WnYQhdnfhq+rZoCiXQaD
fPhc+5izHOxYHb4dVFHbkkIY70YbKypbO7DorSA2UcvVgKyHNHnXoqVRTdsmWQKlHdjXHw3JEjyK
1K8pr1IuKCBM3EsXIrs+49UgR5r4H0QaN2KLCMpqZGQY5M54QYD74Wdkc95hQkcv8i5jF0yYwEea
+fwrmAwtY70jpIHJm6U4nMdffy7QycMDYmSNDBwfKt5ytjoX1JXDRKQ5L1yeWsiueFU7x5SQS87W
r9h233eMDLW+Xkt/99FEzATePDca4Lm2r9zZl4ZnHHoYF3UhAVVHMnyOoZcDk6c7i1aSxepzxLxr
1f+BXnqSoPJ3cTrMcGeuURk94HLTzEQyeFuaJ1n9dejHwLTPlgbmz0d1zXG4JHHRgqlzdGaF6h7x
NTPjDbZnvk/YeTBz4YNZ8ADPn5dskAj313fbsWX7GWoN25XkO3kfG2C9T1O5Z+SqGxbx8fj5EPGU
Zg0kFFAV4wHNTolpsoywz1MvSVGH4z/ENms+iTtpWofLATjb68qPSm8bC99pICBQ18uTnjxgRnvP
ND/UYY25LJ8y7jx+C0jCYOw/ujHNkPOJ7wIX/+djX5PiU+lAqUcZnRMhO1B3jEQN4AEy8qJ1kr9f
sl5rRscZIMRexZF9l3MH9GFqY2rer5tGZgjGWx8de1yj83DQefDUy/rXTieMhCTF8FgMUDwKBIY/
ty1v4arq9z7KdERicLQwh3hzqVltTwqxhxqv2Jhp3Sju2ylJn6avDqRhdy1YJchiyi7NrBi/G+Ju
pQC6zJD3fink9GUCUp7npmsw4RQo4dZDzptaQRXh+cLbOhQJOm5W4S0Kh6phe6k5kthZbetcTtQA
Qix0K8jWM+Wq+GcLRMisKTYCByRPujOH5uRZESCWkpwaXAnqzbXi45KYvrenZavDSXtv+5fkAM0+
vxeTUln//zqpnPBWvRXE7KSNjtJ0qzwqeO9Wvn7ggKAhVRBZLpvSq3U04KdBafT5XWyjwGDvgqRa
wAG+QfH7gn+GKcIp4lDzjDO3C9q/LQ4nKQvJ6QMv+iZF3unAYW42GGJZ5UcpzQVbUSNXGIKUJZ2b
YnNUdibuKfAo9wTT+V4234ZKAAcl8eF8wGRmIqbGaLj6Ers9ComudDqZPEeKQsVzGpBb1z6LF2B4
UbABrrmOetM9zvqrWoIrWIjloFKVQ4lT8Wr36fUDTsN0zvC5r38J3CHh5/wM4zRpjBHhghCYZEXF
L23ClpQdYTYdZ3OL6qZ94sJM6YhRTfRUvEVr0i7Neb/AU1h4R7wEZdQosf0ZF0zwJ4bJRBiSdNDX
vC1pC1XVc46rvGFde+iDgwy0xFH/UUyLvUZybp7WVmChmehvSX4Z8dPDmsuL9gILN8Wdq4Ch5Sf7
FJnWJR8hKF2LsUCgH7zltl4RzQZlHZALs6L0OXgfT8XH4WZ8IwrreSVAe+1iFVU+4941O9GVUU0F
yNoDfyPLqQ0x65hcoxsqNkFiS7GCWlbbxmQG088jceX46CmmyK58DnuaurLkPKMBrV61RGprrcUG
XnRGOSIEIhxR5ykkCtZic5jCniq1o4NDVEgkGwIv01xSm1+dcoF5lZasjr5HwMGapH85QloQiqZI
zYKQutXLxbZGUz87IUHKo1qctXEtwLs5LbHq3aUSxgvtkZGxGLHQ611WCE28sdM1P62bxn39T4CH
tgYktZtzAc3d4/FNy3uAPIN9rgFCAYfg9Ftnp5nXVqQ4vISg/ltB3tLoTh6Jg+6S93EQwfduByZ4
/EdR8HO0C4fe4EgEWphX5AN+5sJJLoht7A2X8z/9Fc/nq0GTFpTRg9SG1jBu9TGbdOyR0Y/8gFpT
VxV5XTKR9p3RtfHBInJSh71unAxw3CjMomN0LzltTTLeXjWJ4IZECbS7tvBpZMa0iOs87SmsPj5o
j8MGarNMSPrkRhOnOkc4IA9OSEZdalaWHO1YEu8F28+jYqdn8AEe5FaQUyQnUHtldD0NqNLcASZM
HyoM8VbaKmLhxdzN9F3y/AqDpftsYfhmEHYDR3ruQiUNf8Hvi6/mk0VeV3ubjhshoRTcU8EV3ANa
pKnjOIAJf1F1oCLRjua6YhlY1a1QUJtvwP7hofpUCp5V21S0d+bh39wS/gzV68i2AACxumD/MX4R
jmFYyF7djbFB/ml5iEA/X7yrKXet61V8phfzaemIyyAiAJxWGu7EFUJ/DiG5Eqg2Ush73SDS83Zs
58PeL7sIIZuru7yB8HykisuHSISgXW7BZsMmFnPZLZKCxW9kx3VQIi8t5fg/Nn7sa4ZKCN9s5K6P
YEiIeBDJAsp6FWD9WhSYh4leGZ5meMLE6RcaF5E+V3zdKZSB3U0JlwObg7tUPG/EuUOqTt7d69b8
EKCr8HWLg821mqnO53g5nUhS34L02z30Ffef/MKpG5HvCnKZvMfo8GaIUcYDdsjAuaDRN7CYtF1d
dj8aV/WAexukWH0rwPyRvYrrllXtCP2v0wFnIfr35W9kC1wZ+wEobYqfq7MRrG4FQej3KNhYq6vW
8nH7kftNKuC+4r+hl88rt+fpcz0wSiwElP5u5Sn8JGPODJtByJITFwe6Md5Qg14REcXrr6As6c6g
Z2WE+pBobkSeR3uNbArkTos85qqRN1rbbMKGqupU0URME5Jdl9kBGKxxUNKRvlWWjfitpvszrRDb
BVwiYHxMuCCZtpbQ7Q5ozEAw/vBKu/s+eaxHxKId/2QK4Vo2Po4glD5en/j+jpIwijrewZwPtWK+
gHpDYN0AbhHR+JuVJKmJgky5McAnLJrM7zANzdQhHR4I+lHU/5yrNmq8q+fBN2I29FVgl6Gn67aY
wqVFcNkxKOAJSjPJPBr1okzJjgM4Kuei0hfhuy3aXGfh8irqv6taUvVDZDWVg3UHc5n9GipyGvBj
V7V3Ht/pFwiD8bJHn8Jx9EMJswOnwhPESZbskClS3T5Vk/8fhCfT61JWs0Ce1zinCwUgXQCD7aL4
LBAGfZwUV+gl5GpfdDxYFxAHJnYeCjqmAFDuQ5xNfDAI8HnShVsISyz6Pxyt74fURnIsJFL2ubEP
KinKdavPSUIGVddodbwrb58lo3QDnDF9FP0mNbDzdrRcWvQsY61my/lqwJNJYNGeq2LHXdb9IFFC
WtHOeeFMtml+N/T3YFmC8G80Z4e2JhuBRUzWcLy5a9jIV7NB7HTJ/NFdomKYQhd/PuPVZ1B9a48k
4A6qlkuF2DRsg/WIpN6hdvftwpZ9Ddvhr+O3IQn7B42eQ8pY+bXJGyQd5q16NefzmHKvHTFNiy7q
H0ZvlLF8X7Jm3a4vfZqcwav4yTEjWSQA5UmSPN40INNzqfNXI8/Mye6Vv4shCYajYgUi68vu2CCf
qQibw0X8SDFK1vMyqQMmZEK5g64kMYOVTeEhiGCszYTUWy8O0ZwkJV51A4qzRgnCgyxMQi8BsuxX
AQSgb1FS3tWDgNhKgX2Bq9Y7bxjBNEjHXUx8LxUfPOVpBcaXyqB2gZitxoP0YA1N2sDi0NoJlke9
U4hMf1F38qOIRNb4XJcNMTOK98srGBgGZ72bPc205APEzw12yqRyRTBOyRuP2DYF2z2j0kVKaPD0
7Othoht4FzthLdeNrvZ0BNYPhv83DoephmvcXKvKe2/wMldF+3nBwMOlPQRhzyv9QVUzDBGUOqwm
t3Q3Xg/jP1akuf8uLFPoYS67HP6Yy8PLDGDM5vlPft3SME4DjIIzjau2vyIqxbitGK/crIoXn+i/
WIYsXFEmGsJ7VeaZWq7vuoQMxy3hqnpqRMfyR1mcuadGN7nXLLTJk889omm/RBisL4roULqjg2Li
YPmq8el7RwA3hvomLu1Mngiv9VFJVIx9k3Nmf7PoDHRsqr14L5+nxi+mAXEfMunjua6qM7eBJroz
U+WkjqdrtwO6KFtxlzj9eFA51A23qFejd+iRzLET1+Q4pR1E2G8OobBsagt+UyFX0eNJ1LtILTnL
OHLnmSN6blIh+4I69xP7nZ6OsNx8jL/hmorRtBsvx0/MpEtzyCs9h7iOi98GuwI4QVxge5QdJfyl
siLfFOrolp9vu/j0ohL6pq/Oo0fKzyT56dYqmVkm2R6oU6sXa94utIlNrirwjjLDRyD039xXTSWd
fFRoHX6yALYSROW4XYKXDplP0F35fc8KmbNvu/D6h4vQW05Zi6RGKMFcBICLmd/6xzISm0qFmjty
32rQUh1AFOhxCHRmJM6WpupsZxT4Z7CyuPwJZP+XLDNnFLsjqUogHNsieflaGKS4+915nPtn56Hl
ZRFrWVUx54p+DaPRYNIDfvWNh0a0TiDpLwUdy4aosCJDxS5ATLTwMmxbZ/c3HOOHyCCLiK1j3prx
Jxu7QtimtRUSbT1RpB42LTIQ/SNlsNoK3tdcrwzre/ogW/7ErmsyRkaVZA1xAVoQO5HmSsi5Q8dZ
i55SfQ3LprHhFllPJZU0AHgii0hy5xmOgteJ6RMo0IDRwdXYna2Oo0bN9xnNfX/aLUopH9Cs7yyG
9cOkmhYWFUGPIRJcoqCcA49tNfRoV44MU92aftEeLKu0WjiAl8NXQqFB4V5sdiCry4QhyD9b08ZQ
N1cfAKlvESdjMbXW5w5G2YQnHmAis6h6gveh4C3pGvq9ykhVwL8Lb5izKWZaIwkR4ctwnO9Nm4QI
3GKCWNwA0WsM0feyPXonakHDJ5i07t3mmCC7iaw/4ICgSFz7t6toJIpNvv5TPD9Bur7IF8kUd0gn
QSiEiUHPXkGbh7d4MdLorOuHMY38zUlHQIW0HkL1bj8X+bI7km9Bjgs98V1dyAPqk0XtgdE1EPT/
oFtqOUw9HbCrcSwA6DoH0JTapg1PMzzTFbBzQm9cqiAAQbwJjLKVg0sxduR/ikpUBu5eJTmxHDOH
r1UMlgmcWL98ZMz5FBieR1zFSQR2Lw7h8DMaz6iNf3v26FvX7/8F/yexnyUKnxxvnhJJnW4lGY+z
+dkPJIYL5j5hUn7vlNgplHfomEGr0Bz2ZNVMP/mR5Nk4lydjXdyJc4gct80tTOmF3ZTuSkpl0eXP
sOxD0ZkT/CicgFJpX+1TnZfFoFRoJtA8EG9On5IR6RFHAk8Uewla9IMh46Vn8foa3tftAYJ0N1dU
joeShlFEoQ6SvYBOE9BP4EFjHwUiG1oHgZoBOlDNCp8ySOFSzlQKGtMjemC4emBFbRfGQuC6fnMx
lXhUkuuQOfAi7giQmcg+WvgYWQ2I8rBXt2FJ0Wz23gSa2oKhjZBgXfODYDvcHuvV+iuHEjs8nlRP
ox474wqlOwNR+8c42hfI8JJZi/wzXQg14C+patJFY34t8zh1QsgQ+kfl3hOTgC/7ACC0SEGqeMHT
GvT2Vpxgr/Y6TT5yVeSv+rMjsp1QTv8+H2lRbMuXbqVTpYspVZyFfH0f1RaF1JztoDh8ymD/pB0D
zvLHYk8BgoF7WMxaS4uPS00uAEBpvlYQDCfDSHVIDWd4gWzKG0YOJGoVxY54w5pkD/ofP6ve76ZY
Z2EWsEQsTn214XKUF+38pdb+aRFEvDQOFmzTnX4Gl8dm8OwANNxJg/gGPDvI3IOw1nPkvNZyEo24
n1WKgSg2XVC5Cwkts0O0f9qtwzSOY2HR/dP6qCGu7XejBsFgDpbUFEq5idBp4aQ/cmkLKgaxk300
42vO5xBwgJMkaamwfPZL2j4d4i8nF6VCMYKGXOG65RNnqoLAxp+du3tWwKrqsVR1Xrqc6kL/RT9E
A+qr7kwHmksrKTp7jRYw7Q0hBZ44OP+2oKuxK6zWKmG7RPsajXxqE2Mx3D9X6G1qjoTpqu1NY72L
cOomKxJ1B0Jp48NFQRjpDaXgJFkpz80y0jopwyWhiKg8E3cGvydeOCv9w0kysltFsKTfi2F4aDkI
884jSCHt2kc1p1rW9gUhLpKuByEk8qrEGeNDiI0qzPdoz8D2b+ApKGckxdGHBGEV+2w3FfH+Pa9n
tDwfQsj3wcyG+K7u5Tv87KFPYP7tzxbQ+BMJkzwXfCCPEicAV2Bp3t2zFytU+mmKaLczaiD4ZtHS
2SMkIktrlAcSu7AiuxUhAREKFme3iP9MFsae60qoY6azsO/oUBex5fWmjaRQvmtLdZu1oZq6xuoG
od5sAdqx9aFiWJPZIHnCGhelH3Kuk2kHdzfc8zL8YXjkiPsxKT3V71Q7WQ0nwzfWn3KVWwyVr9Rv
2zg/AWOaoLOWYYEmKehgWQHYwyIO2WvvUp+0VXI117Cf/mSY0/A+ip48VelbI2vonxWnYLPQmhA8
dcajlNfhG95I/uqCjZljRlgRRDNjQiS/aAz6K4ZnNjJgSpe+5jKMt3S7ovCII/7hNByvGQBB9Ffe
5T0aoHqZ9YD3Z4UO6osl8XYHsYwlk+LYFPfa1AB7gpazeEmOwinTL45B08K4YuBim12aNA7D4cMN
h9JAZz7VSnzi/ypdo9lyRqMkojdDPvvWcOp5O67yboGHP9gFe8EnZqmGXMcbs7dkr7n5LfV6czRx
u//kh52oBRlN00Usshn4c18Dxhe5ReJEh/rR8IE/2VO3Rg4MX5h4VDMpq9tQmHl48CvaYlav9pC2
0uVMcfEALy0NwVwSWACfdk56Mm5Z04gvJTjPigXG3zLXxev09aux2S4/XsY55VYQGLKIHGBRY0pL
nBBdtx07x+YstUgQ454W4qvM6EG1FlxBXW/hT2OzEixRSLmrtp3IFtlU/s4PUka2drrBVRwFaZS5
DHeNPnx1aUq9kAoIWPXgWwC4DTuQOl1aFCq6cMY2PYZEQEJyZWGxvRyv0jppyE4jI4+eGHebcLeQ
O9qNsqkK3v2zNkmX95edDfvbFqTL7wRNxRejJzL1hThRce4fxULyFKoQdeGzlrbe776l01oFPvi4
CcMPS9jFEZmXmf6juCS5JRR3qEV+XVEhI0N54lJ7WIb5sSgNYYE5WkRZuGxXZiqJ6a0RFQuHyw+g
81ZKnIGmXtsoZkgg16yg+eBha4YcpQRFgG+IzzC/Qr1z1DAjVwh60q31P3ftuvm8B7iCWGvY9Dqq
rZ4HvKaKvrjh5Ew3NtPE1JmkwkCXIk6FClfuazqRT51/USlUr3a6g302jbeEOU9IBssasfLFHcDc
uF50EC1TlK0aYNSKY2Qi0Pm+RBKalHs8sNW0qEotHJNYfjlxgCufu3L0iylUNaA5Qb5bY16QwIoW
V5lZiSFCRzFXARaxgoTWGJuHmmpgOHxnEKEPUsZ5J7QeBcWrYn5zIhVzgR57QIi0xL8MNRrjO1ua
LJjPG5iSdZaC1hOQXfut0kEuF3irDiUUGSphGWWJ5JOuPFjRjRC8vlbCbjCnhk+KxCvM/XEfEkcA
ejPQ7qn9KObvZ3U0syI7bajwVCrhtrMmwquw+yMAQoiFNhfb0JhvC9mpRR/axTYKoAnJJJOhRqz/
zKiKZkYt1slg0pWLfrauxyLKXvFP85PJTf+FfIB1e/bYlff7gl5liffEEuWUOSruTtcGTbejzNs5
MWLJj408jgqZ1ME3Prf6Az+hbuSRP/erXLP4R7miuhBHJh76cchGQg2Smx7llvjM/0n0rXbF6mIE
r13JX2td1C5N78eoIz6Jh1v8DPsd65EiHAN+xWcbqCg8vEkSnlnO2dQR843CHX+tXdP+hLmzOeZW
2yc2+IhvZ51HsFijHngu55GqoaKqpVW0d57C+qLA0u0umsm/FG+VKMDu258/WY/vcScO4K2bft/h
eKXoaUVCLqfYUPfgNfVJiTVJqWWqsjRkCXKtuxhVAzfHUpkFZeCUvRJQBq2842G1CElndH8aJ4tw
kKgAemH0m9z5Oh0h8lMXn1ATkfMt0cBg2Q7aDJkLzScx0RHq4LRYGT2Y9FLcHCjp8RG+INMj5aiF
ZFVmHqoCFu9FG+tKEXp9h9ggUpKeQW55MbsLJAXpiCsXVoofjDL2lOaRbvXC6xAOwHaTxKIktduX
6RCG4lqdl/V01PLq7ZpoktTVuoydbAwn5lSpop1aAGqwDkncOHAcvxUEsqiRe8UC3w48OHIg7IbT
53XcHEukZqGqo86AqSdMiGVxYmOL7xkQ8Ht4MGgY0a6GMVmSXWMH6obvfDr4h+JwlIYaVTMsIywj
25qam0QF5EgajV5t+BJxNPJf9MAxEf+ZUjBNWVX+24xhEkLfEV+Q+GDH0mC9E6yDbBrCwRoJ81Tn
Ch7C06cgkW58se3O2NKciSaSrFt73ZDS+j9FsienJwYhAXcypqas6/AbA3415/9MZUCLCfu0QdSi
Ko2vKTmCB/yue0pqw3sUvT6gOwFgvTa5KLATFwQSy5tQoknXRyrp/C1rl/tn+6zPawQ6lJFEXv1K
4CGW88IET/d0OZWs/yO20MGN2JE9xFy1v4AD/PgcdlbdT83brIvdC/VNIxFxVMZPre1/jD8DnXwk
e3O4p/yr5HOQQgo0FTqu/mkESeYLy5a1X3ksAjmGl2GkOYLjHbdCBvQWJwMCTP/4cSuWdiSeXzN0
gEFapqHhyBEq6NapcmbI+3KtHw/SsRbJZDbbSu9xESKYFVI+0xu2A21IaPnK0Zt6fVokCdJX4Nuo
LAG77r6Uubu3IX/hjAIvENBP+ByNM5O42x/UrF7VSuoSmhbk3Ijkuhk0yBkYlseEnnkSjwD86hWz
6XmF+fxCNywQrFDbkJh2v12wwsvI4mfV4ga+RRccSdaS7PATUHpLswRM31SzbSJc2+0d6RSuzMUo
5qQO83jyMPKeWw+Vlnsx9uJqRT0dA+dUMDAqKWANxESZtGMdcpyjtIFoLmViE4NlrtoIMNJDkBa2
k5UYgL0eivVDZ37l+H+P+Gv2xoEZKPHeqajQYRa3Av/amDawDj+rzL1JmMeT/caNd8kkHjpkbSYr
KoIq8phpkkzCoJp8Dx6ssxC2PgSkEjvxtUu+h1jBlHOZAeSKqBb8McJYWZL6Pt3MLjlaSiVsy73L
79t2NGyeFtfAo+ucLYPgy8gTI3TA6xl55RwHT62eWSO8gnNBc+pVYkbBKZNkq7MmmoZ/ZCzfHZFG
ZfTr8WenvqoTdmJkG+3usymQNF8xd3YOVx8nV0zxPFhba29BbNHwURJXrdNQLUqWbNpMI6eFgcqH
yDe2X4Fd7Z7BADmme4jHf4PbzIFCIGt+s0cisDYkiIV80vX6g/31vp+FivYaMMgtm0MNXcDmEDk8
i8gZvUkWV+phTQAcLN3+KTFCIeG/EkBBEx3BHDS1/by00rxW74Rv/ae5wy8z+/xo+gi+WWVf7uze
FgHsPOIU6rXsjaIl5oTBAzIcmCsiyH4hef6/v8UJ/zfcc/orhtrq5AAbQky1Xr/6PvAYHGqq/1sP
N6nbwkWUMzheG+iE8lD9Iam3MpwcXHKlFr/XtCsVHchaPApR9qiUCLwPJqhfIbbmdeOAghnXfZF7
7OYICDVLy49aCEmOD/Y3lvXfKWPIDeWkD36mMNFJzQ5CEHtRPCc4YK61wFMjsftCU+wnJ6+KkmTT
nsRqAxNJZhQMq6xYbfYv1469WfvhPtqfEsgaIlz3LnPIi6yThY2T7Iq8f1Jv3j1LFcXCfmVHMQUz
2iDQebpouozkWNrYjgCuTuJXAwENwTf14vV9wojMeOB8AD1JbIZWtZDYGS6PHrDUpsy5Oigkn3sG
vmgn4PMYln/ljQUZMtP8ICLhwJst9UCKsxWF5Vjn9tAKQim9PWrnBatTSjcbShkqD3zCBoiCzfBP
5n+W806qc73sFqEF9wmks3eBMezZu4hVEWlBPFjNzkBQ2gxxBXaO+fxXberJTVWM676DMd6H1yBi
r+OYKv4dM5cy6cqP3iKk7JNoW2r8hqatUriTrMMn6ybtgzkV3iKkZ+qzNUw+SZNdalxFaXWxOybk
1zClXDaXEB4MTh2Vr8bWT+11tb6Dh3XTU4I/isqHwqfz6H+rrl+nxgRth+PBG2QIs4rSukm1twz5
Q2IGDruhgEDxq/3geOEc0lBD2TlZ6lbk2RSnkW75a8fh+KxocMim0oa0B37VNoZH1VqkbXIndWVn
ZVsT4Xw1v3YFP3CAlrt7Vk/E1EvDK1O06kNqrnSSAjiEYAu9615mLpAyzYzobt4fMO28Q20a9sH9
I68QQH9jH+fqy8J6nG+X+3OPg6Y0IN2DSxzhw9wkxen1ivNHvTF/30TL5LRx//TQEj9VBS0rz9DW
VEK2vjwFqNl6G+22xTCqqLIIj7rDgYS4kd8TJhLNj7PkSripkyhwlEQMmuhLcz6xn2yheEFXgQWO
ORmJy71Ek5Jr++x7ZYxrNZb4aRAJrqFudW2fp13M1EIW8BwnFmm2DhCcw5sDLpYsmnKR09GijMaJ
6goNzrZilB2o3lfU4wQC2V8ktrjBiDwAvJvFNkoLDAEXQMrmhTTho7CQ5sdR2jtyd3zzR2WbkvVb
xFKrbtMxHCCa/RrzFK0YjWi4gfmdwmmlsJ+9zlM5IrwxYhlzbAESQBgQdG4Km0PG6p6NKZV2ukhF
aeYSub5S+s9CpmkFY1AwfpSyvHcOr32EnNLrSNcrWkqSTzN2xHQwxdv3MwrmwkBJ4ErP/FKjEmR6
yYkyHr5gFlyOGuUpaGB4wSIdJNASZnvVzXCGOcuTpJtg2hFTXl2g3kt+5ZCSF3aPu+14VEySl7Eh
EUJxjPFoKqcct784FQk1WmF/hjOWu6WFLBL+qFwSY1AublqxBRVkwdKftFv9e0VBR52HUMm91xOI
EY6BVUYgEkUmZBjzwy+iy8CpgGGjQsOh3r0BZlmpYbKz+EX3iQMCm8i7SXrHo8tJX9GW/CPKL6Ky
YFlNUdjFhrdbesjnV7DaU/zR14JpeVCusiFNJtJMXDLHJ/m5WrW/1KIRYR0dI41qmnc6lhH6kAf+
DV+9bDn+50UPg+SJqlVKkeuKicFBCv8zfs60m1sM0TO80vn5RCtPVwaPepE42SegtWzhf93bIxqJ
zK7UKlBJYj6oSA+jAPg6qIj68XrNqmeTpltFXS0kYIzo4h0Ogu/hoAHUG5WKKwLQ05nNeO3rgdWu
ieY4fAVKBXHFdEY5Vlsa0Gq+VDFJ5ifmbGJOPaijOkXkHdcuVG1Akta4E1pKci6xlN/OiAwtgnGh
JNaSbmOpuPcbOcI8epEO8weX/jcUpIkp403ZzPJAZhrPD58j7/v1aK5bITw+c38kW3zfHWfTwc2P
tOUb0ObaFcPUm8m7Ak+enljcTPkdY5Vo6NuvvbLoNDKQ2Bm3kvE5Zrxk7itfnnarjkKe8zVO4bZx
x2M1Zgtg7LhKBoPRC1Yc4zdbWG/t4YoNgCEpw/eJH4igsq1rZoZdhhjFsySzkpsR6lRBw1WqxR4O
jr/90q5Pu1YGTx0Ig0arAJsEGy57MBoUrc48rfFS0HDQoBP8YPxW+V9o+dPc5816l5LogqV9irIM
LN3pPeusX8bGsOjjnhkQBRH6Mrz+BMtdfLmMiCDJvBLvRki9JRObLqQ7F6gticjjDAdOCmIT3R6J
y/ycXz9l3RsH/W6gfDz7iugm/TKU+mdcBSjtyAMZoXKVVu9bznOaIly/Lzy+JnXXUS2eTnctqYsh
D/UGsa2YUOa9Hnb1zqZFr8ur1DswnfpvlT86Y9KzTIH5X0e8RuJBVvrRSBSl62wYGoUY//oklL8R
hQL0nimPNpt83W6sDerEtEM6Q3oyK/iEEKZl5Hy8vR7s3RvlQA3+QVcHYqH1xDP2akA7pQHSCCZG
Hq9ANabJh1MZxhUQ8QcPXkHEeQbhvNUMU0enxLLjfLXVFjFFTO+Oj5lEeTED+H25Lymhg7pb3K7r
zSp1p9tMfAHSAjOtmden/jDM3+JNQ+43jnko1gFTLkV1qb1rlgOt9a44VrLY6filiyKBzk9UTVug
aC+WM/qVQQHB2q0DzcSJ4xDHCHL/6/XX18Du1V0OJJCMijU501elL0/NBvzsv9YclOkfZmcdang1
7t50dHoHEyQoABtj61WW9YTH6c5Mdg/oPp3xSVzyH6vBs+BO5IZfx7CyY+w/VsMvXsT550XNf+AL
i1JsfxhH8MS6zwSQS+aRUflIITLgfMPTHzFTcM8uBkuj04RxA8hs7IMpKyJby3MMtpik9PVBoDVm
aviaDEJ37DDh1Kfl8Owq17lSvj8cjJYo0utgUKBH5AY+4tOv/evu3dNbH84fDHulG2fwRlzKNofG
9NyDP2WmcDaHfoo0GM6fbh30scX+3EP1ThEUUiOEmVrRDZcBqaLe/be5csN8b5y5t0v2RHpG7X4o
t9gOG2sfeI+ruBoaXM7mxgJoNG0m10+rQm3qWVmXKLIkBNcee7K9PihXF1POit2sDoFBJhkXmFBp
Th5e52E2t4AkS0G5I3CmLh4blgKF1ZmK6eaZruWwqDrXOMDLGUz+iqgKTIdGySpqjxpZYsc4LmOa
0INzGE6F49RRddyZHGv4BsROuuk9bOzXk2w9RMrjsBFgBeot8yoKvmS4iyCtdc+mYJzXMse+TKi+
NEK/YfJ80OZKktkapzZlM6SQTMnjxAPgKSYXVF+B8tq60QUxOG+ZSgRP/aIbxWRl+T9MIUo/IND1
QM1znhouqeeXEciT+q8axlrYsfrHjPmlHF/Rc2GstJfqBduj2XBjbIrtKk29Q1ZsRoDfDMCuAgri
cCNQL2u9ArWsOLVkpXbV66vu0cRvOYlZTyJ5lInbde5b+tVQlpo+5GJVOm/afaGbj/Pov8J/pnnJ
7JdrDWY1InSub7DWByYOYiBGZyhb+wyYoN9gqLFNRxVsuXO3yWk3gGHvrRUjW1hFAyom5v6htdE0
hZlxuCFUF9/stx4tpgD3abXJmScO6Rxb8OvWk+xFJg0dieAFpEByU1vdJJjJOgWDTRgbUroejt2b
zHNubBNc0phNjUc2B/jtRLY5FXNUL1zzHqNYlPYhyJM2bO0P4Ra9wozIxyJmTjzYrYqEgzq48b+j
zJqvz1fDI6dbo20P/NxU3x30/Z59mNAIZElgQbe2t99q0SpJjtfm/yxQM5hnBBpCZLtl0RIwyU89
fgJ/owQOay2UKG7EfTDN+6QPI3DATVtR4fqUsKV3CbXer5FQyy2vBV88aRpMZMhhTUL0ik9pU/t1
JqoPmoSXRX7OBCAt51kwmh7LwmXSUiDFZ2urfFwFX95Q260+Gv+r2YkIxLvMfY24e0id8FLG24iP
cWQnmYmOxuedd1bmrrXdb5yXgzHIkDl7/EVdYB8yX4taw5Zz5WJSISVnCRvg149FDcSLppN3E33p
BEsgJzfhPNOqjRCtqN9k5gUkQ3v0zXj5V9XmeTxrzWeA3ROOIZ43HwkCWQ0mflJtBK+d14xRmfZJ
WWo8ywGtUHvc5m50tZgNEMknvuf38VfWc/goTpV/PfFp0Nt6l+2ItPme9nGLR0uBrIOEYMNaFc1K
hThUg5kydg7gaoa/D2UKU2HDlWB4OrwhO+r/79Pzkzjo0/uF3StJolC4MgBzHEqYaGVdY5c0in1b
yxewMVQNJ3XEYYg+emIueYEIc8Z5zgC6vzzlW7eINc67oe01uTchKtQpz4WCBFaB9Y9Mig/GCSam
iZeLryncvORdAxo5jryxfQJaQv7amP9PXgcWFqGm63QYmRnaUehAmyReZ0vNOzvWAwybKtf1seGa
+Ay3iTRcwEUjB3jO354aTC7Dg95GzAJnycHmLTtIjwnvtwssLsvtczhO8YsGjn6tlrSiIM+LXhDy
LnPXWs1kG8WuDIkMTMx2KQylP7X7w2NaVuuz6EatHpIWKGWahR71nZDUTHcmt9nhLOcmb0U2lIZy
qfme05I6ICtD1tkkWjJkQuAk8EjcRDWaOyAtEGi0eWIfiUJvBmk5NWqWBGvgoykzq9PSbnP/Ts4C
XuSKzPBstdWYWwTntA1E5pzbZEGOVgtVSJoAhHg7LOZJzUGrvmtSK/fOCM7nkX+NWXpq6BvgDvRF
uikcMT8AWfM7OvIB3Kdqvm6vSZ3swYQiDgdYtGx2vXsQ8HuY3AR8XaNn3H63vQJ1GF6eFfPh4CBW
FiX/lYDU+JupOgJ1xKlCcR1LaOclvs4psKu0H2y+TYTmWlx5meoZdYJX0I6WVxSA4YVGHIxr5CU1
oCrocwsO80CWV3RlYZaJrTkhkAylxpItnIRcrJAhBDKmnqDvLUIJ8u8qFPAEAcn592vU5GSnl/qe
DbV8c15qnuaTgoFDiAapKMDNdzJjqRXbuEvP1yjoFN2QWevj+oFehywBrS26epB6o9YIAXT4PnbA
ZNfIdn1cptWSh9/G2J9LrAXQGnUqx6T1uYZ/wilCVUCvRNcRJ20m0DTSdMfwAgqlaUbemm9UTJuA
k5LoWpBnNZZcODF8ViFyrA0HNvGmj5dE+d0VTD+69FWTfTjlPbpiAf6gtgWNWLCLS6r2bZtxbcKo
lHapfNR0/326xRI82g71SduHOdh5V82JUkRf/MN+ABcG88ItiamKP9WptTPpyFc6KcCMJzQVAfMP
mTE+3r+pK3UCKz+mZ/ZsXHIPRvjbtmmWRSkZ0u5dHTXV6bLKO7V1BrxkV9FLr2seQfjg7dS4g9CG
bjecuSi36axtuh/i4YRLvefb628YGneFsecDtikM1X90g0cf4MEXv6P3o+7HJ4iqfHBfxq32o/+Z
WQMaD0YfQrtI/GrrbD6B2/XQYuHHdA5dyeFHGXCX2/D8R8WZfVMQQ95TL3d1H5YbTnkRnXjFYwVq
eck/415DgDdLVu1dv62CbGn9IUE7WykSAdtjDoMpryHD+gOekHfWoDixEXNRfIcPRY+Jq5vibAAE
FhEzYsd2KgRTOaZr2gIun2YaDT2A/J2ssuC50TOOZAzxCrhBasXM28IA4nxI9vTe9sxTdwPbgxzq
1MNRgrARBhU1YyFInoDRg6q+6woBBMCg2rjg5O9vrweacctlOgl6aIJK1TcNm+MFWBQlm61Rq7A0
bNP34dLlw9ZQ3yqehG9cEAgeTnkuzXoi3tWK1QQtWwY6hZTQCO3NHSg6ckM14yob4hoIKmIi/3Rn
7ztTxlkKs4E3p2tpwzD9mrCrx2ta572AUjTAHbR4GX9SX9ALH8ZQlDJxRbzaOjuindvlv4EpH2eI
ncVoD9wFqvZ3mjtbLNMaoBLIOpUnzihQouomh7adR6x5hDtE1wsOVyDsdFBkJnzqc64cbfWQpZTq
aMsjGydbd5mqHbCVqM32WvZGo6LMafflQd///LnXKJWiQiXj46HFPgFjNV1J8suLB6VlTrH4f8Jk
1y7qSl0euX9uBRN/wJXnIRzZvFNCZqOsYcwUHpioQMNUAD84gfinF/BxmcZg5V0zdiJwUhzz5n7c
tR/yRe/ewQeSXv34PXWOuMJfyJ+8lLkNY9RVjohNzZcGFz7yLcUtS+cgjxulY7RxisZF+uWdIodT
9a7VbQ47h6Bav7sqLjVyD9/6PUQEJXKxI50FVaohB7gRTd16VMj9as5rNWB3n7KmJHOVRTQ/EaXg
NGOOWi+y11G43/brTAnwl/sfiHnnaB4eufKukYeESfLV0xSSZip3WYwkIhi69smzYFtrS/X2jrk4
sf1JZtioqU+AFuNHjULSwk6bkvFbc24BmAxLWhF1p2fEZjRAUAlQVIEce1p30Xqmlw4zO8TTh5Qn
ZjkXv/JVIIVtzQiPGkZVdWPIJfBWAUPHHH+39VCS7tPULpKEFjxZI7EN4NMi8fKfDbCsHdJVjO85
afcGV4l/gxIZwPOwbLB1VjESBEzk6pdS+sbW1Iw31BOo63Yz344fB+92mQ8ydmO/GDuSK/7t3L21
to0OE2zCMFJdoVwOU+pF7aKAscULptOEAXbWo50GqeI5bX1xubQmBM7LdSuMK/yU39a00Smt8v0B
WaLjlthXEJvxRDHWmsNxzUgVah1dejc61/fyZcORiGdNTCEI47lebQVuE0wWKfw40dHpxH9+hhHk
N5b3z8J8R6w3DLtI8xKv3KXvHqX+t5OUCCRWLNFMyiCYPlOv1i09824GNVajGzC2KOD8TRZNqbCZ
aZWzhZnnysiDj3n0wAytM9QTHIvA/Zp33Ob9MSVfMNq1yyYAPJEbvJJ/Bx8vIdbosCv1TYMxAMah
H4CZ9UTdVTtDKuV1zxcxaXeMSHtbWfruBlFJE3IMiFlWJZm8ORbloOfY6LBp0TOyckreDrYYhp3K
aJ+RooF7oPbeUQzUPUcJJPWcwlY/Z+kacjyT+NVGWQWjBBvyusj320RG/kgY3xb82UxUnYn76A4G
cjIlY13oYwuP9+cWCC1PbSLJBC2W3RfbysihDlHWLBq5Kn+a2c6Ic4P32Vm4ys+MkR45VxTSD60E
JYofQG75Gun9QcVY3TdKti67n4ngPU6mEab6EmoFsApm0ne8TmL8Y0kLgIe0vaXLPWxBn3xIs37I
YmJazER4eXV0i7ouacCjz16ttZ8E5GHLVcMYujmvkoySt6Txid3GPwxFMnQVKRy4i3nwpwAh+bSl
uuS1z1OO21Af0+kesO7hOnugd/xwEinI2g8pQuON5UsPIe/5zhmLCqw+tCUoaSI6J5H9SItV+Ptu
ZyCWmtYL/hbq+Up6mfld7G8ZYcmrXAeaQ/TJ6cXtaZRTeBNirC7wVaGVJrnFO+VTJfMmWcn/L1Cw
ROiAtVVOkjnv9nAXfYTDE2PzId01FyA26w7t5Xr88bigSs9iEAMpqm/qVjzm8RT88OkWI+rXJIie
6Aiur6jzvFIQ2Yl/RZby3KAa/e3F/j93cyP0/EsRKUH2ugo54jBRKQfkO8IT0v+Miw1GbtorMFkG
5MMwHL0y0Va0XpB+PZBCwZ002YJCpbVsNe/MWQEx4exknUlqpgUVspf42blsaGnu9nhtNGRaE4rR
Z4U5Gsp3yt5BaR3oR36qO/qiHt5TOL+miMRECVb+cgvrPjYxqJqf8gi+2eERTcVOAaVdbMR37NYL
C3fL409WDrL66zwJK7oJvu9E1+Bc5olOLLO6QsJMAG87OU1RFftanfEHVLqBKqeYoaRER77MbPVH
Smt66v1LG/h/rOCNR5j9j9RRwOI3sA0cpG1dkRUnyt5qBGXmsf5vtAlfivABhnDQ5lK+6tNjrJpz
WGYB1hZ2KuQ1sABl8LiFWvjxylUC/eglzjDpUd6KoVCxwQgjhH+2/QeK8yNGYBvKKdGtOioQeZOq
owuuwTmPlQPbeSF1sMBbtnWaBPIRxr48M9a5S4Tek/Kf/R6r4sTwh2UpdGaJ7qFXQeON9WEclTlx
hgZvOlw3qU0hO8l46X9DwZM0z/d4qjuWxYrCA1vp6o3Y83B3eqWJWklUW7EiwT6I8lIyUFW9QcQK
xxdYmum+f83Kpdce9iOYC3bRPLXAuiJqeC0wgxjHfoGhipbwUbfFeD/nqwUmJy1Dy93W9hUs5oMA
nWJA7BVQtiujodSKSwrSelF+YauDKhBSJZK1NUJnj5nWeXF6q4qZZblGh6kYZknLowyDMfa3xipN
H2RGp0F32Zb7ZTHTlzW/0nhlr0I3jcKkYVTkYyMNbm9VGPTQEV2N7IkWVhr/6VIiKoNJ9AeQXtHU
/Y7JC4UXFkPV7hi7cN0Mk1dIPSsjtD3Wve5jE9LtFHBNpJgZ4t4OKMcx9K3aBlG1O35ZtYoX4uAF
aaLKuAH8GMyv31K4Xi/TL3BJ9/hFCkA+qXr73jeLqNEZIsbbwhGskKrgQgsPOe5X5eWsCag8iSL6
ZsjQCJANyVhTf58x2ZubJ+SmiM449T6PA864xWQ1X9LzEQG2/8OYf6C1SQwax2QiKAgp/gz9pDu7
26DdqmIVC/mLwQLhx3F8xX9kD3Z3LDYpY9hThjyCQRA+eutjKbAuA7W3/PdpM85IUosKyEAs2tmX
eCgnOD0kDnidMn4SlRbNvJzziMdqIMRtZwDDKXXHkSzQsWJq2VG8YGSD164eS+Uwt03hhUI6rNGc
n4HrnKkZjT1eQMU1LvtcTBjfoynS4d/Y8tTdC+V3GnF5zoHHF60qsyFbT+OyD8kTBm5ALooFuA39
8miTXjanXhPlDDXzQG4FlHd4bOVsPqomztC7rCjNbZHM/kv0jnEgPqRCFqFK2UDqz9ZmnixGp3CY
1+eTvEwTQgN1lIoSGonIrzZ0qzqJU3+ey8i3eu26KgKmD4z4m1rvf0qX0TwvdTNvi4I7u+Mabd+p
28Tm9sNntuSQfOjavdif4f6LJXgSnnwnbVs+SRLdng/vhhQsYPnKLxDXkSPvjVbh5KP8q0QD1WkG
WFkPHTWLTEEob2Lx2xUqsehpMVXsLP1TZJw6Y4csnpOvJqqFDkm3fystlSUDrtuhAJBdlrKEl2H8
SXSVS5kGFFMKsFGrUTG1iFvFZ6fmstKO4jCvK0a9c4AClcj1VGp06Fkop4AOuOxz3U9LqZ/M4I4W
c6Fl6FBjY+cJgJV8/4HU9qLyASEhPurlfNpWaZmPGsGObbx4Axr8MMogWYp5NWtatXKU3KWotOmC
oBvNghKwDSUVRD9K7IOas/Yl+Q7vhXKCQfekJzyaZ2iHkUmPobdL/Ij7bas08gKY0c6KOnoX5yX0
Hc4020kehsb2GZjKj3vsPVQr2S212TpeuRrvWGELm7XbPHK+pJu27q4J9dW/UtJjvm8JG1xwa98g
of5u0oyPeEb2vShaQWqIsL+cAbPsTmr5felPK6rPrX3EF1/sqkEdCi6Ml6K1Z9QeKdiYXNCQpF4I
qLMbvsJVelSgl3adxOrGgjTbnjMRqBu/mXmIT8e1EYikJmf/aMW2xxoV9EmjqJ2oIefeKFOkeTur
aic9o7jfOLj/exz6nD+i0yKBD/uS8UFfCq9RefINAI4MzNmgjKOsy0BqoMmhxQEncjSnW6tIyrNV
+qV3NB27yTMxQQZLNxmVbo7UXrUZBb7hnQjkdg4YkvDne8IUzJP4X629yE9xzATQ8KQi8boqv/uj
8ZOoC7v5VAUHfrHc0mNfKvjlt9jKqrHO3PFj6P9i+sv0Dtb8WT02FSF53Y91NtTVvDTFurGAoruf
ixaOjvELmd80gPGIVp48iwCtLNJPs9se6+4u7NZKf5hsKTx7JG7O1Y72YUe44eqmlqjNEW8uwbht
LM/ALo8eN937tkvKBFpofq5K95XHO3hEzIjfUWiSOarl/nHRhmqzxIvaW3dfbN4A50G4Tv38JqN+
unhNHSx8uMRswuD/hltAOZipJ+VlyU52QnK7uVAzZ18EBC/dV93OnfnmxyhqDW3ifn7mVoEfU4pl
/aW+I+teQsMMXqrKHmGZiMn8fH6DOTgf/Bb1gYLvP8oLASESkjrmnDionxOUtYopZlnNgHpOB1So
xFQa5PLhgXIWJvyxDudfWOsJtVO5qd49zK10RUjCqLoA/GTG4cEdCIcP6GbSLL8u3nvkcdnchfX/
W3k1xZYWok4udLKALGNkIUbKWxYlJam2LiF/L2M7zYOz1CRfcKfkIadzXKOx0o0hW6w+6qvFqgiV
CueFVOLHB5Iop+siN4elK1gUQAJ7NNCOcBiA9IfCp4j1YAm9mJs3aoC/2cGDCHfD6+u9n7Q/nfjt
fsS3SsqgQdAbH1U9MIhViB7f8dEiifNDtJwpwByaUE39oMTMamm6JpdDbqk0qGDVMoD9OsT+b/MK
dQeIUwtpHVu2d6HxYCpg6lm/xB0X4QMWXrhkx2i7d2y869B+zVFQTAG5yD2zw/FpvRMjBBRJJ4z+
cst8KFT3mjYMugaMp8pMAnnRxyhW44rynxuF3DONOLZWmcdTOQb/mhopyhPlB5ZPvcruGS9LeSP6
X+Z2jMn82qu/n+LvmOMFfRdjEWvVoXvk+xiqkJ092yUm7Zw3QDg1+34mpLSQ5Fx/zQ5iMUt8Kah/
i46lAty0GM2SRd+F2wfupYDQ71mAvLpIQUtOBzSHFtAzhq9c6RjWZL2rtdlI4Z2/BOS6/y5Pq8gN
QMhUmVTsDpEVrdqjSd7seqx/mvazXJ5+v/N4xYfeMdYvm0jnM1NG8cjXKH3vb+4FEbQDtygnXr9u
5NnO9T7ru1xD+kPAafRJ50J8//aot/eNoaryBcEqfqXBBTtxzwRkenqGxtisjJeA/VmAu3eRDDIO
yHizSYu8t6ru2iH46XKAN31da1s+mb76OwdLibCrTM0pbc8YprfHHfih8sH4oblkn37ivMAoHg3S
e76ugqdLw8AB/l663TbjpLfrOKytxOBpbNBhdSF9fDdPmqmoXdS3fuqBSQK2TVglAl/RnWK1Ch5J
SxMwQwETsbe/iPwa4df/hGiD7FVQtzzuwNcqZVWqmfk2DsamMfPUKNq7A2V96EqDT95haKqh6ol4
rL1aEL8NbUwxNIOzYmiKC0A8mUkryQKjNyPnPUQwkZdMJFGmN15ZAel1WJI23ELHmDeSbWWdh/pT
yQCfW2pJF+TjIsZpryI2+yWcYkuUO4PYMTHmQsiRiHbAILC35lYml+vUMJFl8pvFtLxDixOzdxvT
OhegWzbALdsdl+Aznt827L9reRz78Xt0lqzFey2+R/C8ycblYABz3Pyr4ICVRlfnWZy1SW7WVuyq
ecEY21U5z5vUMv34VcXpSkjlnt5raKo2142Wbg3muZ+UXec47xGN5eMiDmXqu8TcLJxhD0UxTLlV
uBcikWaHniCycYb7/PrvlvrWttgb31KThsm1J9nbgYbM8VOkqQQB2pmW64iXxrJmzrr7m7sb8E7e
0qz6kJtUhKITBQJ28SDNFrPQJvHBlKjFIx85PKiSFzZuvcZiJGjabu5BcT1eG2g+hWzJhFtUGrfu
1Ao8dHYIg0zM7kUdPEaFlyoVE+NDra6j9qk4KAN/Vb3AcwyVCDAA9zujpWq1QmQy410sGsQZ5C2H
Fede4bIAkCvEeADQyuRBB0tb222/CxVRtIwMUs2GcdimM5MavOFkdpyOZA+ZesOFR2FXLErtEXS5
ZED3n/hf/WWsSRXIvLMTeqKJ3uOY5MoxkpO9BVorZWjlcs651OgRzTbiM3UC0RFAl4DHXGKDDLQ+
GzomAXvpZnu6B3tEAvMq2eooP937nZhj/svUh/Gjzo51n2UDHLcCf24ceuKuVSea9iDPga1ORhBU
ihHB5DUbZSt9k/2OYINm5PiypdE0Hasii6mCD3DTEAK9vuGFJ673PPvD7EKUxybg4rpDu7TM2GZf
Ky/TehEKmBaV2bgyJEMMokCJZT2CH3Nbl7PuQLb71u439gC6NTv82+is8GEhb98ATKOgFRegBI5N
7SiSwM5sP74H8XAnKaqcFUdy4MnqlmPiBQxJTf6gbOKtPhQx9RyXh+R1thkPPGdbxqPYXI3sMEVd
MceQl32CVHkz8FbUnTr/htmTg41OV0CNc936mrYnmFrWsg/xuncn5CScTmg97XUnELmgtAw/U1UJ
ckULfDHVLi9w8D4P8ohLhxdt7kltOUkbI5QX+zrh93YfeNy5uoTUA9kaD/1AUZ3ekNvqHkXOtdsh
zp/u9VPfNUGuO2eVuRXN2556glXW9tiTN1PO2IVk2KkRjXExIAumk7x4pemLzHS2+n/Sv22lRX0G
mVE5iw10MI9v3aEhV8fbiDKPiBhKIvgaXzvkuRugjOQJ416JP8kagEIBMY9Wm2wfPAE2tZ9cMG2G
vWfTqiYxLft16FGFOFGPWjTlLe84MUAwo/GoXhnOfR+2jnqnu2m0POJk2VP4gtMn/odhyMIn9mPC
SocLkgVP5VkOE04PeTUf7n04NoTy3U9rCwaxacb6A7gKtroG8PayeWWU2bRc5LfXMge+PzUvd07J
xgIdVa2sXDd8YgHBuYzLwbgpSx5C6uMS+Oa1wVmN5Zfw6mDfZGx8HUojLpFKlcRd4+hzzlwGFpqJ
b5RHE+9xTxOk9T5Z/sbv6BjQapC5qg76KTFad52Rsd9GWsNgy3R9SSBQa/Bp3O5NoLDz244FFhyO
9V0+fZwAkV2M9OXKKoAiYB03We6QCr4Cq8WxXnb+cUcEgVbAPgKFOeHWa5mNM92ymX49VMCRvOyr
umPkykITkPyg1zv6cg/ej4idvmREuFrUsL79JUmoYPG3AxyKX1lEGGSN80KM62DuWccwLlRLWcLc
+qFcMd+l0g4Oc9baFArSElcrnHZ/Z716VYvqiQopE9MN7ZkExHMWKm2v3w0/QrFSYa8hdTXAi3V0
is3WbkHbc5bNsirxg40KfSRUKhR7Z0GSFIsWwXjVTR/bEdWYTE7xg4zezcWEkx7RWJ7vkoGttgk7
dUK2j2cvoR6YTXeSP6DXaOVVNPVKov0ElTOX638hWVX8njGeFRQpb2NsDFXW61ajGCXZFAWEV+y0
O/ikJfi6Ayqe5wZ4sm/GvBPiJnwn77lEVNsxX1XAgTYxIVjGyJxrW916+O7e7vO/1rqRJFI8mbDz
t6tdFFNqEjRVaUW4VjJr7785CHznSXjmvg3gADdfGhrZ9JEDLmARWXj260HOtC1l2IXy3lp3QSvs
bfP8ksHmkRiBGri53LCgnARR8u9LD48TfyR+h2maRLYIsLRg5WBu2NgHDWJ/JZkG1V8PKtfZs0Hm
98I9+44I2+sGJ5YKZ7OXc4XLE+ap8oPy/kyPSd4XuLzi0yCphU981ppSYsn60lgbAGnQ0uPRHLuM
99bv5OI2SgPpPaROhiJN+6Jko9vG+auIeU1TdiI42/yuEmylyiluVynqr+gNlFI1I1cg1MlSJGwD
JRI/+j/Re9TTv2Q5c43Skewy/vt5NkqM+AtG1tXUFkLVPFz6xQaE/A8bWVe4RnVOjFlSMUAt8+FZ
djyzPXRVnRRqoU1QVsDXqKuFhSKIuXrA87r68tyAxVtnHn8sKFPir/LIexQd1l8AA8h98HmJmjBs
teN6HBC7FXkortcIECqfJq6mHEoIOZHSxwtaGkHOtnAmai6URh5qz7BPH5sHwBUGyCV3QAE+iL9K
lmq566u6Vh/W0OrCHI4pQRnHmaSfyF3u6E4RkkexezctxuZMP8J4c6uAJ83lW7opoJNKH8qjCZTq
0XA1H3Jmq2aUxjJdFll2omFdiWLa3h8aPnHXZrnv4a1XgWGggEkxzAis7Bh2v2mfBr/YfVLhZSKn
uX/+f6B7Pzl2Ovb+Dd+ttt7DhZuj5j3aLMECf4urVQvyoAPlKH9PXSZEOXhhpHeMd5NYGCyeSRAd
dutg3JLGmvjfrewD90H3zW6eB3KMme10vPlDoPWHZdGkiZTThht1rm+7s+L5udfk3mFkHoNe616j
XX493bw/u99jO0EACNfBNlDaigzc/ef4Xq+x91N1MUfWafDrTkK4wK7aXpo6qjuK8qoAdnWRlnYU
DCtPqDvoMC7sfO1Apnf9mNinjI+j1SNvrTVQ+j9T/IpgA+ludl5aTYcFe1u1yQacrNso3GYCkCOB
wznu4AEv1CH83nj4Hw/u2+d6L7PeUiMJ7K8OZU27D8YMm6eU58DoC7qYqJeIWzPk/64A+Frxmq8V
ofBgsh8E2AX862OVuOrI/TgeoB3T6++gQEKLqa/7ZRcPtlNl7lWBmsXyEkpAHR8z4WyVwkHIXuPK
QZtwUbkLjU4aTF7nGKB5fi8nfesq18YepWqp78CssYlPd0bLw3OjZ8KNKVjyoeVZsnQwljpO3mpM
CS1GeobX6HFzt0qX1++xBD0JxQfOdtMD8mTDWx51MYE4wJ0ZsgoXn900sODcu2CTzEKvdYVDQMIE
1WZAu+qKEuu24kB9fFbwcFgihq66bb0R7OkwII1r4M5Tq9cNli+T5Nji0Kc3qtr7QBRj1Jqi4gEJ
YPuBSE2C1YnG1pmeDH8bx5vc+pKDyJd0gxEsrok1GoKpn1JAPB3t5qV6ICrADK3/0pZxvpHtr1vj
zKLs4ATsjuv9e1NlT1j7KoJyDxQR85HBYFTKcbo7QtmSlKRLNK3P+o4tLnpsSS8xy+KpsHnSI+0u
OsxNx/pWHtKl9bTgGvzUDahZqgjy32rp6AW1BoSk0K2YIqQjsQ3fU5FskGsJP7/aVOSWYOSifke5
AygO7YLZ20k8c+czW047l2qhcmAujauj/wc7E+pMhP0I6k635vq0f9AKz/7JnUfXTJneenFqudHe
DVKeb2VjNFhhWENIxXDcSwZr0FpuV8ZSRRwI4eBXy/+7VdrWFufU3ZROwt/X5mgxdNW1klbCZKD7
uiz2sdM7dXOME8po4PZFNvNo9U8Wcg5Y351Uk1ZRHwbDd1NUS+KIyYZiUhPlS0JSiVPVRc6pmEcV
Kj0/Qc0e0Ebw41eM76MHDp6ONz6inxCrrqOqXWhWE0dDi1zaXl43WtFro0qcvY5ESPpKsDwF0pws
MsmI7ZzV6gcbODD5AeIJldNOZUltXSG9AiL5rpFQ8nJMj0X2WKX33uN5z8ryKjG+pbEeQFrhKf2r
DvLNFhZwboTSYdQJEj9N0kFYeATNYzPw9kE7N8rFlV3x12wTYIioPZxYjYGfvREdolOn2oG2dgjB
mxgu2jyrb9qnESMmKytwj+d6vgHy+VBX1gd3gTG9iAqlPQTVRaUsq/auGl+AQkDJHsTCiKGPd1UP
F0oo9w4GsP+3cDgBecKh9gJFVqhU0MED8aStSxsjXzVr6ZltQxKN/oIa1/Rzev3f0M4iPm/8h053
KdR+xBhtD6UPLrhtFlzk85ZB67QCFT1zrjHrqrpZCu5/tKQ9qv0IzKP8E/MFyrgpNHHZwp0q+3av
nRIgiHCgI/kYOowKK3M9vdK5rcdHzAuFLjeZJPT6dsr0Ab4zqzddJPegXOxSRCSY3vxUS46Q257Y
jylXJabsJh5KOwsKBeNr6DNpfhYZlPFbQ0EDkjVpWkehY+4Z0v6+fgFVc80FqBnB6g23JSCyAaCS
whmcMLaB+DxD6U1rsOjKV7aT9xCpPrCtu0UDwOSZCT6Dio1S+GHaOTDd84+wjkaCbV4/HIrfHrfk
MnmxHOzDg1NNIBYa2VbmHtxgdALnmzB3jFXb+fy7RF60lYvYrFOwdFxHFLn+OgV9yP8/yIBbmtDv
jwmYLoNycr86BzskMknM5wLV4Xcrxo6wTVCGgthQL1upvt2GzJmd8bkgZP+acV022J7Jq4ky7lz0
CNRH2SwZ1PYiArsSkSQuM1oYbL2znMF30H3/sBDMJDoj/eKgt6mCMYSlIEblVVhUaa/hwMqeY1jM
Yjk6xNq6i2/EG3rEZmRy1riwVBvg5UH8yL0p6kO0wVj3UBXP7Sz+nDUpHn3T83WcvnWripiP39Sk
wLjnyxx5+Tq0C88z09fseLJy41ZysIppjqtmQlgIIc0IrHw50HRYHXOvPxnby74mK5PZKMz/Z2lm
aVb7A4CE4ZQw526fBp50VmiibjMPKl/Y1Dpq1oIaX7iL1tNHmBtwoEWTWmlvpJRD8mQdGEDgGuW5
++0aD18BuBFGVvpyX3NWG2Zp3aqXybXif1EMojpTgkFL88ydoyMeMO581umiuX5ue+IdeE/Uxbfm
ujSuRIv3kObcYEKtNK9zSZNAN50WgpCoiqbjLdjMdKT+6Pu4K3DZ1qw1LX95ydRoxoiMoPnzILvr
24Wjb9B/vjKvT8nsl91HdIRoa5qgKqaFGqFAvryLdhipo6ZwvthZ/MwxYfhpFoMhxFoqrOEO56am
kwYKle538o89ivDhW/jPrdKxa6qv77oPE44uQwPcvSuEvGb3OYaVCpiGOy/Yvl9mHNEjkEEXOREb
oUmtORgfOTqGghTHTQJoILMF68CePssD5NPQy/0Zka7qigLtiyVdT1qXoZbKpQLe6c9YLk5a8w4d
FOpyNp+qcw5Oyp/McZkDNUk5PtPBi8JBF3IL0OWq49f4gFD9WOWKWMA+LkA7/g9m48zP/Dkw8CZa
/r22MasZ7aUJjUgWyuoxIJ8hMfY6jItj8ZXeZ3hnxqtcFTx+vL+VW1jEwxP7lWFBDRdIbLdzny0M
IO/gMDhS2kLjFWxemGy28qND2jTZ66Fxi6w4B9MhIZSUlr3HfXzINnEIxDopFK3CAax2zYRLhHJX
JX9Zeo5iD8PBTZJIpUYvb+XyXleIBkY9znXoy/KuqcgWgJ+tZOf2QNNWrVK274piVy+x0S3/8S5n
iP4Wrstl5Wr1RowEamsFAW4asIGZ0/is4COCj8OY9N7Ic4wMdl941rwQdvXzQ++KeyjCWM5lkBgJ
fdx1nx7N+9a4ybU/eRZX8g+aiJ4CZEx2L4ZSF1eiLd+8iHqsnC7R9xZhFQfyv2ExNsQ9MCiH53F6
/3gQ5CYu7isjDakP+DhGH67YstHu86mgTxYQ4bTS4bkmfY2EC10L4nBb7mjIJgCfhgw/y2x7gwXN
gXfOyb2AH8ChP7QAcSQRnI95/V0WnEgL6t7awn2PdhV/59GUqKdvGgt4hUHHD9u3iiZX3ODHbHtF
ERypXgJ7bgvUPqgh+riDN5lhvmPJbJzSQAOyeh3oHGizrSp3E/55O9w9k+glhjrO4xH8yfnT3zcc
1/iBGKk7E/PO0HbXpgcw/SRNFk2pYpisW0y4NK4mc5FleEFVRN65srAJhGcLrSqCe5buoaRaa7Mv
aY3Ai7wtv+rEd+P+U7Zs8V9CtpLVYhhYd6w2Ts6QCwO0eqoD1I6xdnJGD5oJdTIRJ8/BwS0TtyY1
JcLASJH9zuSoqy9G6nvNndQphwUGkm68gnAv4GDB7Q/V/h+491BaWzp4vwWJ2RY6flaY38Y5TDS5
qFPMFg/VhzQ95HvO/pyQbqWt3jRvSLi1hYSCu6cCA07FbSZZU0TnIbAgmmz+BEZ7DUppSYk1mWp8
srcYODoqsMwA+0q5Ewxy8Aew6joGxR5rXgSGNNPckJSPYwgYEmgI17W+1hQimWD5wLUM4hCRy9pn
vV637j+HZmYZtF7j8ZC2ibmmFecEMxJSDYzijwtu0dNkzXtyFgbahdHNdcoGTehbHwaQqYKuYucp
876f7ZlJodxfHUEPArUuKZCEtWdkoOz0zjVOOPwJHM3PENkjlOWwGvO2CP1ymaOPHN9vMnpkBCBb
qsdufh9CF4zv0Lpt3N2zQ1l7bzuYqg70yRXPSilvsG+8YpJVMTiIGZNyUVEodyckepIybe7MgWWB
yhdbz1dHQMgBxHnkXntsNWE7pgkvpD3qjjzaFU9bc8RGs2zwnNT2z3J9uGdy2XaWXE8XgWnqTMZ5
kLjbp0gmj55JGH62dStQaXIitT1Et4wlOp9lLiVnk6iY86QWxmxwuWVBuHyplSLZjQM45zYQYUHc
3ETs6BbBhpEwII8y3VJOH3BnFmaIUt6XObqIh0u3ikE4P4LK3btdAislv/tTC4JDPqXtY3YUpe+3
9F/qhTSJpp9t4t+DeO7aGhiPTHi1907Wmcl/ozFjtWuBsZV9Xd0MWnjN8BV+X0bNLQ7bTjmDDXmK
V1J6Tr7fnP76OIhOKtWAV2SsVv2EwbkoRwaKEr0g4Msn8Hb1uGumsa16DZJ74GnOBSKuQqJkQcKn
CBrxJkqo0uQaKaBWBsNebPIY7JBxNHp8cPBnNAC+iaF2A5UAaYjskWmcUePby1wgRWIO3MlGkCfP
972PlDsoxw990BDL9ACxMsUBEzwt1I0O2az/S98r/ysLlxAeQ8Y/zC78sRbr4exAodIQknCbTbNO
vOTRTYNKT2TxKuBpEchPQAYLW61vmJdfYHv/mbKm3AAyCuuNp9QHkrnk3HUt/sDN70hKvHQ+W9Zq
8hWBkP2YbElUABRR5fKWNUsbw+M9GDL84QA5YSSXo9qG6zXm+8LFRkIIaIiEGeIkmNA+XAT+myz2
XhbaoOzui9g/H8vxFALZHnl8rTuX+GlC96wBXEJYpdK1bCsDEdtdYppIz4xXQH3D95CfN8MKPZzc
0wu696V02S8EM9haBxvjX3ELw8BNEXUr94g+c359eQ+ky5NY/b7GbUq5b4U1sPtIj1Yo7NoN9cd9
dgOIeUPfPkzQ0c+3DgaVJD/pd3AsdudpfpBA8tpoHmN7plGPYZmKSt9NSDl+ev5uvD82V0G6OD0W
e456hEoqBwuycl37KGkrCWfrwVi2hWDUjuVJxBW0+wu/coHQdR+j8dFCMdgy15gBL4E/IQHR1kmq
vJEe8b4SpZyJZIbaqyfoKBviIpMP6J3yy3QA6FjZ74MsSYfE4YSJTSZqEWCAxYS5lAlRwNln/FsR
n4pD3Sc35NftPx9c03h8vWTSgcW2YYHnsb9bbsgrb3XaSZoQ9jeDagNosb9nL42y3Qly/0zmzCbn
FcIk8kctbD+zalHgLQW0Yl8580obfE/bMhL+1mgU5Xkpq6gEnoDdb6AT8zj4Ip2alkYA0ikmGZ+f
UFvkqGmFTiOgE8mbYSSVchArnvyO0VDGjDXlp7AGV3oarRyJRHPPLNOYVDi0KkMfP83UIjajpFGh
gUkEDlxEHqqtQLGzZ9usPRU5kxtayiGyqmFpEHgq43530rjcOC5/S2+YSeDlbqyo4Bmt4MzwdzYX
5gkM66XJZ7PjcQ0Jysej9D1jsXY0lBYsHu9D/czXsx8H2umRyQIvWM18D3MYgBB2D/K9uTE2kFO7
KSa8M6ZBUeEQe3ixjofDvDhs3EYIThl0fUe7f8S7ScAxoLwqiXBVKd5lOqHIPCqwUS73oT8IR4Pq
ni9p8S5tQwZS0n4Lq73jITAyMVIkGU5SX1lR46NWQFxhptvai7SS4MBfwZWlKbM7mM+2nrY1Iexp
t5e7IPGaYk1apAvXEQKjpHC419ePclh3qg4HTpM4OsBc+MVIv6eAhvIkgWAflKZqq/Jwr4iwVdEd
iUddVQx6dlf8JLaLqMpyeOcsHzS8E53Z7H6HNu8Z/pqJ5w2BeD+H79tCviTA7H75IfB0WC5vQeBi
lYwy0C6O+utac0cgRBDtW4wLhPwKeUte5+oYJeV+kky3PCSuf28/Y9BDR9YOm8hokBsiNpEXh8jw
ma8szF4x7JZy2Tl8uES2RqaIuB8tFK+kYt98k/KE/KRPX7x+5VMbIB+3B5Wn6Mgw0uZQZ/c7fi9Q
Sse9JIu5ygjqqnQjV8BjxS2a4dCY5qUCd0BLkjzN6aGtbBUhTiza7Kgb4PtpkuN979gLXj2WLHwb
CA/Z6+9ok3cddDIdTaKuYLxjJy2ZIRRTXFzN55klgny2i4+qNsqkJasHHKWfMDezuTJwlnnjCRSN
KQben57b2zLIXLSPqrvB3axfBQDartVw5NPAUaGczTHj1+QuFmLR5IJq5ANz6SwxEx0IUaOhxLSQ
DsQjLahTCK6aLxePcGqsWnSHkWieoO0sy72QIfsS++F4morKfTRSN7xR79NM4QKJV3ZEmIoX4cVT
/gH+s+covHALtdMbhlZia1WOc2WZU1jp3LTNiqJ4ZyROp6fVV9jq6hC1J7H07F0/cYSiwmP549Xc
KdmukWyFjIFrDTS5stgKRY1t/O0Ckdg1mvNV1pKpL5+bYNIeqKuif8VlskVU8wnjFBpK8+sAMakg
Gy5JkF8xZk+mMk8ZjYMgtenKbOXSluOUnRPZcjH3AwoAgv8WuHv5b20mcRAaBGxEjgKIQ4CaOASn
nvnS/vKWiQZTZZobS8fC5Im6w+0NCqWbRyJ7ACKbsOn3yITHCwXGnlHb7E/hwZdr2+XuCQqt9oDx
MdFouFQWSdtlgvv4qbNs1CMJS43BKOuj5YGug5y3W/4Yb/kQr9jWRZciMjDZwGjL8BFNXjkUPqoE
Vomjr5jV9hdUZgAYEMt+ueGhQoEbAPTMifgJJusG99RmYZCs9tFDOn5oaX0tt4wSzLbS1yT+Qyuw
zz2Xsel/dKPKpdPH9hcHAQzSp+9hzKgG11QPyao2MEshVwaI4CwULfVNOiqy+f0BOqRfOcBsbXPb
/f8CmGt5YfzeTtsvq99EGH66uc3ZV0GAa4XTNuEHq1muwVgF6lugRp04ilCF8uqGNKjSvfpDFSuU
HQ3rvQZ5uR8XW5PqwouSq5FdWJvubq+hTl7ppqOZfWtyTi5yMQQyE9Z+OGUVWSKao2SEnJMwtEXl
7Aj4E4bOtDLV1lmTUC9ZWnQYd594NND0F28cSctaYPvpQ/lD97kbJUGYhHGRfLHB0s5ywSO3vixv
woGMxdTKu2wJiJdgIiTqpDvrkCjzu5gsM99E9qf5CaTmrUU2qk4DZTNwR7qj2hu5SFNHpEqwTcl1
j7NWmT0b+KQ8qcD0RP1W8ul4OLpU+XeqD//Xvaksac3D/DMX/JxVJ38XniwGYXkhRN0OtjtcXs5b
oN6PMR7WCRXaiPFZ2Pj+6+7JhuUOtqAQ3yJP+EX1djd9M2i01C0IbJSYzyltauua0cVn+yo1Pn4S
6Khj0vsgFiL1gjJV84JtVXsPCggJgZW+F5FTXUVZirxJyZJM8uizMBwDTYZbfFANNIkOT70WVLSR
l1Sp6QiikAk7okIXLc9q6/T0Iu9HlkJZpoAe6Mg8QadbDrEwzcJ7kXi1lVtO3nQF09pjUUrKDSe4
6iqDPFOzpYYXx5HFL3eGo3MXefwVh38/gkWecQ0vB71oCK0T551V6vzF0MZoGeyXg6lDFK6nHerc
858Is8PMQQqDlG3JjP8trMxvg+lH1g2bWnDj8DdbhO6E7INOqfeHTW738MSl2U1yGSQMo36awkev
oSpeDk/sNkQg3jDplq3YKMekVm/QHQNeaZt1XWH1vPI4UgfS+N81qpovRM8TMw6nDb2RYri4NiFc
tUqRdf3Lx/9J1g8I/CkiiyWCcGMbeU9IgNYZeM1e2ejo3yBTRYgX+u6fq+eMsOxn2lvAUy8p2N9u
Ox9969buF6mcqrsM4NG2dqiaqTjRJmdDktCQDkyklUYmnkwP/ekYjco3VtrIQnFAhxscxYV8U3bD
EQT3Ma/X9gNckOZHqb0TxmcHcrPvVmK5Mh6mvREz66g/wl5c4UuRmdCUxydRkJ2UBo6CbC+Pvc9g
RFcbcp00SAkT6SBFvZu2LQU+unzPwkG2oThWL8qE+g4BUCX0wxFKN7kSPhF4X41Ayj3IZizJLWUO
sx49m6y3gyJexjW3edHkKk7s5I2NxNGRrv3Lk13yD5i2BcNy0IbgeQDjbpvWginzOI5N94h93xbP
UjPdWrBhkpLJm4g790iU7rEAYu58PE0BSCpwbTgQL3Kq1+9nmv1YvrPgDObh13I4UGGUYLDT8yAH
ADzeDnCxJLb/nJitIt7xA9uusaLkpwgv45Vv0ILEKJzhZ2IShxc6Yz6GXnSClZZmUf9QKzcn3yua
v8jPJOXj0780RGiGrfFRHEHGTolckkK8E+IlNX4Z0m/NfKTzB3yNY0K8Cwz+cs/b/3+fkFhYXjm4
2k2nuCx9PmfrDZrzMeALKKTWnoQnx4Xv8ai1TOjlMzXeiz/rIc7x6dEJYAGZB8fWHZBnkGP6Oipb
WWLQh5E9Py47QqShUwz25EYIZ/9jd6Qfw3C1MMnRV1aOIn9VaBXOsOvpDHOYALgHUA4O6Onx7QB8
lbqtQZ1G+VesymumcEszDWbDvEo0o8HmpwIxRrvy3wjxkeLYHS04N+GIiNVuVX4UaG//G1BMungg
4Ecx7Rhjks0AKH07+JpUkOWqFOMZ6wvLOoW/QCnLH6tEz69NmYcRtngrSep44mJbpEy+H04gR5Fy
5SVFhg/CgGHLMPLe6pwgwQ0FmhVgGCZEgzIDIu4XH0ZviRJ4e9FHyl2CN/gvolYNYAWiYQGt7XtI
9RlMrxiKN8wF7aCzZrBBRycSB75M92yxwSLp+CBkY0ZX+MT1eby1Q44MXwZpBzlu/BLxLW6do0LX
8HozT24JOfjUMgmW3cUSQUcMD8mGVnCiZmuEnPoWnPnLw0hMMU0etVbmJBnPJeA4+bv8yKpPXLPF
oXPwM+1ZvIA64Eo1V0jd0iB83VDUFLlFDznUEOnx/0AL+0h+LKaB6MtCGzS9+k9WRd+r7ykV+oDe
Kt6oJubQnoGvptaIlWYqQndyVT1HaZNp+OCJ8jh7n3V1dL/8l+cetgv/8kL8ggxdjMk6qe0rrg9P
euwYIt///bmwq04LZPUrVlExKHyvjKux0D2P/AP5UJko+CPoZBdpQS9KslOx6yagGXiaega3I3w9
QpKCZ6rCLZFUOS3N/jkizZibRJw615DruMbTsAiHF6qCHzVn3AmTqkQzpyKVIq8pqMZ+H4KkIuF2
9yGqgOUYQB+CDpcdJkFlbVBGsRr/NkDsl7e2SCwJu0syCT/MaKVDJS6DjPewyLjBKK9reHiGn3yr
EtCRuwNPWZbzp22So2w+ypRQSTb4MuZbSF0njdzeHjxozlcMIW2Jp6XtK9Voo/iI1sZbgiSxncnv
u97U4NgmIQ2wT9gj66AQuhe4Nz7IX45quY4VXH2sDI8OudLO9NgK55hJX2wMDuBeAK/yGZUNZJHs
NlNaiL6OL//JU7y31NPPFGcFb96F/WTfBedqgL+a6LPNHPtpFL70NQ0F9cKX6zUJ7LJeZ4VOuaUM
hesiBpdQ+36jP0zD8D4DYq6G6ytdyHHq9Rr/zNbNa+AFlA3uX6CADFk0IrfnLcuo3sUmDhTU7FK1
5mhGeU4huUo5MWDdil9okwACfsbxvRmbdzs1c8Ciajsx2VBz6kbuouGVZeZz1rfHafa4qx+6WrX4
y2dg8Jy+/9HlTdyuWJAX0pCWB33/eZZRUeRkhdO6JvTKKHVkxK7DeLIMKVzXk5i65PV4Z5T/03m4
HgrWIc+5IM9TrnYlX3l8rKrrue77fFWumLNCiigseAWclLWQecclgb1kLyKD5nG8XYx5TWXgUlh2
TehSXJ3ize5GtJI7+EBFWfZ3YPZQOjnGRcHFVStdAFJPUx6EgL/QZlX2LSmUjHppv4ao04i/qJx1
CdC/kTZXPYBMkuhwdKtCqa/yc1xo8dNchjb+rRWvNvcT7/OacyBfwn5FmO4ctfFcPT2WNKmZSOK9
SIY3TDQDLPfRi7Na2stIMNL6//kpBNSrcLRbLftK+c4EcNurRuJZMvPsltcpom8c+0eZvflh1/Jm
bGEmAdrAJKxIX+FlF22VfXwj7Ib6DYWFg1ETh2mr6KxY7HD5wxlapl5Pf+Ia765vRIJADhhnk5SL
jePiDXtY000mH+S6KGl8vm+VLeJ40EqfCsWhnmNRBL0G5kvsUDePN5Ub+UHRJ5MWi3/atUQwJ5E4
zNlYNtyptPxIBNrHlHNzZZIdnc29/coTJvrtz7QekbCjKhv1hxYheweAsUtrCSAfX0AbjA1qutWQ
m3MCZ1p3j/Qz01ZvlmyB4nffIYjVvsn2jf71KWpwuGCphhU3gNnORwvxafni9zyJ632aVf07EZnE
azZrSdEiMXYN8yhj+CBxzgdXskdoOTXdMrXrvm3tBDuC7wylBkwPYnNxILQAXAvQSiG31zEFwnJ8
NH1yj2dxklZpOIM4gyi+F7hefTIPdyxL0mBj8bppkFviAXL7HdlKyyBHO7iJi2P/K4VRmjQlA+lv
v6jw3wnlbuWUTam++293lb5a9lFNms+K/yUIpS1Imq53y54wCF1r+V3xzOG8BMOYUfl8z/0Ec3az
WKlOiAMu0KyCpvpzgj5uESiKZVaM2uNPiryiIgcic92FGMmrBdQS29W1j5mbOiGk860Uqkp7dqJ2
Sa/Yw58nnKrlcT0gxG0rLywAcIYUIxq7G5CaE7gvHcF9KB+oFqsPkcizD30hrYssc4qQV4sDKVHm
ptxkODERPK0YmnLGZ6GpGFRbPiaIMZxxWM+SqCWrszDRqVAZu848VwplE6fNTJ+a3nwP0O5WtXQv
VN+l2pk5vAUh2HHofL1UbcqyBIpAsh4kybIy0phwkMiUje8YQOTVLjemL4uJO8/lIgDkd7GBmYwX
2Lk3TOdcCEpfh/LuaBuBVoV+90DD09qVuC8jsrANLA4ZIdv1/MteHxzUy/dFIeYbhw7xy+jE0N2z
0W9159NHgAvuQZEfVLgnA4WTwTQ1LsXHQvVx3CHssATijGY9Kn0YbY1s/IVr6qE0pnfkEed1Mp7r
7DKgzv1JIjVpJLtimSokAfy7zG5oGmAIDAKcuubjXQxJ9tI30q+o8d+s6HvbywKez+w6GoHyucKA
8tfR+qyIhv08TiYOB3dRDEveJAV4+1/Dk7Cu9lkBOgpaW5DlDFCyx0mwTxZSqRgUoapilw3pC/Iw
8MimKRJoZi6Mg8xeGirTQw+0wCiWYvgqaErje/MzYe5OyT5jdX+PmYPvBN/nx4IkZomUav2ggPbf
ZdOQc5BtmYdjOmWGxISW6epzjdlw6OsQo5WmllgAyci8pusy6odugG5FX4ltG1Y5/MaXLjDBRdI5
20o2FgXjD0Zl0GFrYDdaN2rvdy73NdXWQm15o1VWQ3bnIg5MVQxyDLwCFV3Ndjq5xzgLLsZTTigd
HXVl+OV6VgaKYeOf9DzXFhtSXW24x0yAlwmhgS8xoUCDe84FnIeLTg6pwAeoogRdRCqbEpHV/dH1
q5cDMMoe0JTWd/P14U4LEibywBD6QME0vf2z05tbbbTwF3WC8gnUiWVqbKolrQY5x10xlP14KeaV
UDuBUoHrTYZXWRvfITqiw7Kd9yC88ZPhlBxvV1YQQ/EFNzThYanhNHs22HUh9/XV2IBwx2m42d6b
FLvikvE2ttRCj4ApIPQDY8rmnKRUhY6WUzUiAu8y1n8B985l0Z5KAP/7BnHTSBbao6V/moZcjF0A
UJJkUjZ9objIGjv/7M9M/O3N5KEz+P6/T2RPrm/OkKBZENQvVCqEkiltXYf4K6wZAQvzADY7sSgv
Qa9P+Pev/YUptTgGuhML3frLYuNPgq5A+zk7y7YpoICiGyEP2lf/i6jLKtxgV6OkoIPHZCXVCiz6
/qI2wLNgWyoO/3VxnBe5fk4kWFz5xCyhQdLY7hn+JIRcK2x7ZvalxfuLat/KfZOPViYzjKvlkdVW
SoJhpPxIX8Fu1nUI5ge5KhvEHHFfFBsxo9G5AqR4SVNpxJPXKReDgSHvO+tv/VgvFd3P5v+3iS/O
rNZqTyutZKBCwD77UZ3ID6gRn+jRXk+ciYZhVw0o8VVgdcy9RUANeEhmg8CpEqmT+RMANmkDmB7U
XkFQRga/O4arffu/gyBZGPr7/xzhhbNQ02ngjsJX2/OuUIhGa1QinVuQ3qoyBL9SpfQtbi+QSZLo
Hjn/+STdsnS8iCTd8AcKdKnyfAxGrQ+hsoFHcDAhNp7RkaVVjE2vgizq5OStrNaIxEwdid2s4+eL
Ja7M6aSc4NijrEVlrYzFMwVG+MarkRmkm202N0nZppAY10ZaKMWh+M8zr7RI02MIPMSb5kBaE7kg
mSVSVKpi7zwmaSIzgVhXJxrLIUhhv7aewDM7pDwlIWozBPFn0j8uXotSn0pmzHdBJSnEonLp67mK
4et+8nt7iVwSppMclf0ffTbdfmhxIJshCKP4FFxTdZllbgiZfDbWRQD4V7lnSosYK559ZsR1GDHx
9Ool+Yqk4BlmMZDf/djh5e0hoTOVgpGq3RWix3z7a8fsY3jxKssp6GGSjOF/Z0zrz+e66LOD66Fu
gLjLNNYsECRbdXS88o5YTsrEtl7munGrEkwXEhzQXVCeAy4QKE0Ay6UjRY0GdJcindrx0MRR3Sql
mGCEU3Lixx8PbZvLIblcNvXIFDi0q1mjCoXp2YArjssNO10x4EFWjRDK7B+6IpehgBXnhyamxoeq
21yVgKrsSC4rGwRn6jrhOlpPpxKoG16fP7TbOqDD4eRhLKQyBoLwKW/PqqVxdOwqTho/oXIa63YO
01+q88VWNskph+pyTBorjb4WxPgqcymdMUrNcIUcm2QmgEfWMGw4OZMfqU5QWkjMi2FIFu851L/l
wr1eNc5XqniNz2D3Td34EhJVgd/hNOkuKUZQbb5irIFk2okhoJxgv22o/QY/wi2DtRzlf9jCp8LH
kgg0oDJ+1PXqU4A9LulHKs1ytKrNiu6KWD9CoX5xfXND014aJR7kNmTYb03uGCTgWLu3IoDbzsvK
KeoUbqf7xaEGB/+LvyCgxtbgcT9RakjJSSXTEOcQ/FGMRwPMTB2c3D4pgK65Sj/KQa/oPa05JOO5
PEUctEOIc0esD2Ds0GORZ+Tj5npUWzIhfrXwUeS4HDbsj+p9j1f1RG+C+eRftshVZP12lF+HwHEG
+mCx505WtEa0KBuvb+wWdFd+NNwcG1NtObm+1C1YBZcN7GgzvdJyQwU0kBRMyYZ7ppnwBsMp364m
lAm35YhDSHJz9T7jipdulTA3+0gyMr/m+ApcE/PsmxeS24Zbh56VfTgVJEfUlmQC86AUJ9VQJdNs
IDHSXCUBd2fh+Ov+AY/AAnMQj0X1gxOvmOYq36abDpbBFpzfwdgU83x5+zYp8B1hDP7OBDSaNOh4
oZbXfsaO17Z9iZdyPf9PqJbEpUp+MiX1/A3lMC6YToPCLOkVWL2Ol+Efy4e2/yQqVlcpk1ynGJAs
fUmSPzfOgMDXON+VbQRwjmYKUzUBsAoUXmIdkcnkOcwECeIFj64vgOlpVYoEW5qrQzXhuvXAbges
h4PrQQHCEXJ0CCSwiToHiOoQSb6WO5B85n77z8CBX/wIrTabCT7ap5I5ICWsVMA3XhWvqr5jJ1oW
YJ5rUWlCvpDIbUs0/wpqzyPSQdR46zZru6D4SgHxQ5K+eEBovgSUYQpvTQuxPo7/ShGosj++5CqB
NnpT3cIkeZN1v811htcHR8ITokz4WmuGdHRoO8V7BDj9G77EMMfU/GZT5vcAzhkqy9kOtaNVaIBp
IFd1140ZWPLIidj129oePp5L9xmRzTiUnjBlvEDcqu5x246RKCc/fH9McusrfMuH291PPHyA2YxH
Qd5tf5IuS6Xyc1J8AsPkjyRIIMwrhv6g7CapNyylx0ZuFwyC/MeHhfUfuRb9iLoffuzU5A2dtt1R
AViSYF69imPQDZEGPr+YrBke1NOfaLVE6suFkZuRzSrbx05ixl7YK2jlDhdlDh0rSk5ruZg8wYeM
GeDocw3AyxCHTfCaFYOd5xbIv0oqZpBrcBKrR9FFodJwmFQmEyGVLVYcq6Fzm4jMWraiSw553MGX
s2GZIwpyb6yfXiVARxSWWRN+x7PsH/lm6GnWVWXdxAFPf9kxWAOWrwwCuVTInKQmtNK+2IrTNEp/
q7VZAdnDB50vG4GdqqQ+jR/HXN+Ej5yu3YEXWqdQTDTl+JXebyYR/hq43UrR5LC1p/qfIY0tVcvJ
LCBjN/7r0mho4Fd0iYAL0AAGEKygUbIf/VHL5kwknaPs0ooshlfYiBkeREMf4IcM6F0TKkVwwIhf
1iBBuKaZnKisbGsjJggHCW1R+oW4rY68YulsHa0lq8q3TTxM32QrRqfoZKwNqCMYdwNKSOUmtfyj
EjK6FqtbWyITCNtAfZJ/Wp7EoIMYDIt+s0U70AJgNAMbSVDzXX/1cMVburXjLO2hH1QwcvLdwn/r
/Sev9i1Z18105FG1MZ+0szz+ITHR1HMkz5gzdly653GXBc9raUW58IzzXjyyHH5YwIqp/K/q++Pb
dtUwp6RFiehiozFHfrdDyzpul7Z3EVGdsahmqDd8RYKxLVVdPU82MJoupqxOze0laD4Ccx22/Q2W
VyvFq41xw2UCUx+Z2p4DMhpDSmUnOpP1FDwU0GjighGD47FY6YYRrDNaJn+csG2ACCodZzAVM4lH
07UYX4F6Ti5EcmZM7LQczbMgSogh4o3MfyUma9DGWwKbPqxP8wVwy7eOh8GefU46Cg2vEVlWiAi3
VAtvY+Gjc/Ztve183lgTjwwie0qpM34pS7kDz0nxXehREXuCm9gQfK8NEj5jNxSCgU7lVYYF3NEk
hEagimUQ2hU9OQMU9TG87AgaKEwNI2F2nm2Ya1rmg/IDGPI7gZCUpQYSlKK8R9sXZn9gG2Arkf6f
pmHcgcgtOoUd24MR4rteklXJBiKQqxAq0G8wgbxt3zMPh823LcupOoMT874vVmRoWdKXZPRGOdP6
bTMtTEh8KlEx7g0PR/zKPGHunuAocQ4MjUe1tch2ZOqIJ8AQtOSvC3B2MiryarvWZKx5GSyeNrbs
i+jaxwcirOBe3Byrr7zzWVRmV/fBVFthXKI/7CBR+6lIaJEY4EkQjRajn/ttH8y6nsbjgS7K7/kZ
K3f+e206fm11dIg2PQ9fl4zHlNOnP2dI1XtNcavuNHCpZQ8elSqR+sgMGAT86AXsAQtMXGl36kne
l7UaZDHyTZdKX8P5wrcoET1d3cdm32qYkvW3L3ntNN+LfBK084HyUz9e+YOr+IeMoV5pMRZSAwwR
fSvA++BOScXEtYgEL93LDQq8NMdm1xih9Ip3qjCn8e72N2Ll9ZJOCm2nalTy0DacXw+t6Oy1ZvzV
FX9ZfnQD/txUrN2Gj4O1kdBzklvXQJdL4Xl6pscSv2r2y3yGzXF6Ngn0ePVq6EAQ3mjHxH05Mxsz
C8qk1MdlQDyWAxG3IyVUPwKiVhogcGygCm+TosnW9KsZcttAlQ6W5tne0GIDOagpxbx2Qyj19UJ/
JK5HZC5ZdtCuf7g+2JqFBpyHbJ1H+VND2l2M/shXkEroQ45GtwsodgpDfIdjDRDl9NlGxFxdp2jb
AOBlQXXT5wpWeLvusTLWdB9vATRkw65Gmmy/olXuJDWoM1A+afrJoF+vU2vS2+qjkylQa+RJB63t
t2FOtSgMdLfn144Ij9610kG/Gem7fPrg/eVHXlPRhqq7y7qjpUnmkn8zwSMpRnyQkOP2IynFQgdd
WNbU94u7fENeQf6K/cNMZEzvPr3VojDUs/fZypLg+061+XJCpPAo19LOp4jbxerfMUr4L20AAd3O
VFJgLtQkvLABojeXtAn8lKAp0ADHqiYrR9XKbRAv5+yjTqaHSIGc4D4JwxXdjwHIF44ZIg6kgXlN
6dWEF72yYb/4zVKSxen8fZiEAbS/a3IeMNStmY2csFXcW5VR2eA8hwFM2MwMfK55sFFwn02wnxPJ
maM9r+IvQ2rhWhZdTkx6rbe8kF9rcprv6rVwvAO0XeSgYX0scy+yGt8Kff5ZsYsxzp8yo8hVFuKY
ztzTAQjoMeZ55cJJWQZKHVOwrU4t3E4MCNHn8Y8P7MuhmBBvqV37aa/4IzJntWdCavptgzpTbPKf
RaPVzdYWvpkBSJSN10uRL3B9A6ZIGHF20dOYCbRpKqMtn4ZPf6p5Tb/GCPVvv2y8yk7IskED2XeJ
3wgHxaEFYeu4jwy5JU/mkBd6A1Mx5SNhTmTlUHa9/e2OTGnMqJu+9fPCqIW88/pTMc5ONYNA8GG5
SRK3cAjZERgEg7c9SQzaZbQZ5vxQGhk2DHiSQV8ySKaITcWj9vmqHWPeOnR6VDhwugQ+DlyxXDzq
n8kambL5ybAs2VibwOz6iW94t1Tbyux+vWn/f5oIxt7zTMij/V/dVZsaPHo9Iz32Ap6zr6DNoOI5
yJQJKRjGHRw3vCVxN4BoRFhNntA1GoN607Xofj+16z/XzTlsd/CWNnAilP61DnZTzhGb5ALh9xFz
xZf9FYLt+haZkJw6wa17WUemEL9z1vcQyFRJ5QLjwmibfe692jI3JCy32AFG3eOS9IBIgOgBtDg/
banMdO/y1fZ0xDa3yxChvKSCFkkb4yjwosRdALDwe84lTAAclKXAFUb1L7IYB18gJ8z6yF1vK8Gz
wk/t7FpcRFXUX0lLQBdPEPZveWjPabyFZYLOW1LJudiy1iBDL+TNtCIIuMay098kisSAi/dQemuN
+EVix3vCoTUnv3wvqakJps3H/8XyNsPjvDRmEgM5y4biCG6Qive6IWj3gdSTbd9PrLwESTD5CBZW
A8+e8aFdyVuUi31vzvVC9drn3hP7XvRdy1sYdBClvASv1lokRvCUSzgoBC0DyG76wDw7ccN8+3I1
y6zNFoGz3jASljb5Rg5Hm+GPMLp+jGjfWY7sZDpPJqHKU4a1j8gIjSfF169ZfDRImbut7Dk1RgPu
7IwMqiK4NjKcLcTLaxfxrcXFNYfzvz7LAKd+aw9iEvfP6pmT11VVVfyntBpG1VB5SUbdkd2zgd5L
6XwcgfX7cwPG1TRqSqqu+MIRdY++prd8o/28bLhooqOw2AaM+n7E12LUBGuZ4eadTLCLSsd7Lh6M
3bnIkY8tmfppUHSzaqKTEefp/9F4kgR9owGxe+DRLydvAcsYWU/7zK2XJ7PRYv+5MbVOhuSwAre7
WJRfPddkiumBT2+b4y4v3Uchv9h++ngqHs9f0t5SsdWc6Q5fZ64hfhyINKq9iIu9rgTSAl9J4t0m
oogqpUf8o+A/fAM+dmp8r35HKstGLuSVkx74ZdSNYHugUKj52qFzsNVIL8UppGYpVuc1v2gt2X8f
opAGVYmF/CuxwKvnDWaKmzAxV+6BXTzwTUZjBoWvWsZXkUqpMkZ3VrA+vO7O+ssiphDgPA+jzmbJ
vkpjbV0ddIaukVnLBezcP/SWrvex4cYU1Z+fNgDdPwv7Xs8yrOVYqb+nqL7/nYRUZ2+qytPrGlSI
zdL9ThmU2GBbX0jxEhF7w9LKvhkOGWkgqitYgurIIue91mUNxLiSyQJtV6LApAmSkL3kuGR6xFH8
wDelZPhRgp8oDieJFgL2/Fv+umu/QIXhr0fHfpGumm25g/ENxyLM1vPfToLg92RRzoRwCGNA/UMB
5lw2qBvyN5BEIIbfScC03qfvjdvU0KZT4F+PjnibcUfh8LmO6zYLc4ccgD90vwKKBbekow5cCac0
B+SJol0O9Mk01FJMbYoSPXQjDO1jY/i2Neg6Jz8yphe3Vo3WsEgwf203PHrfwh7ly6FiHxK8mMiX
0wwo0h9sFteYGLIv19Tbu5i3xBQscHnF4Saz3z1TEa7L3NPHDJmYrkGGBgkf5nadQg6LhXhq1Wkz
Jz7g6MxVZufsVD6kcoR9D69GvMPyLv0OkMJxcsKp/TkG3MifDeqT5Ln1a0rNCZ3N08ojNUqAyQva
GGFMtQJGIFMEE8yky7Vt1f3SPdX68TMW5Im4wLThE9r38+3xoBhiSCslqI+qYE7Zr0wLSjyMBDGs
Poz516y/3udQ6fBUe2ZGu1drEi7TCwnCIAgFz39QJu5szCn/CIFgr7oKCfBX49t0EY3TpgR5mfPF
LbKYnICaEXYHzW3o3zQFY5jNb/yOykjgBSivKX/+BDfCu+CRL/ZegpwhlRQYUTWBbXuIo9U1eqnj
EeSVd3ohAFxsnwarJYi8uEpxo+gEJ2+Hy1PFWuLVphRtdwmwc0ydDvskSMr1nyoOzKIxFDtUwY3s
tse1C0XbvZm1L8x9ie0SOsgNeWyKc/y/urFGmIvf4l9OidutpYzfhnFqxmHr+GlUwUsvK6wEQiUP
hhvFzbvdMH3FIMvAyYwmrA2lYHOho+SxKthX8Kz+UtDRxwD1AlJyR6gznTrKdhLrYGtrsRZfaz6L
Ymm7EAzZ51UeChm6DSHEF5clz29ywjXADExyOGzxw0BlZWjVTJQgLWFuQZ3TIOnKDr0aags2YcJx
8mUoHOKN96Se1otwf50N0qpk8+hbBUyn8wqfpke4fNh/wc878ciLOq1GegXAmD5IhEaWdZCFtPi3
YuiMEmnL+57BCyQbZI7jF6jbtIA0JWca9L/qZM7pqyk5szVR9d1rYBCw57VMd98BSMv+r6tifqm1
IERsnIK2ItlPZ67y9Yg47dZ1lao7shqODYNlhn5IlLnVJMhMHD3Ckl+oBntRj+eQ7oVMRLC5+0K8
LV+5MR3b2LTNC59ZnoF3vfD++9XhWdNbKjHIMe8i4/bM9TfE7IX5JfTcxyOicq7ay2Vl5WBHhOyz
pqyLc49ytIkHJjQqTQeClxFgwXDa1oCrvUTcoCFvSymIaHgq4gHujzuQlmUWbLSVDw0wKTRyuwaI
S290k9Eat0kZAnhYK2DtR5aZjAnqu15H8jR9jlB2+k2OcKUKzODbVSN2PVZtjBMRSZTJhg72ujQA
J6+PELvs3iJ6xsaWO7MIof4AVyAU+qHbxKDp5eyghw2nwBX1yXD4cjTMWcIhi1gC8VxrpCOE0HT+
pVhOA6EunxUdXcfXphVVL93WzGyORmGqxub2vT5KfaI92y785f1amYJXabOcaJf1me/XhBQYl5WU
OHVxaELLb67QXgAravMG4Z8DDKihaf9aDFSq1WCjIMnAqFFEtiQAW6iJB76SbO82Cy0wvK9z9Xnu
8pfTsNjn8T7emeLY4lZIjd4otpP9fiKhho0+LDBdmOFZpaYTmINq/6bMn5aM1TCnOankq5romP+R
r8Hcq0ObUZGbuv+9FZWl21NmWIeR/kvjrTRMOPz7WbtLxd/cB2ZZfKxZlLa5ePYqKJf2WwpbUq+f
PC/etuk60GnTokBKpRvXnJwS8nCHCvXcnYQxwMVgNF5EMn1EkbB9FsOaJV0s+5087gKPlDkEoJCg
uHY5rp2JUnntPrlltHlZH+8J4f8qGlteZq6jqX77LgiRKk5I+DEmThJny5hexCTXVwD4MCurZak5
hV9g83vrdUS4GkQlC77yFGwNhV0FgXOFxWJFpSX4dVcZ4bKztYSCHRSJY4OZbXpFGOnqbaWShB4d
4SQogd3cOxxNLMH7Vwl730UaiyINlqiqVVDWwaNP2xPlR0nRnILkXNnVUy0zQcDuIFid+Duq8ikv
NY64d3VV1uXtnVE3fdCWkhx6dtUIiYjHNEfEL1V2iVitSxBRKBUu66XR+trVcPnfwnDgr6sPvVrH
wY8IsCafcrQpdjjSVlAa8rflVlp5s+ar8h5vv2qC0olcYjb2VtGTYkwJbXVxQ5cUCmcwGtFiM0u9
ybGhnElKgEapFpydM7qZXRcshcDxEdNLWCohSJWQ3mrBcY6MezbY3v8X2AGsW/cSbDFldhiRUdal
4v/FrUdhLh5PpH/SbB0kiv+rGpYf7nkrc/fezSv167e69N3c0FTYackblLo+f6rApXehxF1Qa9yd
L0A86oDPAuQ36UpOg7qWur0q/9tZ+1jAWZ2+dwny3oEaa65rYB8Wab1YbVLfGDpvCFtUNPmpVjYn
tPvLSETzGJg4nNV3S6rU6HfSLaYvpl29jzpzwpPLi7shS99rqtBwmqslOhmiubXvnBeFQAWSPlU4
13ALmptgg3Wjk7BO/XXBfbrUYL8BkU2YodnKcxluCo7gQyC+Xv2LSTuKXuheLWBvY/sAVSdlmdsL
QIlMFJ/AUlZ8O+YOcpd1lOcAjzVD031DpcwuP3koUixV13W7op+tWRjaaOZgIeS3NWr4vb+eBp0b
U0I8BtQLYinLmMSigoOjno1Os9PYvdUSFWCW1KlohhdUH8/pwuEW6JzNY9ZYjE3vKYeUwJfWTP8u
vAgEA/TTIXEmMK6ClUp0U4u11upkRD/A92IwDhYiCLIwpvvaUBUAkjPaz1hVd/dWPOvQckDJWT9h
HCZjTYBFD2h2tT83mMID/x7tA02Myvfcfdj6GUlqsDo3RyoZA9iLMQWkaS19I83E6K6iSFP8Np0y
OiGlyPIbpu8hjUzj83nNuW9T1p4bDQExHgFmp0xZIcffdNRqIaPOb3beqcV87FpjLrT+IxQ1IDKv
MjusDQ4d83jZddQu+0l/q9Gir1cdgr/ftY4SAcChLxqlpSdLjtxuNRliSNFR1YiV4ldwjoo81Rfu
0/SieBVep9OiBJpuFc5SHBNw+MZ6ej+gkVM+MRFxx32F6g4ze2k/qR3TOM1j8ctOsNQxNV69Aqfp
eXZf4fxu88t8vy6RujzfVggcud2IF3DUYeG7+0+8+5mEOvE/eRlsBvHToXs9VAgMypVud2fEMvWG
vIOTIktKWU3K7IF3pzV+kUP4VfueQbjjCrWhc47YMk2Pod2stR9UgBI+7Xtu+AYugBrIIGGNfbn2
ZSkNnjv/DIOP+Z2WZhVm0TOGv0fDVdwu90iuBbwnG0XweQELKh1HPTdcITf+BLj/VxezgO7A+Izk
GiJ1N9KvYGGUK5H0Y/RljuBh/rKv8fogRkdGbkEn4LkJ43ZjftZpu4Bqq3SbNeqbNhm4kNXOq3LQ
XCccni4fNZsFH83sEYSLgaIqX0vOQE+FmzFI5tsnpnNGTMq14XW6GYDkJM4nUHUrTY92OVwt+AYC
Y0d5lUcGQo8yluyLzwK590vMsEuJDZ9SKHJHXe3alZvT5M7V4GLNqa0s+Ssi4OxIarz8/LhTFHdi
vlsDN30Cv9qSjfsUXX1x0oWyD2/60B+7JHXmIQXgaKSxTwEp+pyMvRk+DzNBST/Sl8tgOvXa5XVD
eqg8YasPCpU3a24UKa79e0KPrXtmIHMy7gJy+rTOcrvmQcQ5cpn4hbLZY+LAwsHq1yQeMlkM3zXB
XJeRQ5DJiN29HURYa7qZKp0jUjc4XnEi+qhzVaDXh+MdpTVbeYCdlFFo5EJiiSYSJgJBPMiLmwoF
M1gd2oq/DZ/Sh2csfSqBOWQADCYV6bwzLTH3xsb7kgJbS6aotJOHlxtyTn8P27Oa95ua8PTqQDID
WuYHi0gGRaQ+E2jE85fi6+bsEvSDHKwVzhwZFSeRjq1IVJjwepHq45nT4YsAcm6EXcCt02ug9hK6
wlNB+apTwqdrJAr/Z4ARJ8ReQphWSZ1g29/ndcB+N1YxDNdl3IueldaQyBiak/Q27sz7RXtejWsl
L0b+BfmIHuUvdaAiHnpRgLF+6Le7N1sFzXZjLQPtxOQw5GIVOuSufiIgfscIfDo/8OmX0Rwu5HQ3
aRlAt8sAHq9qoR+gCNgjAFY29LNJ6+AEVk0nF2kTZ7xiATu9QwClBnFxuCOiXVVM0a4gjkityA/t
pQvXD98jcDDHKGhBoTZRQ6+tKztipDs6V1NAlR9fBH34126mph6cKCQbW4VAoQwVXXhlkgocCVmb
v1kpW3zWpFM0NEXwLaPQOMDxk3en8MdhVkuoJAGNRDDNlpyzo3fsOs8AZ3eFG96B6O1hWpsKjYhQ
MvmgIfYvxJkifnheMpBieh2/1m2sPLXtWVX2wMNy0IYM5lyKbR9q4ClIo6yk4cCvDJi4XuhcYAPz
rPA+rFY4yQBC5Ve0NmFwv28gRondYe+gPmpMkeQWe6a+M6L3+cIxudoakrN97ceSw8L3WNDQlHWD
Wq69HrG+tC7EwmTvvdUimADTUFonq3/JNp0iwwZ4745zwQRlfanDF1cvdB9nWGRRAWhSkJUecFzU
CHFc9dILIVzid1O0yuOX90ecH5vZ6yoTyF0IQmVxWRAcBqEJA0MLgmVJWYZqowbpJuDU+sfFoWob
QjeybOsixZpcrUdYU9fE4n5xqDdazCtJ9IfAs+V92etSi5QIgCFN10NNyyOijQ8gBmhLG44d6nqc
JUt7q50e7d36vXPrx0LNWJi8wo1Ut5x2NUiemwTO4K61UASTrYYPQdwMuaWCnTS7O26AvfVrIU8m
Dqn1zPpWAwW1QZm+MIGkIyL6kp/Nnp/9zH8z8/+zkDuJ8VBE7pm5IWPDsXq3Jvd1zbMv2suJY6kW
UjtWX49SIeRD32NxokyRoN1mpXTWEBtRmn8Poeixa/hizQ3iZG69SlhN4G/4ORcebioxu4qjZhBe
vkZwvX4z6larYjI9c97iaMRo/XPJ4VbnUmpj7sEBpGJP9xONVjt58Bd4m7zHgPhM5y3DpHjlc3T2
VNwZrHKjEImvsqH7r8IZbCYTaXoFv7KdrPVCfEdOEyD5EcixxGqrTLMjBtz1m/FCHBx+qC7LY33v
jKuR6/WZwOQeRwYcN+p/OaCvo81K3SwsnNVIIO3zF8HelDxPq4yXzWSfuySbNBs6TBzbdxrGNkNt
v1rjMJFFvBk1KTzTOCiWE+vtycH6rW5imyyBojgTtQjv3edV55gZrAwGd5Hg++Qshr98IHaie8Pi
esoDcxYhvR557dRTEH1R4WF6dTSowQsOtBlDDXaKBh3pKN3vZex8QBC5uvxKQj4JNdeNmc6ru4hY
wUufM6WNvNXaEBNQwjdk8PAg+nHVFBUjxlKzG7Nw//dN05DLX16KHrZ84XF97i0FP7/+4tM+hza8
JGrvSXsTIzKNUZ9WqyGVhmU1qRj+C2yhNN4vaFaZe0+7sMCVRTxZZZ+PCeBREldeSScMjxkGqSgi
0EevbDYKtUgpoZXT2y+C2tYLUgxj/vt4cTN6BOyNG/CW4GZcsCASYxh3nNrt3JQ9kDKE+TBvmWGS
ufyfORdWqUieIeDz9SW14yHHi44Zj+fqAvPZbfasbQZVDqSiAE2znbV3ZrLXN7KUwk/b6XEbSR0V
fuP+xvzvuUVCg23wQSxJ4QooWIiq7xTgneFmm7AUIGf6airZz/w4M8OTW957A71DIyW/EpDBohXD
VqMDBcrUd8K2KMzLLAVPZUustyV0YGg3GHqvtyiEOlwVA4gSrg5I3W4KqAL1EuN1CP6kEessaNf5
LutB4bd3eMhHTOzewKBwOGBVy6pN6AirfYckwg5KmQE61BWmE3CGZQZnscSApQyAsz3F3UmCUAC7
hLCQvu8Se4LEv+9Jga6P7kBP13uDnSlGng6sTARjkgOvXgh8Ew67Cmrj7rqthhtpUzc8l3gA0Qko
1vVOnjwR9mDhxMu6S0Z9sjIsNbeFGIJl8U5Xxg7E6r55Y1GD5HKcqlRQ79NEF1LO7W/bNpVUOnXT
89BCEHj+P/rF5SKTGzuqQSrL2c/bf6ikjJKiylZaurpEpOM5sT+w5BIgmTPvPzxIl4/Qjvyklh9H
6iChsGTUkkDFkulWtZRNm2c2I5w8amb2C0XMTjC4DiGtevTHhs2UxJqoj9hXuK2CZW3rJPX3wPQ3
ePiG6ISFkamR5AfZxHo/2Cz5IjSMYvGU9kr5Pf/22gOxe2YNqir7p54E4HNCKcWM50LU+dvyXxds
851kdDorWfE7G63eNH1ygnRmjqpZKoXz8ZH+c5HaxjGTs77zq1SZqgcbUE5ZrJS0gSLaAC8OgB0c
Tv5y5I9/u5biGmR4me7WzVQY+rSlGDarTeMFQCo4cayd9rgjwqj3IdSYK0XmR+wp5PiiCXk3npCs
NeYkUSygxSVBA/sY4U+Dfdmq4YZXX7ahUf7NfTmxB6s07tNgPb6SmMDxaa2e8swpQ8apGYEZ5dH/
NFzo1+aSQvjU8hGrj/2TFQ07F8cCj/Nuc8q3Tm5kdnmWnLtaKr35hkb0U4rLFjLyAIOxH/WTgG+w
gba6j147WAtkhwkga3v/kE/5AA2IJsaHr/CJz1Jaxf4z915icI9wmYSC2Ss3gFlxgv/XqzFCCavm
DJFlJQQArp4r8rbj82TE5mJfJLpkQVUYq/yxNfy9CZ+csB9avc+6qNZlO06d2XSmmW42R0jU6kj4
RfRieOQja3C2Q1oy7CAPli2dK3VcT9BN0r8QdtV6GVJnGMU7VQxK1pzjkRC8xQ9eqVdHpjJKJUg9
DNzYw+h/gKr16KAiIFoMYe+go9adKg7pldiZbx8s7E17iBNYrOO2GMPO8e7Y3aI+beRCCao8QK9x
eVD2mmk5eh1pOtBYxEarAVwhY6LMq/HyDDhEMaFhd8kVEIk52Zpz0GTLFtN/YJEFZRCS0IRuTBeg
Dqdq9js1dS1dsaOG2SHmAN4oYjWTXdtewJbg/CcXsucooM90khSWdUlHf/fGDTMdxOq0CxPRxoPE
T+Juo0xMfYgrddRD6wNf5KtC4LDqWPahyPC87sFtBuj57qmpize9kqM9xXcBxDKoA5QY9TJGDhR0
nKMVQ/oi5M89iWIlgNGeCUfvRwpuoPvKLaTH4pscMFYJSNjGJVfv7/69PmY98sv+A9tUq9Jg+ymB
0yXOPqH+Xg2mi2RAEFuqN7EpgP7/h0LZu5kdR+pB+V85iGwLAw5972gXjXHoy+bAno1tfTJa1cyu
yE3Y67vzjPOGtPQAHwiklO1YRl92GTLxVM3BgnK8P4CDX1SblTLnZUO93j0vUAqXumHfXBiN/ecc
uD6/Gshr2kpz1AneY5Aqmmc+7MRcwKVwyCM96qQ1yYThRqRL+hPzLqYg+BnVOwtnbHvUPPrvU8iE
OLNWavqTi34xZwleSgy5s5kqiUqiTT5cpFfloILVQZ6FC2wZmYq3WvIRyvYaIT7FgpgMOL4NpMx1
26UNR+9POjJwCFumJAMgQCmF8JFILZgT43r+Fszx8eGy8SAps+dUkLG1f0auzoM087hUeSCFWDGv
nlMr8MMHw16H4z+glb81/VqLCvZSrt6M9+R0T12eIHsHZw0hYgAFYSNANquKQvSwwllgJZqgsJPS
u2FGpaOJ+WfkkU5lQ0O1axLJIAiiNafvXvm+bE99HpHFw86d56LslVXJZ+rkzmQFpe79B+XqV9Kx
b3wl8w82Ah8j0zYcCk29daMhn1X4ttRqUIXuHQhhEQEw21FDSUsuzM5KzIfoHMtSRMPHfPTRpv2g
pN6n0wH9uE/AfsNVL6tXWxbzcQtZbu89qrmzGm+yLqF2DgfpMnbGvwlJv/OQaCCWhBFRZtOXTAbP
mICHqlmaYSxPyBSuDEmwqCk2LFGfAYPuu7LTULk2z48/YcFFpwXImRtgdJr/RqBST88WjJZyzuUr
yJfasP9r9OOmOW+k5EOyMEteqSetxRThwcKweYuN0+5jpXWU7V1eHwqcIz7txXD1EPEEhsOn2VR1
r1hNJt7nDw1wfmEED2ZrNaTfZe/7gqKuudtIRa/4uy2DJDdqzr5WWSk9TGACPl/NxF1v+WybXhtg
HRfxxklKuLIXUOB93C22ItxpTKJfU9/Mi7DlNTIjKGZIE+4iq/+YLK1k4ne8TymVMKnNWuE0LtxD
L5oKOBgXSRk9+8RdkXMHCG04xPOJx6/xLM8+ITPn/dhB6h1x66WNpUVbAUEj0zBEISqigisr8L0I
HjtcsZ/NU9lJwylATrxu2EMtjIpjMyGPlR9FBTlzJBVlH04w9Yso1rf1j/dh3ylJ0kHVY/TPjEsV
V3FzOAQhgdrYmI+sM1poxVnEZZkUGWWgMhxClCyZHDh15tcFtzsVnVHOin4PmamTkLxHTi+usByW
GcbTgBPbIRHskM6TBP5yObK3smwRiPW3ecvcQSTfilIhiVWYYP2+owh3M4JiYs5LM78bJIqG1LPR
ty47I3aRNZs73+IBqlxzLz0RpzsBGSRCDjJXTgXxEMNOBEszX34fNPOy7Ip2yquTLnd0t4O0GF6k
tEpnfrmeYBe9udUVw6senW+175aCKLLZ8bVw3a0ccUJLG5KnxEjJC9TRZ2LI4IT3fBtkbJmCuhdw
S0OvVGJFxOCQmmUF8nKuInp9GRubFDZtLOwgWqlHLQ5g5QQG1xHcR/BvSLeqQQ34ndxPpBmDKWuy
mNcrtFZgPxo765vNMUp8HYteNX3YmLKNSel0VQMDv22woDXs97xPfR5aKMTEATaUu/rKTHyD2XXv
2ruF95mSiPg/MjCnwqARTTVtZTonSnyBl6H+QYFwoRQOb5q+gNPtKqdkSyv16TJKndLCSdEOSKiI
uN76Vp1ZLQxd17K1oPUKFojl5pAKh3ruSW0MMag1bUYN2IUC+tEmA3eri5VnkSEVBGEXJL54OV4c
MDwrm7MZNgP/luPSzYmT/nsmDkNj8knB0YF4v+Vz0ObZ6+e5vP02ZANssNeXTQLqeCLhVUgdX3nS
zgHG67rFmmpdBJ/BgmKXHlFvhjyMZ2XjfR0AfktKVVdOEifeS3tVmC9eNTKGF9GiQAiTqMkNOzSY
JaKN51UXh6EaYmHVW1qNI14usWyrWdIbsaz+XBguPU9Cvc9KrvK6s72H1sb9qlYQ8SkTuC2OpRyT
wcY02MEE0KGKr5uX8s5zIRLWoYILiRnJp3NlhoqGQs+ccby4juyPlQZoB4EFI6HTsFn95Z5qMsJB
FHlPJ7+ZSiVyvv1R35ct8ouKRP6QdPYKeA55MREI2+dyArvdRhavhY7je9hPH1YeRIw481mcIfjt
rZEBGwP6W3lyjxzxzpZgZBzpFAdon2TW9xP9ygZLNYUgLp00Y3PKGkDY1rVHd7gTGt/bOhsxFaQ/
VssxD3cKSWzib3f5xRu5wr8g5yESXYsLaFNEeSOZoOHX1SPwg0WPGuNGZEjsG384TZDme9yhDOTo
92NdIfmrbapznpJgkaGmvk17rcaxj+Bwoa8WojfdWkP9JG8LUC67blZdOtczRnIBn69uRgFh9BM7
NiCUdbq2XXwcbsfsup8t+/Z68Puwa98xBfukTd0or+pXfzc51TKBtyDpf5YY2cVUT3rvFhpQdSN3
PImGEyctgNykaMbvssRCo7QRLbu+6qwMPKxMnYZp4G4PF+8ljP98GUEYBzooX6siV6R0tkiCosgC
lQRPyIUQTkfZWGxR74om+z0QMG38FrMUo5DrM2AOmYlp9SYWTy4xL3RTk+IZG3vSliMaxkas7Uvt
fq8Ksc+7QGFADF1RaAtejeZg0gjDYiuFTeJQ0mVEswS1/nxXbU5YzAzsp0xxr2bTJJDRiupGqH19
sh9LRZlujuqCYh5RIJR9EHfWYXyVBeQe8vhYnX6UVFdV8zfJL4IuGW1rjc7uci/YsXEjY5G9IJ5g
0QMQLIKlsF2Pn94E0Lc/LbB/Q8RXF0zNiMHtKRiZnW+tiec1Zn7x8TADCR5l//0szHVX6SE0GBFi
+XVIbPxWzQXWOKoSJF6+QmGkxwcJMgx/5G1Zm+ZICCp7LA2RCRitDCcHDhInhKbj5/qnZ6TMUw5f
tGWz71XWMHgXxKdYKobZkz9O/K0XtnMdiZnPdSTwcR88m9tuhXTVVoHI4XTHnbeHHkWW5K5taz5L
kT4e+JO7y1V7X9rx3X7b/jn3vTo7JEEEko61inO9hnhEyeNP1krhrD14wkII343hg1fqkaVdj8Pb
gDYNUzqp36FRsro4+w5zIlNx7P1H5QDgu2sWkOtrY8tezrTbXRh5Ox8w/bwmSfq+zZjqOO5Y4n8+
mKSry+m8PKDRpyG199k9CMZB5hxaW1jkYkcDw/7RiIrLW0cqXHPX35l4xnOu6QdOs0Oeq3SaiDOW
99szjlUda5DJTl7ECa2IT7mDbRFCxYKCKIHX5gH7r1RDVv8842exVqVm8B1uH4QhXde4SODiTh71
3x87Vp6D4dwj4SLA/xayM6TWwaLJlN/Xbg6dR8eS5k9wCmPrR0hPMJ4uc7n5pl/APhh61GqWoDzJ
AMb80k4BRNss5WETU2opKhQaxq2T46R3lU6OtOTMBcQu0CkyRC+qK7sGSYyZ5VPslsa/xmFa/X+0
VDsmFqg8AsN1oRPn3vQl63XtDkPCLvNLPZ1xootx7PlXGpeaLSweep/0wQQRhS9jPN5zbEdUrREm
yfwva16vQdiRr3+PM1aLMeA5GelOAfX8VL7DJAXbCeVznqOHVGAsFgQnc5u8mFk5seTBRaJ5Clxs
6019/UdnDKalUhPwlyak6nNu/EsBV3XI9ER7AkGRtpMPBmPqNgGivdzN+HhRCwTeW9wVhVjtiLC3
3Y9v4WoMTr821nLnY+etK/wplVvpYWBqRRq1ngtg/L3fzE7d0V2m7sSyaPOYE364onUsxJUd0mi/
/6MPkGyyk4QR0PgifzrIjAuJxn4qkwqyBscH+5GNjhzGFqhM6tKyb1EONvQ/R/hiwTSXGJmihrUI
vbvvTjFjjuAQgd8bkA6vzFdreF29xuTQFHc+hHwlmBmbxVARPGMvKPtU2dvo/tfsxKQZW6ZDN0s+
AzATv15ZVzadBgQvoPFROHsuXm4hmsfbQ9+WY6NPYpGDvQ7Ozubi9w2Lq/9LX1jIeB5LNXMCJYUV
z7XxCiWs+y8jm4ItIH1/gfUO4JR8xb3uA60QLuPshrVkTdp3axbszSlWpkhlPam3ioJ3E3Bjuajn
belyxxSv5yqbQCxM/Ug+MMihoiQ+VVJJ3vQJcIk6WgNVVBzriTeVqJUXdAScrj43mMVp3jnvjnU8
mKIXTAg6dERNRiuOqzmaeXs3USBEkVcqcBioAzdeIRDJ3ZKRqWmVQWU+EQEyO3MjhOySXrM7l0bS
7i4XKzbo/g+wTwYg5Frcrfvz21HvfBPrGrqbd1ILS6xeynv7DMIFEZnb4K+MCCR3sEnNnGNKYw/d
9NWaiXns4JexEp5xymai/87vxjENdMy+0k/KcHNKlmiiWK4sF7yYV+gtfTd5R8+LaSUTsqEOezPu
dJL1CPjySK7pYPzF8nLfi86PKk20h/XfXqaYdhUFzRDuMuJ2aYo7QvrP/+UgTEIBNINFhO7xvT61
p7KreT4RcyP3n2RNvriLLqa7iqAOnJaGCQVIXxGuSE7zJMdu0dI2dG/OSfjZQJ6jxomj+OOqzzRT
r0FVv3qow/ZW+0arqAT3dk9zU320xCLw1fSs9jrGGIpqvS81nDSeKO/6KDE12PDYEM2SjAIsnbFY
53bfTHBVCouC77q2pgW7wBA4H4LjSimZc379aapf0KnHnDoTVwdU1F4pkgQI7xQ+xqQ4rgQO5WxG
MFnWoxU1qyeIX49VCYBaYzKsA8iv3Q9C6+2LkLA1L/eBNL6gmHn+ST8hSJ7mw0H79z7Dx3DVN93w
AkmaAHtw6GZx5yFIGiwO+tx5aGHG61gkug4rTkkqAvarI+ATUrbUyhEO14/1uAUcFZ9HASQRXZuC
gHEnAW4fpSde6r0CkEgg9JIBOkfWyuxvLnVSTInBjoyXtdv7n11t9ZN8Egg7kDv1fxBvaQ1O9jDY
RmVHJunyM33r/bMUpQ6RTCCgzUZMNWD4vTM6tr8CRP75QNZFYafdw0oaJlR0OSVwBSkUvOJ/gcGm
6y7c6H34uuySSVIpt3JWbIskebpfcWclkQhJsg0lg105lrYP2lXtbQ7ZY6u0S6bLG5EB3CrBSHJ7
n/7wcCB3HPhsZ7AMhrlIuxE7OmT0LbFNKA7Yq4mwAVrULI3dtDMF39E/el1rYeu+SMpNtgizTpHx
UTmTiAqMG6G6Y5DQ9lckGEHEVT6Zys09yyLbbXSATDX+lIxLOh8VdzWnYFvAbEFszH7ZuFAUXzxB
BoAQB8fVWhqCFmoJUrMA1K81h3DBaePDRPaCLtvNqpaizwadk6gceHLWHfRvMRXzTe8fISRBwKsf
tgQSx8i/TQ8fGsBLLTxjOuMjbJ1eel1M2N0376wW8CihrfasZ6TfsxvTBBzHMVNvXvKT1G7URPnm
3HozTIMuR80rppkY8Wnvg0ePQ45oRpuvW4n7reDFBiiuOFMBtmt1wXlHg+BSh/YsBhQdXyiogyjz
CGkeSe3XwLlBe89St4gg5noaCiFB/NHP3ppPwm9B8p0PYyy43/AWfu+ulXO2suiIzLtIN/YT6E6Q
unyL5VkAVA5iDQh/o3vM1HPKA/rkVpiJprkLnE2Wg2X4t5blwonHH0ENnID1CL639FT84emUHb1R
3QzMu+mqYcwW9mqHQ3d41YiqU6GVYwONbA0+zBQyzlmhM+B8EENSH8lLuU983z9q/g2vNCN4NUaC
3FbCJDH6yaS321O1puvPTCRH9clfVDwUuSyZ1GWaj0pzY2nJ+r34V5xal1F4KgnovIhmfe8cBQYG
swMma+w4lV0NJrz0VyXFvFVRx2OFcbHmlyDn0GhAaaj2BT1EIk24E2slZ7iKSAiQjID6zeF0nT1N
cwU1CPG47T3Tk3OpmpDrWteJKaQvoHPlDF18UdYgucqDgjgy6yUD5dqTTTTm6EYFoIqM65Lq4zLs
QAk3hAGn/wce8FpH5ufL2B8VvgBDB5noNy79C3cCbPmOXTtQeaOckGTud9xCBpa+3p4MeFpb+dK+
hcs3gajothQm5vbXMoSLJzIgpzpG0hlzTWp2/2U7xbUqor3sbUslt3IHEBLAc9mBRqFJk7iEnwcr
w3SZrtNHDV6Ulf5+D846Kl8IhorZ53XdIJWw8yoo07jqxS5po0mgUgIxcSVs/VNrOdYL+iJ5m2Sb
eHMKIOhPyGp2fGB384AWGsxmzSAOXSgvVwom1YSojN75VtSCIe7nwKe7HlP72fx0R6jYRvGWVBxS
si/NFMQYDP2Mww2hioJrosJTD71tsLIDacob7cZHrvLY2NOvDOn2zg8EwfMZmzbEs3TlXPggKEga
tWvzOsrQf/tzEUL3DV5H1IUwJnYYpO5s1GQ3C+ENvd24aPjBKXVnP22/+vTBr1ei6Ndq/wzN0/M1
0swRV/Z4BEKTizWOocq3GxKUT/txPxIy4VoOW4Wbqn+XCT5PoXPKSVp914Vr02XxSx/7/S851dcQ
E6oIIjgJOFsjZZ6txhXCFOyiAIF24ZS+ztvYlt97itTS7JPWGYLAs8Tp0PDtn7NSonVXHHFZu8EF
bckmeURIdtNfwDtAcOmjmDfT+a7H9L25vqn5hL8EwwJVqX8N8usJobKzWV0QrPBz66A1ZGdQWbCj
yB+XhNcnNWCWP82b2XdDtD0VAjx01Hkb4hOR2ZedZO/n5e4SBYQeQeCHAeyIeKmQRxZ7ne2uuRnY
d9q3YT+AfCfHSEmSkVDNuWBGafb2MUYh6vzwTym0SpWcTC12A34YAVX3jfWjywMN3CIjjCC3txCo
+VmzeJp/3YNjxNzo+1yOHQUPie5EAHGa25GK6oSVGP4kVHqHlAv7tFQAXIkY+2moswdEMsrORsjl
tA6STdlKZdeh0s9gxNlNC2r2ZuGcoL4/JvZindyWUqb4em1KjgoFv9Ziz11F+lE+X35uXB++gAC2
Fx22/vcYWwUH615N27palHWX2pIh1B2nFkCYKBuG+CjG/q23lgDgJ4usb+kJcaffcjLe+OzlJOzT
AuIpZCi2vP8eh8RLlZXxPo+8zB6IQlumVuyL5teoV9uHYzMiO6u2MPqgdS2eH+9vi4Gyr7DngV+D
a98NTMYZrBGuRf1JKxT8eKp1VV4d6hhS4yxbOEKJAFSU/vwbqNsYYL991MXwud0FY03e6KHk+wJH
oExFqzfRGwLy+GNaqmgRg3WRx6iZDqYiuatNYG/G8zq73g0+Pag6MDyfv/G9eCaNN2hn9ovt2EQM
U7iBIQXi97FfVOYe4G6sbf+Obr9/MVq1eUIXS/5kafuKs5YJbjdfrjeveM2asv+NmKq+PtX4lzxc
EUQQFA3GOctcztU8my6cRSpteH3aGx/Be66Y01UOYG9oDBGlOXxZDZYYSmfD9opnEVfx3dLORv/3
0VhF3Uk9jT4mcCxZuLRtXvHroGfMywwRLVjmJ3HJcMg31VMXtEwD/7EsMAHyEn6bWmHxtYY1xcdU
dn+l1FBAwNniH/y3eztFMk4iHXGDpZRyxFUVqkE9SCIQi9jlsyo6SMPnrLU1FdpYRCifmaOR1Jyg
Dcm4GlPPQ/S1EJ4nsS2HoIIfiid9EKuxJmAmd73go0fL8EF8sMPEXT0PebBGDSJ6mr3EitOE5HmG
VmN76Bbwewop0nZzEOjeNGGssD5AOrxfZVQISYztxaRC2TLWhR4Z3YrsebhSY5u4+v9t7IuHA1QB
0rFekG3R9p9oNMXWPeyn6lOr9ZPLmO6T9LKMVXDTYlz63Kb+oyTbdTdol47J3wXpxoeUMpRyDdzG
JBxnU3Cd50gULf2kwvYQb84RzU50eRCyG1ceedp0hm+kBxnZzTbsXUV0eBEUdSTcwTb/ImlFkip2
oN9qPCc/TUlRV27O14vG9BtCeomqjqZkHJXKOz9OKW5e8sf//DpdXbIhpZ9JMV6kmU6tyVyx3H7s
pnXWsrlfq78YUxcJKz+kfact/FWg5b5XYde+EQLDOEU0jPXDHCmYPE/d2BZKTqvnx7txksaXMzfF
/VE0e/xf2eDhp0DO/N8NRssc5Yj4Evg9n2DzN4wfYSDucCHvJiqZ9ThPK/a/c9PT6H2Ulrs8ficN
HOCD6diacF42IwQsUEv3Ax1G6DufU6xftI+M2bG8zwQjsRT8YLTwzzWh3XFgFgOx3uiWCAVQbTIs
OwdYPEgKP+xwQ3vgC3hDzqLg60n49wCAMXafIjWXqqsImNEn4MasJIl0D6wfdS7tWehbgSHTCZSs
2EvxYEtIIfMabebBfbrGCWAVocT+6p62l62cuNeTABWRTa+W2UZIyvCa0c9Hh/odvGhg8oEw8hqr
YZe0cr6DRm1H8Roll1PplKKL8GSYOJI5pYZ0qtPddCZ7XvYsy7yu2mPfBXaKdRUU1FfEQGk5r9c0
fTvxW+jWmJIObs4TkdvaP0GMFC41m1Q9MSgqCwINg6+EwozCHCTJlAz+RYLzIhlkf22RwIJE2dKM
io3LevHX9tpZXkrFje2PMCOMh2pyRvhGIuTZxgnYDEpO5n9uIpoHiQXFitGyIftGYdgk82plNSw1
2DMSanU6LrONeulGtURd2xV6Cjxxx2239lTBlNyIXYWciOx2bhEeOBKff9xKcUP8T98YL0P1fo+R
Gg7CEMhj6p4NSqYG90CkV2mS9SUjLjNiUYECW/BT6oLAQvjoZZsrdxWFyFYzpDV7TDP5OwJzNTkD
y8VeGfoLgIR5Mh+7xvEC+y5SkvD6vtP4raza/oyEFW+kiBe4RPxmmq7nkksNqNEbD6C5gJxNBcJb
1pTLIhKXO7lqOwxPuIJNaj/zqqjqrinAmRfFwfhk3gWHii1pqwb6p8OkAYl6S01KTnokFbnGL/ct
FAHQ4byMSqtLCm9fyAAXSwFxqhBSPwMvKCC6omFRnhJB5M8gSeeKL3te1ahRLELbkD8JMgR603C1
J6B4RxvYVynWNwylfAx7niOPTAAy6FiI+LFswrqGOZLbYFZaDeOHjU36oa5K13/W7G+Q3wFWqnmI
b8Qqxqj4lIaXExeiHk8TRKOLiHfzMj9h5Ju+CUgQ7UK3MC/ObcEj/kLYN3cy6/n6CPgNHx7XDvw7
o0kpBDrIzaiMMxtYOgdM9NKgkjR5H7CekI+y7U26KBEyBOiVGAq2M3WoDbrwkbmLYLOjkGqycsRV
UGSZGKGoJQCLdYS5OPsB2qtjowHiBtSp7pxJCmKholP3I72Iuee1/IRJA0OU1yAN8wiQ3v+lqVYD
EdoAJg/Qe+pULj8JuKuyriIwoQwQTI53qk7Q8/WqaCNX/t8e6SKX0dYHmr2t9EPSHOKKE2NEZ7c+
PLrpTGOCDB5dArKkEU6P3rIKo37upX/Ipc73QvYpYAAzFg33EeKcX/rUCiufkyo910Vy/rTIh6D5
hwTTQSveH543KecCyrD2SWJdRTUOcpmOSIlFrWteIMTaIYB53QD2wFgNDfJwS24KecSX5s3XlCSp
KgyunJGKZ1guErI9BGmUDBABea6zl6hkAbU9LnHO33HJ3zemCjeM0BmzLv+XUzVq8yi+OYuN0c62
K7Elp2KSzw1CUT4jlW0csUYUAE7uI8/MwelVh7Xmz7hf4DcYWx3fsC2ZrXHqAMHN2y3D1ordx5ri
5TSRAJJf7GMEujtAG3TEyWzjiuyoBS42FUzDSqbsWOdUg2qFjwuo1w1z1x9IklVklE1FxLePPI0R
c294P1an6+dOelhiWbD4tG4RdzEhY4+ZMCBxw0Zf4vOR+XcfbDXUW7LXLOlUSOxmSkFjoJMcKDRK
aZXeb6fjxJZXT2X8q5Ilvzo5QdWvNvthEs1nT1DzZoZePEcXeqV/fxliwQejGCALsDlhHVAHiJcA
I73GoxDcC0YVOrRKEBpTJ32kx0T4kHyMOVdpbfHcnGVNO817b0ZbCaJGRuLIpdFrzal08S0Sh2fS
qbPE9c2QxTNxjvhWz/omkfKFMt9aAQZw0I4ilIVhMyWQbtOiZW4/BZReEwPyGfBVvGnmO/ZOHAKC
jKFXyGzkeE9ERXqOFNdXChZE4A0F6FFiR8FPrCF3eX+uzCcAvuAVMlDPBJBmrpqVFmhl0Olaz5v/
BBRpnStHx9M08Gq5XgAma800yEEtu0B2gukAIMOWQhA8YBGQJ0UXlJSBbHpdGqXj/mTHGtAEO6SF
lvUjhnbBqAo6MzdiOeEpbROIwqSE17rmXe+AcOCM4NZBNzTrcS2JiP46sqptV/h+5RavkuKjYYr6
ufdstHS8ontid1b6yUuFeMQk20uoy+ISaib92NDCDvPdFcvpYf5V+HN6IAs5UHkJqvL1txqloHD6
3pzXKrxqXqc0VlLdeShbiJHJMztBNOU6LahdUHUMUJpIit5EGjGpN09ljbnKPmy6UN4FZ47twCOB
c0R7G5CVve6t6ZNHBwLfk4dEGMSdWMee+w6Qrgg1H0IhaxJJBds9BK3F3MugOGwJdWFE2E397UlM
JF3okl6WNbd75TL+O7dwAD+R7HqtOnov/LDuhaKwTO5kngvC6BLfHkL73K/XObz/R8tnLhAiVjnM
HP8zfGkwS+iQSlmoO0kbfOHjzFa2NYK9k4miOzCzrQQ0RCAvhSc/NI9+EiLkp76iImZw5YUAIIwV
iYZv4I9quu3G8aZaePRYwILATwl20pA+QSECol0ZcmhdlINCANnvpk0fyeOpc9bToMBs2L+wjpY7
NZ12CbW42O6NJ5+T/MtfmJPHMPZoBT4I13EERPI1yAuusslCPlzFhDzMsFXmX3JcUenzYWK+n1YA
TpO5ZtOFPM1ctshfeSZfMQS3F8IQrDrKmlgn21wF70E/ImmUOOe4SEnoOY3fa8oTjfYZU9uCfzjs
8AfRq8vRYIDWVZbDVpfrG0/EI9JxBwBat9xRI4gox6WQ8g/5+ukFv9aRdulpZ3k9rEwZwW2U4QhQ
wcg/zlNAr9pP7gbP/2PBXvAjdOMQobNsadwdQdRFlk+OGAvIXo9tUXfO+uOkBwRwrlVFOX4Otwg5
cXUrnHyTUKvOM5g3WaKBqRNM99DvjwBLpBpXu43hRJ4MuHwHev22yjwnZQCG3EXAaiT6ggdqOg6l
HzqJMT3yxzfqSV1BGrQk80YmJpb7C1EZLRkwS9m2n0sbaoCuD+NESwipi1mXDESLoSlncd4rs/f3
xyTtb/WrzAOqc32vrbk93o1Mq79kL6KzA87E+IQnW6V+w6se6lKBfpGwvuWsfDEHV4Ef0L5hEvBt
MOFDXe/2f5QZKGet00bt0NfCpM+xF6RKT5SLfEzrmRnjWZeBBxtX7RlEodPAEX+0C7hscJLZG4bm
fgY5d3yvN9nNhD0uIa2Xcgk+uI2lFwY9HLQ3TJXbIj4nGYOc53fUj6DOrzvF3r0Y0tHrdTAkipTS
+UWfMALgLdzxKDz85hQts/qUWtVFemNWrnil7dPfJ9WZTM7EkWtUfTnJmqBeTgCXFL+0/3L3UgNq
Yz1iIw18w1P/wi487C0U442W3vRQChMmzXTTGdxW0LdmZyujXAFNlkwxhwoi6sq4d5cK2ta3Jgjv
TekPdE7JG5D15FV5s0rrWbFcDWJTKkf7QlBALf2CN831WC30c7JQY3M7ymofypad/Tj7cIUjutg2
q0K9eyqSAQ4rzPK3zPHiMYe/CHz2C2ElwUvYg3DkjaDGYzWUABlDcHsBFqaTL5Udfe4C7qYPRYSy
LmOZBU6rjrCxewVCPcqkJb0A5bL+U23TjkgWJphClpCE+9/vMjj8iD+idETvHdkZrIsSA0fHSFrL
R0esng+O59NMVvt4zQqJUa4dMWYA9dukTYnJvE3T8GP+FUMNNGAd5lJrTqPywA44nHXjEPbWHRdA
882eAj1aWm+1jsGkJIrweTdEXUzYgt0xGxFj+Hy89jSfojWKh3yVdCKc9qrygrB+JTtE3d61M/eh
Mq4kIv/Sbn4QNn4LvUdVCVskgD4piYclOo5yNNV3+nNdJMzdUXNn2dcw2g7EH+XhiJalRNIJWHpb
NyOKSq/Z+S9UcFh+KeUqdkX7xQd0QJhgobctsSRfyyhOMtme7N6rB/vwBFaygQf4+dxNrif/CHEB
YGyxSeA5qpPYOKzxH8//DyWEEe49gXjDSGDtYxur5NHrnBwPfBSZmg+ln57SM8i6u/yI3Kv4o0li
1KLyb85O0DzdkZfL9/JVVpHTi+/r3BB8JlhRGUPKE/T2NqNNCIgRx9BZ1xiCoeoqgwZv8QRE8HsZ
219Xw9k9sQlfvCZjZ1k95uh/c4u8Rxv0F9sXoyeMSniuPQcNTZXD/sSp33IwOUXiCnhoKrupw6I9
ByuWrvBnt8IHWzYSGFdv1r9Ai1fwj2OUxjjYZYOnZbS303gpCm+sTEy5pMd63HesyySX/Xogn6j/
C7M/JA5v5/QJzSarcvwYMKRIWK0u3fbmI6e0b7E1I4PpXYn2TKd5xQLiXgVLKeWGeenrLawlQejI
TJ5DwzOTIJGfJYSqRwCqkPeoVHzAXmVB4R4Cb9MRq+FgFzqtRETng/AMtO6kisgK9wW6cGjHcnDp
dEvvbAflbwPuxP9rwHJthRW+P0vnztG5cku46IsPtCAtW8yiSvr/iCJvy/WZ7eSNheVpiqosfLYL
ZnG0wuLvsTEK2gguC0J8326F0aEeNr5EvRUDdr5Tv4CduH3QFFTD5KFLr+pLF8QQwZSPwQ1ZPKQu
hOB4eHLY0y9ntdDI9PWVu433pCvOpMCZOlvg7vIm8ZK1MIn+0v3iOJVN0OEvtaFB5ZJTVimiRWP+
77B4Pqop9R3AabAS4xxO9IOqH+iPvq/3smPSE6MdPiuMe9qyx4rG10Xlne4DnQbL7eB8gWe2hlBW
g3abVjIt02VD5haX2NqddLC/RJjXUCMPwBixnZwkXZSI8C1I52Z0lN6hEfXiDFJ9w6on2hf3aHWp
LaxqTLAP/wWGiGqTsOUqo+I1cc9DuTDdA/gsjQw8GPYAMQLmIyxH5hQiybJ8gXVvbYp3LHy/71nY
uMQ9BzHk6WITNuqnUBloHtMVTdGUkSgJtU6Qq0zwGPkWUXyUp6JuHJ6nNmL+TRvTDwdyHFCuwoYY
oFGD114XbvwW4HHLcxiQCo+B8Ndqu5+beQguKz2bBCZDCgwWq9DRJEheaUBIce4jcsMokRWoSjo4
GXmadGPoFVtXJgd8B7sGrMWJqOhUKEqPA1dTYB7j4JXYqYKYsKyNS9YpBNqbikkPMoJ5FpEQvxMd
oNKbzkfl9hXzcBiBO6U4WmoCXWjNGY8hjyspFumFc4anPWnZFqT3eBfP3zfbLWZAmw4PT7okKfEY
k43GXxTEPnHDa2ZQqCWnOzZoYAXrPi0GzXMGkMe5pd7toBC4yOgj978I0iHak77sxEeI35DFPtZK
PX29GTIY/PZtBmJtIN8lyC5rqKFTN2r351zPI2VThMiBg8T5u+R0bRtVkCcVmFyMznMq30ogkTUr
3m8y0V3CgJVgmyKSlJL/+KV+K6zbRi4qoPbQYtorW1UgDk7l+zYtrxOC+yUHLqzlXESDJni2fmQY
A5p08XSm7Pj/mzU4kwCcQ9ki6k9+BkF3dmHVC5bMcQtSozox4ezTumpP7zxDA8z8jgyV1FRvRnsj
s0ziazKBhr1ENtdYA+JcomtjAyklJRshKM/Q6s4jtRGz+9FWP2ZqwcdL/diezU7qGPJ39hG0cnfR
Jh/6yWqysfiYqP5h54/buQdqOGhq6iZvBubmL88irZwAYNAqH/umGQ8n2bT8CgUMOmj/bvkJEJkv
UGutKOMZpbvBw+xRVATwK6RhLIRNusStv3f/bUTSN1SF45XyZf8IGXpqG96HDSHMvHcJnrYIac7p
cGqk4resi9M7E1ivR/k+WVwEpqiRv1Lt+kDX0xIxYLLA0fexNF0UvKywTMUw4KnEiebp0CyqXLmf
3qrPa3HpRGNUcFXPw86HPZjICufKub+/IYuLzQgIy8tJDbT9hIV6g5ZR1cHSaB4dz3xkbEceNzRP
RKRXkZsKdV4+yVtdDZQvvrfxKW8MQhGMCJhR+y5junJ0wYW4hkkPwWoUq8yNIlrpOUGHq4zDIdb7
vGR3OmfXn8ed2JK3LdKvm3x2+lnGhRKi8qYbybcHL7hgmZRUXnGAuHATnlcGO0nf/8C9MZL4COlv
oYHg9RgPOewFY5YjUjSdZq5lpQ3clPIGySZRLcuARuqaNVkBoGg7XDU4RyT4gZak9J1uTVF6g1ZB
TfPAZlMty+seGKddZ+agsXm3Msz1fOXSg+tjtmxhPZOlFEBQaaaJMEzAHNVEKgowTwFZ4P9oMMRz
+S9vdqmkwDOH7fPHjRBvkXzkIzN+nEAYIz6XnCdfiZ/64Kw9qJWVWwCWsFi7m7zjaDDZnuOWhU/q
ZmzyRm76URTvhOwoZp2QE/9RBFiS34MXXY+ATCKa/5UVp5dVqjOwv9+Z5Ei5Hg952o35hfX30oQX
XIY3KdW73VTbywH65boAJ//jJzytV4ejWRyO4RQNa7+GBJRAuz2PjVhmq3hUd0h7VB++kQ4/PRsr
z4pYtv8XXLE7RtKsgb1t7+70efL3btUoofOYyRq1E9UCoPFXFylOg08JMuyPlSPlWKqw6uZ/kYuo
UNfw3jn4TjpqVL7yXsTxcOe7vBFehLTPhlfXTKXgkRHeiT0UH2HrgeUBjqHQ4hG/zAmts7MK2F5V
Xj/QsXR5QzzVP8KO6kXkt1zuYSXV8WqNq2z0T7A/W8oXNixlQwJAKUWp9YOjo/3tX+pMMxdww5Ds
6tvdynhB1j2rXmR6bNw+4iFJVVFpJKeuxYZgKlvc9XavTmhqeB0TUfhKGlfAVSVDv7cqGgBMwTg0
nrN+qusSvq1Ok8o9uC0epWSZMFU2oL3YVCXXHaO0AuC5iRZtf2PSWLETnL6/3c/kkuGMXuOvfACH
Uz6LQyoXyfZ1dmonikk9Jw/hbzT3zuEZEHdbID7Ot18ZoVMyYLOTTEEWVr3baFOz5wv7FOlEDB26
DNuRJ0wn/+11KgGDyOTmisbLgHANa1wXjJKxOe4SHkRCXnC600TPI+LRQfpf3bdx2SoIMVuVPqCc
6XneFHlOgzzTBuZV6Fe756SV9O4Eh1036MTbaEzE1+D1aWw+IPy2R/jus25QkxBJ4uvaJgFsMNUi
EPOaWrZWUIJafEMTvVtSLfXI66ZO0IcEc0gql6tKm47Y/ShJwVO9cK5p1zf3z7YVaPIU/5NvGM+K
IAxPv43VLpFL2yTcCRrp8vbS9O1OUFI6PK0bHwdrJCpg5oNm1DwiEI+F0GkuGavfjeOqHPnmXBJg
5f3whKZRVAfFSsrETymEYZAW/kJhdpRn+Z2b5U2mFeeurfHuClI0bbcsdGL3588LrXMolb4DA1UW
wotPfCKdJJOlQjWvKyn6W9ydilOL6Gtg1gWc8naWOr1E8sX85+IJPwkgzXL1O3/G8nmANRutZsm/
yNPfHLdk0FGQA0/VXP/H8sg9eZVf7F33ATAjxi0MCvmT1VtBsr3qgJ5Lj2mTu6J3yKe2G5k3E0/N
vZEPTSJrH7/iSS8iLtYkuaSHHPryUUBpYvPUT16Sfkk+1wAyo0ahsWtGWlIfOwNFslx+e+bKjqby
iJ69kSVhhqqJHOSHBxd3vNeJfQA9s9EL6aRRSWPpbB7NZQfs452OSaR/4/5EwyfCshPRpdJTa2g7
KLyhQelhtE59Lz2I2nY/qPCHjJEsneKP5mbMr3NwYdyhM0ovsMAQ4HsIeIXgpB88eVI5gUIcANCS
9044x5UCCWBb/+raYR57GeIUqPaUkIQJhcKkBcH3MTv7NlNoaXvX1agif5hxlQEjLdcrZcJh/Hzf
82DQ6fzDFNCLBOOwAvu2HDkFEC11TY4XIpYCMtd67TvYOTHUy7b6qYoMV7gHG/MitOSKpmVb4QYi
3fP48Sy/tzpewyS//C3Elf1XSien9UAspn7rA1clYIX2n+sh/dK/wYrIY3LilMee9P+ZnGz6EJpT
dF6kJQl2V81x6LfuK5LicPqbBE+lZ5ZV0vzg0PmQR9G2VMxVmZzDbc/9TlPiDUUVmr2zA44jmpGG
Xu9upFy4lSGh+zV5rTXyKzLLENkY86whid9FOA2tvUJ9iSpKrjQ0qhJvaLHUjdhIY3FY51UQ7qne
z2OfnE5vwP4jc1HqtCe8G+lV98exqS2PsApKOP+fmd4k5l7FVL41hjSX40Gz5EkZNZzs7ipbilb0
sGIb6CvCMs28W0uQs6ZVFgH1anfcMYXBpqEdduoFP5maP6XLFj/IK2pMz7XjGgRVea1NqRDFllj6
0HbIKdk3oJMN0sbd5wcBggCSg+b+14T+jvwduJm/Hmna44hxOShWfT24Jm/BE4BVMywp20DeHYtf
BdRoWeI+HB/wGlfmZACnELHzoUvPmFQVmn4BLAf9CzB8o9+qH+ubumhYDpZxPdzTbtCg5vjA6ZJU
U3bbqzpCjseS01wqIq6GiEgqc5YF2ZxMNQFgxk5TA86BXzP2Om2Yx9ArUCsNZQnxCjCyTomZdk01
GwRT6S3wmBdZpNuo9W5S4wt60586S0Htn81e7BuT/XEeOKh7dTSBhAuJjqMdxNGrqcp4YpSMDhX0
Eru+895Pq4FbIpkV+NTNZBDg+ob9i2JPHsks0RCdzDtNxTF5HOdec6uvT55fIkNdUKDK8k/toBbU
OhWlnFSZgb+SdYeHw/nTV2DFbbumMD4xLM8/rKxkyZtUvziEMZ4yYcmRCIjnsrCBBlS8OMzqviSa
c51iVCBSlD8di++Ozws0QumiWVHd5ypdzQe0I+aBs31+Dzr8m+Ur4vavMDVXNRbPDJNDbqlgrNE9
YWwSsBWeBF8f8KjqA0FyqFLVbSYYslAMCgoBsJPZJFtm/1apFATGMBZwHcNjymYQgFiM+un/AE2G
IRGFOT4aQaX936Czyse48jQ828/UL2KyPQmF4My7EX806ffygO0EkCTTBBKntpOLX2LkeRMJBAjg
DDj3WGgYr6bM2XGC1LTnTx7VkARIJN/3hJ7Rl6sxxAyG89vyXTUCsn9pcZ4rV+lWV5B7s0cuohdn
XcX1M/REVyOqVwFe3Slp0H+AtCMA2LAjkF9FJt6tkbK4gS2VtpB2M8bs6Jg8hZxILxR+nS4XVjI3
suET8NPKzj3njc9R+25uclt2Rlyt9Q6We2XzQVbWRN/IJskcumVR9kJ58b6QAFJ6lWtH2qi+Ku79
zFDuIyxY3XNigKnrBMYvEUUd/RH+CHhWqXaTEQ8RYIYZPrErlVq2+E/srQagzQGYAd4ffQBSJzdB
oG/TB0VMIP94VAYXQbq1+UY1devUYlnc3vo6sQVwwuEd3ATuLFj7CAV16AkGwiXl7bqoDi6T7dOa
J3BSrnt/nWzWa8ueGTitR4Wfs9FGd2P3f9U/JPNwfgwDgRlXR5RXrBobhu+HfO5xrdMtCyLOxhO7
nTqVCs6sAZIBDgv2TXFWy4fhHXShd9cB3NOg4xF2msy+oTu4eDwznjn+hxxLp1DLF9gUjRyBkwI0
2JpDMlk5JWuKPxWYeJQuZ92ufvctf3KfguARHsvMkBMQwmxhE4ujZkAYgSMMhoC34D05img/BMZD
6tzlMl3xg9XfAQKs6u10oJx1jR3KUQIGJtQFjf25R+wrdWcpxvut42JN+66LDWyfpVXjg0FyaqsS
wsNoGNVPtdohp92s61zxk71MnBnufKZnTtvu/axnf9rAeZ71txNqxh9nCUBWyd28q2tW0HmjK3eV
fVkISNqyHv7WoFvJCInEUVwVeVzOHfeJGLTzYAlj6Kf7VMzSoH2hSN4a5l7GhKiuQwscIMuDpdjH
9tGMP+G2A4z/gWHcGw7Zufsj6MrISoHDjpmPDYsBZCPxzzaTs34a7UBSBzIhFvyPfctAmD5OmAIs
6ZsGXxyq1UFc1LOplmQsrkl64O+t4wL5QxLwqX11qQjWm1eCJkEqJ3bm+pveClf2neS8mUWvuxkG
N0a1a2GFHZdmphvgmnGGNnvxPOrlYNc3Ej6II67v41sRK3qARE3TgV1JXgQFX5BmqwGg8TK6aa1B
v+IVTa3ry1FGSZhC48ifFRIojiiz83eudmuSnnGt2vYZEb8fuT9R3o07tALCn6vBJuqJTf8XMzDE
/1RPP9KulhjHT8ER/UEHOF/I1Cn4vVnoOffJG4L0CGpFK4no2D+VbalvWu94q5UbHsf/bLSo1byp
ZZhwhph6HFUxgfSeQRFkpJB3+pUkCNB1kNOt7cV/JL/WUH6h6pZSbxUFDtSD3n+IQd23syB3yiJu
fo9uSmDubtsVKbiTl/NpQNtBZniFQDqXpRq+vbjr07G9lZqilL5QJJ1XIpQVSRQUyp7jotQZtoVt
5B+Dbobvubj2/9urrRfLQhNZbRNLjlmgm+wU29SZ1qTeEE9brU0k4UgVwEzNUqttMQKrdfT4+yyW
kzPwaMuBuslB6Aro8VpOmw3EMmBC9zX7RUfDs8UnbN+1HsAAJcPaFdnrKQrz/REzO00lVg1ED6sY
OnDXokThrap148yyOhA+sHsaM2rlMhf+fnIq56aZVcd8zlrYxPLViGq3fVXVCkcJyUAKrdVyvtNF
+O7CQnGzfMMfhDjBABC+3io0KOQXXw+uSTSfF5tQP3x+b+3ap77ILQinUA67aCwCVH89sSF5nER7
56WSImcr7Qaf+9OaARuj/+INSh16H6hO0S1gSKxRL+TLLhJ0J2ZtQAGC1w6vUzG8sB6TLJXRjQrx
gF13CtnosiG2683Kc9hi0DkLo8N9sn63stkLez2mQxP0+c+Y1E5737+nNVOWfBg9e0Xiaiyd+dK8
QOfTSrrWYj5VH7EPDcmR9kY0m96l/kvLcDkGWWR44O1R+T+MH8cc/WzczcCeUA+8H4KXwtZU9r40
qjb7S55+tw6gYZ2fWeFhFkSXMxh5xi2GA5PLsSSslBucEgOd2LQR0Ya7u5synaNTFnINw/avQyau
FBIpXN9EHPtxFy8550deyzxzmyZSa080jBqirAAT+FjYq5BTjqfIhJ/1pyWqoYQvU+FZY8ixJI3G
xyKVwjYa7clxQcUsupQ+gcrGB+6FYLcbJ8sYvqP0DYUVMb6GNtVSoVvz7NpCzlXO5W6Us4+c5cPs
YqgdSP+dI5xpLfGvwnrlC8WsQko1zhPGEy16XvCbZANq/Cn+IOMYyctfpX7VxCr4nK5qkb2WwKF9
kHfwpxXke1DyIFC2NVWWTAjNzGGsIjsN60vgexPgj0TKumV0BSruVC8Wx5YNU35aY29xgCjj/YrA
UkQXHyBaUMtiUVS5WePmGzBaOkgtINcvPb6JxeLL4HTl48rtXfg8ZMEorkaKBiO5DI9WEwR/cklz
nEWU/SiINBM+NUbc9NVphzts+GqlhzC/J+3ynb0ZQdBAkGSJzb9dtnJTmj7D3gSxIhggwDTG8DIv
37gTajKbZYMn4Bre9pAMJOl1SfPTF3ZftO6/zaO8JS0Pa24FQ8XDosrNAHYJsmu9SnBv9yDd9u8m
6vUbUd5SugnY/D2iDbtvxUUhueJIEAfvSdljCfoxgNCIoUixU03+f8MjeBizqmK+QtZnwLIy4gDv
riNKS242Xp5CvQ7toPN87FAx5INHpn4/3t02p8IN793s3BHiUUDIvvFQ7uPWA9zyG/mP7Un8QLyk
HGMMzYNaFcRYVH+A4ajURaHXkwoGDgoDnU0ToOYWQR2+pVRjmRIs5qC9WeeQfWxO0qkBiu+7jBz1
gy5fYSWj9jLWInyx/nOreXHBtCvZ6AaYPEFCVrPqWhufaWCTOEzsVdtsTMojhpvOYWLVMwxdYr4c
purZtoazc0yysQXMPF1jFrVA02L/MriB2K6wAG3V+rNil/aOcDW1HaCA6KGYV6rVLngdrHieragk
vIGGsXKLEj7I5FMEoOPzXf6Lt19C4ujplH5iPSFwQwSj+8mNCCteguujZgrHqjHcus0hcVIAyX7X
0xiXXOBT75uKW4CyqcdmysAvBHhOI7WsQ1SsGYwlvIsxI+do00QQGrLKZYuSEWsPvazYXJlcQCtA
Pr6w0VuaCgHZOgXJPsqlkig2radurae2pR0YGVgmIFulaPEWPD9JBGxzwL0+6Cocj18yQwiKTks0
rgk6ZQ5oVN/sSASkpobtdZyupfvQiPulfPjzqStpw21JZWCGiujp+MolStdpry/x5/JEXOP5Lo2D
9y+/+vXKaSon3tuuWIFW4PN6wCJEeOLutmB67h7lxYyLLTAVzLuE/GA3aRalyvT2uiCobgDM9fRq
Eo4Nra1sAvlcuiVbWJeDejOwuq0Eyu+Y0U5SU3rsjI8hgWyi8WI2IT2/dBLX57d0XKjJnZJ+e1+Y
B1fEnLBAsALfjM56Kp20vyrl2f6NkA1qmhZhze7v6TvOUYHjOb9IwajOTovyPU4tyBXtHJ0fu5+h
vNruxLB51sSXbZqcN6yyGHU1G3biq/0yaGkwBc/O9qu3pp5SMyCgbjVkn6a/Xy8N5l/1hCdaHdLw
HXqNL/4eGp8zRrUqSH1OR0lJDYmv0cqWH2n5a0LFLaRPS06GDYjxoseMJ9zolsT1GrHlf/KySlA9
OXcbpPQzXAIVBtmL3nU6b3BSyP3/LoB+Yvz8PgKhlM+yck0oJV8zIYsj1JDvBnaySWztRF25gwPB
MnvqgGQ2Pm1rk9JcvRQbVqmS0VZxRNmTRvl1VLMP2ivJ703VI35Z+MQdJpjGCJh+PiBiqYB1670Y
Qg5nj9bjYxRF058Q0JKJcnIPpjPEeNz3Yb8ITKEbzn3ofLTPBIYQprFWYyhHe7iCPClH76FJnj0k
u1S48197BMV2kfvkSQMV+ESaCTDT23vqDjiOjWkm+OhkRuHmmM9IX/h/vBAecyehJQtLq3vEih65
po4s8K6kCp1FcZ3lvkrSZR0dZIuxKroY27eyFXzE3WeiBQ9cqDYb6Uu/ubuo2wIx3mcpOq/iyQSI
Ye6FPt+3FkpvRbJyRWfk3gy9m9bLlLdx6sre8mjOT+eqiCqjueyWDjNyEAJ5CzXcNdbiOnIqKZbl
NK6bD9EvHHCdmheOjCQ1Wkn6wWDdtVmd+c4OG4wJI6yi6GbIXrdsOPHO5ZKjj+zH7lEox6EeUyCu
TyzZYKw+pVjWCghDB90MeaNpZbCTWQPm5WdSZ1PnfxdiSY/YuF/a8wcBgBAzUdeT3IkVjde3ZHs0
IxjOfd1CB1up1cY9R2YihWLGgeslhxfnGJKxXqu8iE4D6taD92VeIo9TGsrtd6HrmnYypcO2E/t+
MyNtUpapdlq4Qm0tRaJAHiejXV8redJ++glqZSzr6i153K5w4ZBvQ8oqLJM6HTHPkw1zNZQxDaYX
wJN/PGZt4Ko0Rq8xagh3HpmJ4jKdDAIddEvwICRq65XvFFf7aOw3NImIfyA7BTuzi/kvf3LjjUjo
rERdxf6rszWLmXSZQPtuv2lzLbrb4w/KSqVUecGKM9yL9u40iKyheP5+P0miJmWWjV+QzsnUi7s7
ZYYppXDwy4sRFIUl2sow5rnFLk9mRmAHKjqbTs0K5xBgaZ5wiyDpmQ8aykVNQI/1t0H/zEhNGLVV
k1ldddCvzQ5oVP4TNcARqV36X8jj7tFGNAYHnbVlJEGnXYWieeVHIVqGQpmopVjQBQg3BeY7ca9b
oigZfvjiW43NAd8opdASdWXAGAR2nIq1IzO9wv0iBKh8GvR6agWth6OVfBXE1ZupTjT8VGQ7E6AN
mJKhcUS9jCLBG3dVBgP4KcJaFnxaU9otOAhR0YUmjB7AMAgmpw/L11L2ys+Dw671l7rZ5uAbTTpE
lBs4GNFvJLzaTA//Stf7t7ulK6XVxoHjEPeaxdYjsuCBqYsgZTzOz1ZRz7cTpUayfxjMM5shxdHU
64I3VHoK4i7LwMWx5cfzqMuYemU2qmSUUqnLneLuug/X//AccntYmqGAoXqKBCmOKFjVYbun/N56
6r/qksyNh60ArffbE92oDgexVi9/AgQpIENk6WfxG0ojdG01QOK+MnhYlWZh6nwAKywNJo7TAf0w
1FnnUjg4MPUsbYxoXaEfUq6bTddkrTXWOBIVYCZQe6k2eVuDTY4NXpbTPrtFETUBUO4IGGAhA9yI
FPS17t7fp3Lk7OMcFh46Xion0xWgKUb0GimPDCPCX4CO9MDVSs6DoNR7ShtUGTn7W14vRXfs4WZI
+fz5ly2dShMo/3m/l4X4bNkYuLVP7egvTNw0wUSWWaRlgaBzkDSSUkune8jUU6/OTxUGfCtf1Lit
hMYw3rbJO+M5rXqR7lTN1fAYBvLP/b53uzUky7N5Blh3q+nJFnbxbMg0huBGq7WGjuuUZtCZzIMw
8JC6CcEBIzraRRpuXsEFnwOBWSI2gMwCNAdATvzb5Dk95qdBy9Iq0mJEawHJnek4quDDAuY+/7yu
sMQy4FC99jkXUP5/9AsiFl/dS1/Xb1ujnRvfA+G4wnCn1xnzx3550nzxS4nWTnJEYVbAj5M2GjhK
ET5M7thRAg0wXUY13ZSlRQl3bS09C2Argmz2qijVDvOzjemb0iaDYvSrS7Qt1+Y1a8iG7d5Qi52J
fV1N3JfqgbPsCJDn92ljyFpas9A5JVAJMR9W+auSenCGpd/ZdrAN2JOEZTJkG92KpX4m/B4iOf1O
KZeBHUb4k3q1gqVj+UBms7DoiNToElY5Cc3kKGuWY74EcW9L2SIojDnMPtCPWoBz3fMyrpsOOq37
0ZHa2XX/b5RAht/O7J1J9iFyD9dLgFXAouaCNIfe7vD4lROmXF6jIBlQ3y/Jp0HYwcssZn/VWBP4
6nscG5FOsAriqWHqOIr0VgvKRa1EXkOKSt1zGVi4LiqVbfk+GA+B3hE7pdYpegV1JcDSV/7ZPttY
MZEp5Ml1wEVPb6xr0eBXOwls06IsL8Morrb6ERxYe+aRuyfl8d9mTKJ3TnqaD3SjMVCUXIqmDqi0
kh2wkL3Ox1jZGDyrEMy1ED8Q3EkyS1ASsziuJ7ZNGz18o5Q0wCxsCFxTGuakfj6CTal33ilwKixW
KjdjvOn5oN7GJf4ONP673OEshvirwxTsRoTL/YOxrf85n1THeIPI2bqAQBw1AWZsgdeHA0y4gg4L
eRzIOZS9dOtTdoa2AOAbRLlA7ADgdcVhwgXVdMY801U2TSoHTwkpYHWIWpoBD1BuMN5aOvqtfnzT
G9oSIvHiKDXx6YoPC7yGn4HbZM/Qf4MNFc9f5ocZud4uZqEMmH9Aut629nmSLfvnZA7l9dcHVOcc
3yRX/waN58+b/XSyFqa3lJDTqU+GEF7VECAYeCm8rvii2KK8CXAnYovPxJ016mhni3xeVOWnTqH6
quArQ6XnHBhnMS3crJgfOz/aNXQQxnOmaGIQ4fl1dA7Gsb/igMCtEY0wYPm4dW6V690NzHefZGij
gliLUluqpdnCD/bV+cgan8mgdPqoWT/MAqS9bCjqTMixsKZr9TgwGiJFKpC/mhlt/67Wayc0Kh0v
M+e+0YJJyYDZZ5uTvS6J3Olkl+BF9vNPPQRHBUBxyIDtfJhO3QHViWVFlGiCrVaHjK/ggbATMqxY
Aj4uqd4w6G7teZe+LiNJQ7mG/zdXXNAgJfnT8XpdFj4s8AO/CMVp6bKu/aqhmrcn8pQ93dtEg0eL
9iOXNqBlU4uxmrlHOXSS0negWD1kHOlHjmI3EFYXCMW3yzP+3Dqrkb+qqO9gMgLCQ/G+ZOQHVxh+
Omv29c9dPP4loqnFHhOAMByYWARY43Ktuab22Fe5/x6d0FumMN8J3MIkm6IjgBxomZiqcpK6eAq8
L6BJ4gBhUr49xfnZuMpRVCQbHH6po/+kXg37A7/K892vwZnRiS2+fCG9zw3Fq59qXa+ayJjmXb39
6JO5YokKSACZpl2KjQOAZkkljObgjpJQSI7dqY/C0RlSjsb3rgZ/+QOhT5gmKU+WJQV6lTX7wtN2
8F5TDVmXdqaSjYtoyyKR/kFg0GRxVPJm+i+I09SJ3Of3KmRh7iADoiA7cth33pRPPvvrLDI7WE27
80U+6EeRXBdzKv9vvbfHd/ll17zjuStbRUw9KK7hTFIUwXxbJqhun6+Jm4KC/afFg6wFy3MsMKN6
Kavqg9ldyjxVze2GW4zMA4xSYZcagrf7kt9/FGTt7SjWN7lGrIRMxgbdxOCKVKhmNX+LsRhpj/Er
t34Xn7LASM/VAp1NhkijUG0KS39hEJGMnhgAk/eJmpLUzL5mOWJ/GvvUcjyIFMTkLyhy6BEkQPmi
WyR1rG4UUGJFuaYgnWWxCsma7Yip2GjIQAEo0JTupa26NpKJDujQCFJ9+rp0OZtTQDkNaR9aw9Z8
RHbbrYhg/33mTXfYHlokqMLb+rrVvbxL2omRB5V9FFinTeLu17RauSQrmZ+c6ikMABQa2ZDdxWVG
DWk1KOfZ1ktnoXwy+AWO5eybstUJSR2gCzWkkWiFDmtI/b1SI70L9N+ghG5/f7VFna1XkDnrMVUG
DCn0Y0C+6lS/kqhJJDC/Fv1nJATjkg0sHJea59kZn5BSW0wQoOSCqqNl5yMuhwlDYj4Jbr+3iUL/
ilk8WsWqhyrIrucNXRFdIgwUWpc5ucQvy1CezdVKKTa5301cH9R+8Rjy26TROdHnV9T4QBBk2/ib
TocGUzWV4mZW1dhl/ntqInbBhN4PQVxlo3b2yMUbXkD2mLVEXR72reZDpGNMvsjTf1qxM7WODSxm
CkGjQXD+lc1hM0xehZfRkmqU173aLDqQwx/SZtW7fsqnnEQZ4wMyhnnIZhJxtcmO3LfEC2/zPtaz
v4DfxPUwOaSvEa58id+Tv90/cdw127Zcvl26p6fuEqqT9dDjDaLIDl838kSRVqiK30ha/cUYshzA
avSv6xcQxcHpJ65MtTb89jqQAvX4QnyvKNTl53bEhXPtv2VZw378tNXmY884XE0Jax8LuHITSBZs
Hmg42fV45qdrBqJo2hzI1kdTQjbnfrY8gawjXZRs6PtygoXz0SF2T8GFzfHqSFiF2695uhqR5r/0
WUPAQcAgbnA+fG47zwvB4TrI38v5HKs8x74fJWBS2IxmKzoqL9xRzfhlanujDSDnKhxHuMBLrtS6
IN4kbYPZdxBMkAkCZf843NKWrDO2CUaW/FP7B5IQpNibOVyZ+SNoWbAk/8HogJ7jEIpiWHQsEOC7
7YpM27bk8Pnj6hMu6LY7vgzGqb99CU3WmlJHxMIkdAgnsoMZ4jPqzFJmZKCU5lUM7gyXxQ2Y3VNy
bLLRJ1QbP2LbbVU+r5Nf0qhAHLFe+wIrUx8qD3N9jvURqUopZ/JRwlmCDPQa4Rb0GS835RdTcNVR
WX0nRHD05mznXsTpZMxqUX+cfog6wmfYAH+koEL2Jx6tvp9TouJkCw8EgAtdTRJsJFw2sgKVoikx
FCR8arfXY++WrksWPJ5wfqyH9Q+lPgtkcZbSrFXGbXMrK0wk4OvYmghUYhfXURn6/5NwMZ58hZAb
9+v2Ft7HPmCXT0A/7+73mH93fqq0fWYzotr2zvrh3fNVg4y56p+pg97JCzvrVxHYccDUGx039NvD
jt5DFkRF5KmMbpV+Ks+mQjVq2p4ndmjcL8U7MDzKbdluKxOkOAySmZLsCg9mObIEb2LtwFuh+2WB
XdOY/om6NqOiJmUTbIEYZ+OAkBkpVZUBP55Als20s623aPNH09OmCdkHf3fvJx8AKsZo19wWs9+C
h1ZBuIaHjF9GS2/Bhx4AYMHGEWll9SPXlcTPkJnLfEGrU4PJulw4eKjTyXy/Soi2GfSg7oUv/DGh
sBUjYa8HZ6EzYGHHr6blPt0DOzgf498Dlkxob6NII0E/2JTeqNoRo4fYcBYFHnZl8kg6g8G8HSpC
/JDpjnGf9kkJA+laDdCqF5u9G8VN97FdWiDCtkkzcgufZVFal2L15jTxjgFdpYxGpKvt1wa3cPpk
fRDlS+jgy9PMsuaMdovYCZ8ihsL2d90CYjzQPVY2Ohl6Et2SP1qzs1ckSqwr8daSU++urGSBA7yH
Oal6e5DwPwAEmYL0gnEQuGtn0NXoBEQYSxmdLCZzP5YtTetrENVJRjlBelY05raUdq7QYuDE1NjU
FFomr6L5/JZM1iEI5msCaW9LAZvpNXHPBYxB0VQAnEwODn1SnVARecdATELPf0diAZbypMPjzmqP
pA2OwfdlNpAReqQtTSOBIOQZ0bSEqZ6EaOjQbN14oHIn+fMVCshUiqtE40Jl015Tt2fuFzQb2BUL
R+yV4MV97qCJXI7agq0j/GJYOwwwLYR73x3BfuIdW8p+3ZtfLbdd+IoEwG32SshUsA8TTNKdC8gz
J3fl4NnpnYh4eN8WYg9Ti8zWlZQaJO9jlHflwqwbIntehiPvSsvBf/vIETzP5p2bmEB6P01BPifb
7b7HgZVbmIoXRnzML+FUfPBdBqr0sT6R5tuy6YOcjkq5w0MezfzuQVmA8elq0OO9Xh0L1or5d8oa
M8EzIE0idAgPVXGaISlZ7IArZGTOcaFytVJZ5RA79iLU4EeL787tnRJgIg9feec53jlJDA3jx5qz
Wafi6Nx3ojtJ5SCYg7OtoAb497X4GCaBqks4SxwR+1JmTwqL3bcDcF4J9kHlNz87nl+S/CmopmeR
bmDOvdj3HF5OsT646dCR5zOkJE7JwCIFNYaTPYAbqx3p+F0rxeGqFVPDwV/nRP2pIX9Av9JTmKEt
PcWXStnJPYpfAi9OK/UqvBkf/cj9TwfkmlMPInwOnfwxAc9AG2M1HJm48sl1VVF8e04wI3dnqAfI
VD5cPuNzX/2IPh8lr8Dwo5pYhMKevFRvEdLBoHJLlrVWsEHMcz2eHVpGAw0dFO+t+AsWvlFr1MjF
xXZEVMXoFMBPK/TOZH05jFZ2mM/uuYjUtxbNk45fYzVmXJMQI+qgjuk/mSw8xAYrw0DfxZTMezcF
F9x4y6ZNbjBW23B2VnzlXz9FKJJwg0+cvu1F8lO1pxdrP2xhmWRamay7lqhhSUiRAvHc/C9NLC8J
Xlobi/gCTUu2x7YAxoVM6Jq0GSIjzzbI63n8AHtCx3gV4ccdjBxHWA+vUatAxdKhCo8D+fp2ZDcf
8f7/8PGVEJ3AeU4qY1g7dttcTjQyLlaYf8CeezU9jqTZNJqgnPYcJlbc4qXthiKOM4CYddxvftYQ
fMNWC7eYj9QyRP16BKkl3oUBW1MlPiqtBusSmcLTC80bE6LjTSyjsr82XVAsUe7Z/KcgSHr37Nl4
pKTtQf6GkuGzQ+3HTT13V1DnAFGEq1mVRPq3cb9/ZpQPmPLBLnXv/gDUeP2R2uSsYjjW1m4xh2V8
gtX90ZWIZmj92xIpM1synUZ2BKSz0naLnohUAg2T4cmDfjTFzs2bBG3M9oPzrBfw7DKPOBbnyeCi
8KcJ09/UQBnnH2Q0bY8rZaXuAYERHuv7Hv2zSMx59+74jsOicD1TLe0bhcdp9Hlw4FLQx0CcwDuG
7B00lOvCfzyk6OJQEdPct2+7M5kFsXvfeqXSdXVbAHfRHgNNiunLrZl2vJozjvEdU/X/xlMBhhJ/
luTx+IawtjYEl7I5smVRVht7Fpn3eD9bnbWEvgR+OlTeDgBHUbFoAkrn1Jj0z7h4spkloVTJ4Us0
r9m9VeMjYlXy0/18XHLbCfkDLhOXZbAP96V/r+fv5BkoUHtZxn55cqMJVOYfOQYHSP3Kaw6VL+ex
ts+U86+CdBH3PgqxZod6t6u/BRHTQjLJyDKAlN1TIAcw3571bibFIpAUAwTLTghG6nFLH4OV0pS4
KwGx4994xUgzbpoCXi1t8im+LGsC5MzYg6jfOd581GBCwqeuCSCvZRT7cz79C/H4yBmsnQc5seE6
ExRLw7BAH2zuCWxfaRwYLS/XmWNjGqyYeNpw4XAOjKGaTneP2l4BwnZt7CVRSYtHDA3lzJyL+EUF
HCNUc1idpU4pmQ8TXiATDJrkjizGwkISlrqH9X6AZboTCpm3JLgsYQCIZhMBa3pzZXs9chQRGyQR
8VttjG/LHNNGjXwRggNHQmVLw4xvyizavI+JdMe8GBesEkPwKjX6D5dzw/Fk3n5foVLVv3Xv8YQ0
CVGCVgxQBwe/WW8diN7VArljwJ8FuVGRtoI/ee/8r0RQYOJNjIS2wUJr7nnvwRctKkaZeNDfmPV+
hnXut+S8UHeZhZF+wQOYNbETYw9opldPs7zGoYqOID461pCLA33sRS2f0oCyidkivlxdPd5NyKyz
iGyu52AegDXAnnDMoNc4IBj9qZ7heAzYM+1YdekJeZmrXuWIE7FcldrMlEBslI23oNaOOZsBsTpA
bH1IGVpxz+uh6QxSKRY6ujDKShP5LrHN/yEK7yK6jejo3w49AfQEi57Vh8vohvVXYBy7X2UOMWl3
I7KtjSW97JnvVooygVQdEpl07A0DDozLOy3QaDA0tNsrkQwBgPw6k8/PgrjNLxQs3OMTkbghDCOA
MmTn1AjCYtubJKk5j5e4Rd9gP3AawGWMHSvcMhw7S1Wm0U66SuzXw7HKerBMEDwiZFkShTZxQ7Jd
yr1wJNhWQaerRwgkHLAf8xLtCE1wX+OO5qO/nM7qnqcy81hoUyGJ/OhO0/hFC6gDV8DS/rKHOigS
Sv3zBZbBqBWVf+YgHZylKeJJ4FUyI4TAa6ruXT1FtCC/SjeXL3A3iCzol5xcIxYzgvgv7tCfaWFo
Z+1+6lW5ZA3t/nWv1hKjpo5IDQc8eqYJ7m8jPrAVktG4oSbky4Ja/Z7t8OnIgmTCteKagut2ApYp
ACGSGJwMb9t+OyeyFGeMw3MVpme+NFb8MpGBljHST0K1H7AJin6uFgLvn8UCYRcoUlRWm5Oky6Kj
veT8/xMvyQ6vIu5XT8iJuYLfeqf68kkeLzg8+ZtNnfTrn+gWKtybi78sCdaN9LwJ2mQQxwcRd/W2
BSIUEkiLFfAGDuHFqbystpT4L2Yg9Yg8Bnnat6V5d1OjwTy4rzT8XREKwZoTfLqTZIBie777+/yd
OHXwFaM35dANS/gcOd7W0BUTC5XRZYaoWOREupr98SSE0QR1hKEDmfa5eGE4PkU3XfWT0cUbCISE
ZihUFu3HWCWeRfMv1k6gtxsMHsglM32tsYGlAOEs7/N30c2zfm28xQHqEzaf599FlkQgeqLtFFqz
r6bSSFw5hCpdJzvr+Hg2jd66prhfTSqwlY7XRJtWfiKaYUPGSVdtC3IqXMe9n8T5ZmVE9FqHvZh8
E8XkbDLJ4kmhMbgsifbE9nsXUYGVpf+2dOHCef63iheitE4RHQS0qEhL7pMXUx03OabAKHnV/VAn
aSLB5Rc91JQtBjALUqTdRBfICDayJI0CabZn6ezhPr3vird/1txe6mB59Pbaojc6QF2qIKhTWtpi
EDJfObrLmglD9pfR5mqUD6XStv/HyiXJGQvviKau8ySPHUqceiqyOlr6qjBDM9IORqLit3wQ9/5m
rpApkeikkMk6K8dQ/QA+k6Uq4hzATIwXBZjqL0aUHWNdJNn/y7yPWWywYFW9Sy/gIjvnVKuCIrWn
kwPScLjg4G7HLlGD4nX6sdm20eVn4XI5iF2LxuS+nRZFQoSAHoXrAaZvode4VuJ/UWtkW9EmnBhJ
6hkrS5rIdJ0jlDlc10+/ylNccjcWcooJnELytz9umpN5n+C+u4LPQrJH4DYNxTE3Ha4o0bHaxS2p
GbLtQ+hBZ7iAnYF3jAoo74k2nzo7LAmCfAR1d/rdJGub5gE0W3md0a7EtUyWcKtKBsyQW7sLhwpY
8sCfPzJyUk7PXUBYFzxNO1sWIdheVLHiCgtDRJ5TpmOaxePMGeTQ6UJD3BZcQ2930cvoJPiYqsFT
0wA0kvu809bWX+tcHKjsq2/xxVZjzFxufk5s16j+R3FhoLcJjq7sJvKe/nd8n7Hi6W7+3H/cP3Hr
3vPMdCWBeCo3UMVTS0dp1B9ibONNc/lLZg/SyUrITbMsMqH48Pei9eNhdwbA8lUwru0tusBZu5LB
xIttNSAv7x1Ir+Hx+uY+QIplYtEUJOMcv5OgKTy06zX3UxeH6O1ugGhqSTvVPfN0M18y8iDxeDv5
6Pt1tDypVjCbEBAFPyNV9mZCA2urIQxl8xjGH4W3k2VKsM9q3IMC1gMSM4lcxA+JrsRlyNPFzrNy
tk/ap8PLjuWElbPk9siO5caHJ9hpIYIuCtQ87/h/J9N/PJKV43BEjXFXY74JD67vO6Kw2+99upu2
oepjw6xgxhy/uLVjJtokKWpG/F5VDXNIfhXpyp4WHy80NWcTtex9FgI117GL2hTuLwqP/PY0xmTX
4RKrG30MgWkepzlPp7olEZsdgYdS3smUgMS3JoxEmIJEo3zzqB8M17EVo179ehOL5+JfXp4Y/+ci
LJn4jKakTY7i2KBYZF1bX5Qp3v2YrTZTtb8LPaTB7leCAvODrMZTeeBqJV0UD9PFWfEI+gpqh34Y
31wL2Hlb9QqwpXSuhK1enRY7kEjgSNugRmzJ9URl/5dmUELs0anfT/V0egMxDP3Gchv278j1uYbx
YZMl62SdXfIJusfgvWGI+/9CqSp3wt9xgZOU1AGp9O/Ux457/Vlug/Et389crr6dRq2JMJvis3d/
OnME0PdnwdDrX9S6BQUGQHmyGPcaXfgyMQaO4eSCYYNSXGOAjlN8mzy2BJAo6GNplxB8Ov/UXRf7
Ueleg0d2If2qjaYt50VOuTLgr2+YAGsi7O5jKpphXmDyV9WKGLwdDveFBUZKMXSf82shaBiGdGuy
/nCto8pzE3SQf6g87V/AowY0iRf3rRLuNqpdpDYJIOlloPtKeyPPSMcX4qWFt5UQ6vr5756ZqMEs
qylY3GhX8hobh+j/NLJxKLH8GdZuI8QgWuOirPkBzUqbbSu7dJqqy6jv700eJqe2HjUC6I3AQn60
41kqDFW8IKe374gQuZX4d2tetZZD0ys0AHr85asBTTuyaG36d3f/ASOC5NrNKHuLlGJeOCe33h5j
VYnmGv61R+SpiaE4yk0yOc3uMQG30+meadDxdPb68CSgEgdsyQWzhW1XyGTgOG67d3rwRaRodSMb
HY4p6eqqsk2eK0RMELIgIz21zCVe0UgaZNg18zhdSd+mSy7V1Bdgb4dnVGbpwCQ4w3zXQ1aKXABz
ScCTbjwyGX7impcNcodnXCcMfiU2K3bQaO5d3Yku12D4F4hpEg25OKt1xt+z8GgB3b0mLecA0G2r
DYv9cRVXED/iLCYqfL6Aru1c5w2gkFFtvH9Z7tPw1e9zA6JwqAxT9fxjSuyF+s3MuOSy6/ggENuz
wQ73r/nQqkhlxK2yfLpC5n5n+vHVVdhoZeBIn/blN84WQXBRefoVVIb+wwUjB5uDM2goRllAafA6
tYiEvMPC95VJOnPKcFs4yLg/eFtj4ZW4L5WdraCU5nraJ8/KYRqBywEEK0l6MZ8VlI/t4BIcOQsk
V3R8Q32hoTGAjida1KsebHnm9EnYentVva2MpQ8O72lNlHKFMSaoAf/xIcdyUDKVpwGgF3kF5tle
g1/nbfbaEeLgcZrDF6k95Y1cyZtvIy9700nyTNuqx/EyD1Jk1589zhAX92HLZzVVbQ/SF3joJt4z
YLbojumrCN+bADMCIIVt53Y6rFCQlntxUcAAwi+zbpsHh/D36W3Nd8PYy6AvTVq+fv5F2pp+yz+G
KKTrB5wXXdqF0bRQpr/xIFABVf8kMbiAdFREkDMLJuFLyQMzDNxrfJ5h8ZkxHGf+bTzsBLygpWds
+NW5e2muBfn7MQ2h5j3cop9xjjotIQfy/nOZAPmQjBo7MMMPpdDhBJYA2ZbxA9MrfGmN/5JgfE58
wEF4eg84ShRX1fhDEIqrFKuHb1ZNYxY145ns8+GAJAER75nnPfx2vtruI45txO5Lvn9RKRl1JEG7
5R877z+j+LS0QsYFG8MXRJBQOQxONt4o+PcNKYXJ6IVg3lBeDbGctctQkjF/w6ulI3h7zpt9JPei
1/23u/LUFEdvjPn8m561Xq5XjIDHQVFrPhz+TgPfR3N+F0gA7gmQzcGMUzM4bqJy2DucqtAwydky
DANLZtgWQ/fa01Ej6OTCvOvHUqN725noIOjRKRD1OeYS5o8ET55OTeN/XBWFbC8H3mO95qyltoVI
bukeFzoPNBnTd2/6jnJL2B1M7GfT3rDiouvSfYT4QWYW+aRIPXv9zTIN1AMzF9JOLkww2GM0Y37P
rOt6iMsB2Xl9qIMF+MjZTLsQZ7yz+f57GSyyDjnz+WkHw+6G7EYD/H/yIE6knCmoGV9cp8e1T+fh
x/cBCUM1IG+8EpfyFrdvZBL1QSlEM+ABL6OH1lmy+gHZEDZl6j0SSXDyZidp8SQ5GzlSYzjEE9S9
SGhvz6ZvBYw/qcHevFLtlKAXrri+8eKLwjRk5Eq2Kb5vBEus5g7Z/UNgjxluhumRsVQgwxS0n1jp
OBoXKQE5mSK42oX8ViISg4DuPtjpF+UrdirdVZ24Dfjk9O/7X+6Hjj//AitdDpPQeIL4l1jXUeyO
/LkLGRbgahK+jncZWw+z/tW1J01Z/PMzckNpZwSFcgvk3YUYLdv4VPtVGSdkWW//XFRTtUX4pTcR
FgSAZUgRwKzrBPpxjQZHF/1k6hmkluClCCTXOcgpxJNv6R2+wshIVboKqm80xyB5S14V8ALYvwbI
3rozVU29IPPD0ObhILOB2c8kogo4z2B2GR3mTnBv83GLHeSBusN8ZwxORSDvG5G9YeXdiButSVET
32EME1dnF77o0KoZ+mU6Ya5eBHbqpYlyysN2mVNJ/Hv570clca6xfeUHwVzVFxSbqxEjp3aDHB/f
oaoTW2NC1aN/d8rlnILBfZxDjZFlNjMF4oyFM2q0koMvi3+xI53oEHwrh1fYni0w1OiZMca9EPl3
BZlNndcFAWaSlYR/e9Z6xUjraASJvtxHjhikWBHuaJcT71JlwWrSUbUpC8lFCEQ6TXG2S7TcFR5j
rK6ZCgIIAKRR+S1pDyaLQFFkThnovN6S/rBsciohNQt2r0ZgaW46s1oGxA14/9gYlEYvafCbTVFb
aUcfI8lHVF/1cy7L/LkrLX3Jgvn4Wme73iVmXdQ250cjZtCjIf6lHIaL89blbE0+nA1GE5ykAJTv
GsFyzfJ+EPN8Hqgmk09WBNb3XKyRJqkkNcMWqLW3H6TiSgIpywZVnqpOPc7aa0s8wJqCxePnv6i0
LlF1gOzEez9dGqnP9IeJlfHK+JZ9C+JQli5EqVWOMZf7hSn0vPpnaMQ00jBP/hCeok0VzQPeqZya
IxHAr4ymlCktDFDyAhb9omAlAuMbzu3CR7puqngAGxY0BN07Z28WRgIhl7t5457mD0GXxkAeDNER
r8jLHDPXborUQuaxfxscBIII3dKbX3D8R04OCDGnCDWk8+g/uXAzuWk3AfZRJguWCGOWT3ofT93T
JOdAjctvcKElHl3CO/twj0ZqsGeUKrP8LQNr72Iw9PkgDUX1TwdylCurVoNjBabhet+uvSrby0Tw
2Al3ENvHYPWAEecjmlqev5RLrO6Sba8jhBc0ADcefnOSBaYAXFn80jLCwn7ZiXFrssLN1ejSlEAU
/VtMY9P4j6LXZ9H3w1Y6cTmgdBjsHoHlxeTjTDpc0nXITE9rsOtvA9QzpS8eQYeHG7SW08Zmh6/Q
MJPh6FK64ChhNi0ZPiXCkE+N0Yn1SubQzznCkQ1plIUvMeJ+axxCajXxBqO9N8WdtlCziyzGNMov
UGbC2Wot/nuZxhWkUjK+4vTWCwR2jfgae6pUV4rIszHTUhUiGxnvkF8PZfwQZGEF0zXh8vEZWwE4
MOyKvEXR9rJvDOelSdQPXUL90tlTeGq+jxop+/lsLZrXh8mGMuUjXddjVMv6y7nFYKGLj5NtMIrb
zOcn877HP43KV3ZtXpTFwMKG8PQaY/qkaGfWQhvH34vDt171qNAwtm87kLXVDmb1xQp5D7sUokL8
JR4nsYZ2oV0AF1e3K4wwDxokQHAHfsW7Jfschlmf9ASm3es+0x0/QPedAcjYJrgKa4LH9qxvjZwt
XOSSvxGIF9VNsZyPRdBckNURDBhvkDWXQ27ZckXjg8V9K05wG1o7du50HbGUUL7qE4O7C+7b9RUO
6kKueUUdyw13Qrv9MCjq6+G8paOa3zLvZzzUcis7JxST2sVWci+KNmfrDFdZw9Hbl27CIHDFZCxO
xLuYHX6mQvd/2Wic2IMHXro+zPncNAmewJKXWXbI0PgGrecFDZeD6IA4OrfBRNGif87Jq7R1gLMr
Luu4LFAoOsBADjy1lQeDiL+zVPgYzVOrHDy5dEWVDUJmXQ3XBuOBWjMv8QoB4Lq6qofkRday9ztf
j4l9GAnBEk9B+sgrLEnfCCq30XuCkw5NR33wXxcs9uOCs4gWuh7DPSgGSi0/8dht6sE0vsmca9uT
/IRNh/khLVM+oiNWNNExofk8/rAapDY9m5IRi1iKJSpAF7dqzUgOrMr/W+2PKKV8K2AyQpOwKytf
Vm1xmacvNs5Nw+kYMiutskVP0DhMr4eSw3feiMyID5QqqzzXcUhb2h+1EyBlrZ84/+kI6RtqlEZl
MYyFB2ME5Ree9nX1vJxF8tzhsSdsnG7kU7xPIooV2WqaVeFOHSwjTl6wf6rw66Kje+6a2nlol4S8
jl5X+SOIhbNb+NwzePcHsUbEKQtWJEHxA2JEydHGzFTz5opWfPfCuAqmMGs+YW5J32+tyeP1rk+j
hRbie/ABLOjWRmzYKGA7y1D4DRCoaMZOu8j08he8a/pJltyYJ9FB5Aryi89OM+ugbnk6USxIJCxV
rujiot0XPjnXlkK59mafgHFh3gBSAyMHcblfs21N0ngWhkWf0IInF3EnaQpqzDMg/IqaIH71EfHF
/uhU4Xbws1BBmw0vMeam4OtVTN1/gu4jronsaiLBjetWrnvHbbWKNg/uoQOYMOWnMNUdOLy6fU/7
vlVwqoQpypp96+bCsPsu9c8W2yrF78/a8b/MmPw9SbrdJMESKvN5Nb4kpa7PgY0Ortu2jExq/BDh
M+ZGv9q6w7b+e7cnG1b5/uaIcUg8jr8ltwu49fttm8uBxYf/cHtXXs9SKhz6w3SE9KeH0yLSarKK
x+8hTkMXTuhIlamrLcridVa8dR4WcNuYUH88m7v4sJ1S/crAluocQB+NCEm4ItuokD9Jrs6Mieoi
U5SsZ3gXzChVULM1zxjTkJ8ZN2VOIEVRdElIIb9LKzyFTDzx0L2rE6OU9bkPZqE2MZmhmZ3xjW7T
uU44KSHEpP9+HrsApTmsWvcFGZXiIUcHDVW/9RP6NlMRPijO0LllT4W4Pp3MYI4r7pLYlsRYiEi/
fw4M0uPIcKEcs+3hsZvQf61FequnsW5GMl49z0klbUlzOqjGAN3l9PDc2ONBCWs+s6ZQaM/5H8io
BmME6736ACBVzJ0Ykf84ViD8sXJeLIAFz7s4xBDdJVtHEgDv6eq1N46kMrE1FfvUmgOfzSPpWRUc
vFj+AQsBBUULCxrWwuTz7GOfC6Nsgi9JzqAeQwNYpyGWVY33K2juAcVLRh7TD70GeBVv+Gpx4nyY
1peQ/7orzreWp+f5N3aAxkzyeM9BVhIdV//nR340jsqYhA2kLySqgtzAa9HwrV8x3WJ215ZVttbE
nC8Rm0fZKUZ+dYv8zSql7AFeQo1jlzFpV08L3P2d8iFgVcFoVTHk6UtBPi9wq3s8+cRUhYoXc5jn
2nubCud3K/8aGJUDcK3j+of9yfkaF/f4Wlsb0X+NF4CpZwaoTYhTHhmMtQAwx5X2ncr5+cPNUFtR
q1FzxXlLDk2NvBx9cC1xIYwL8AVHBllNbNM64Mdx1Y2phOnm0vFRdchXsWhebkwJApWrnvBWGbAV
lee+PX2/gMLXyj9HHUmbcQ0PNE+AwRGa/WDaWV9cJSJu8OhiGydtDoZARHKfXvFwfP24wPjmaXhk
5izAAbpJ7wo7VkuBHnXS7CQT2GaWLT/kZRZPVrQ0YHRxjsviGzlLWm3Ivuky2Kw7XBykyO13vlu4
6qS8gj/VXqaZtJhnp9oQA38Z2I080OBGygpwGA7hmhDdIPu116oJ+rXrWi71iELzyLWyCEii5t2y
Hbx5mAwYe2WFryO0Gm2WU+ofD+lvBtzlSNhj96ErKbV7u/dQfDxyThNDDNM12mrJsj7OVyNwXZSU
jEsDONSXd7OpEbvxduodSEsmOhfBu7L1r4pO6EPjxQVNIhb5tUud1VIHomBuv0pWl+5QF4ODIgsp
vKR+iloeggJQpAK+BTmt3xue8RLT70FP0Yd5ygaLaPDWpP+VjUkWZOMDff0MYn4dhU4La7UFuB6B
xSdTQqlcQPhCTr4Bfj4lH+LYjgPbcUQxDlIzxrAvjmI7Rtgg2wDpoLmx6pUAdDV56d2lWlG+LfCm
3yd+mBNfNXWaTgpDesStpHBM57J0K7IHruqAwmwIEDPyn3I6IcCgnbE2UTIBQP3J0G0qr856Vb0J
EAPmO+sOUSAEjycgOVNPVaAB88yU3KwNM2pjNrTweUfqvpZd6oQD5jTmMEyOM/QxPJXRODMtu76V
/StPveecA9OBGWTweE/70s4qCz8vtj9X7I4jGmtpIJvb+pqtv8IfpGrbHf27zPnJK1qo1dH0YszX
3e+3nImdMmOCTRmxXm1jjYthj13rBJ2Iwp4abka05v/IQpPI4S6zdKHQgXb1wvHuCaI/uGc0uXxy
LrrE6HOCUSkpGoYuXyRmx6veG6sSJaICgJPY5Yi1v4cICxxWzxRDBiJsz5ODdp7XBORky0QIrfK8
gYGLkCQ6GPaYoKkbMZ/gmfb2gvLLGvYQhJ/J4nv5abHnC5rqXwo+o1nNRKEc0sGOIqwfdnu7808U
+27M13FS3t2If/XVr4Pq6HdcFjDsdfbR1l1s6iyrBsgCiPiIgzctVR/0dBGNh4JUCzyACE5teq/U
sPwNwITvPgc8ZfdP6Jpx4NIGZFQW1PL6hfbC5Nj0+LcF5Fs7vtzzPVaO8DjvdFPzin0jquH5Vfaq
VcasX8H6rzzGg9w/2w/sV+4gsOJYLc8X7AsCl5/1DeeonXz3bWIlsfLMx/YrZRweufHkSGkKaL3R
JhqNd2A+HqKIeMw0nThM26rQfric15me+utE+umdi/7Fy4jzxgripuihvTMVxGp/N8bDtNesOHpo
9PD+YsCxscvZdpKFm9tWJnyd8Sg/juRoCQgq1aY1g/k2pxE9dcOKz8WcptTV2FGj2z/GxBQ+AK0U
8CJ7820IbA0rhUiCjq0ZZwijJFDyF/tmSY5dB0HF8oxszRMyJ/aBGlyhbaZEyEB46rG14TQjoYyU
196rNAsx4twOrLTxMwp3RUWKEgM8dyzBQyqPnwIYSxydPvSAkUSv6gn4sRn+Nyzw8puiF06MFzCz
y76j773rPSYZ01Wv1JXdWsm07R8eesIPlOTMBdNJslf7NVr8DT0OFHsLvsNfpbfzQmxIfWJ0nOLX
eKQkEgekt4KNr/f7O/B5UZrULeERpR69mV8lDDrgbnCUaYnWlx3m5fvJScIFcKIQbKCqF0aMTfYj
+5eo/v/+ZlCKez3R0AP3AIERXHW0DUQJKc3orka5czBguzwoMUrYDbapA85bnZaMQHYS0aOzYAyQ
mrtNVIGtPW1KDK6/TNcZb/Lpro1rS0AsqUjH72cmZrdY04eixSxAPakPoGGBZ57x/0ZZDKGuUNA7
4aGXNpx6ZswPI4oK9JFtF1avlTasGJsKjJSvYSCJPKGQHFEdnL+63iH9dMPHdyXy2+6ZcgkxbBNH
JccBJUpLG7B4Osw7XztSV9qbJPaXQ6MYW1DfgmPYYZLSqE7h4O3nJSD52XjKlmgJXsUSY6tLsfeU
lDS9pC2+z03lSnxryOrfxM1g+A2Y2FF3xdEtoCBK/4Lq9QMRA2a73Ayejbpfc14UrwWOB6Y/eLux
mCIFTMkfWp7+rzOnwSTMTeLwELEZPQE6+YbQRs0eMllc8o6lcvdTAJwewvWHiMEDPxya394XD98u
IwxzHINJEsAuAtzljl8tQdAVYbi1ITL/CAZaOQ1Y5u2dKWSL7TMqlWvQFBT2QJxMwl5DmzOcaHfl
Uc0usodXmUzoFKIkDgWZ+tMWC0BAGGWcrj55LAYA4ccEU0L/sa4N8UjCBBQ7WNgfoC6kZy+WM65e
bRQXlvEJ28twQW3z0eCkJ8hH3PYmUMpbPLZvRE9yRCouaGvQXyZilvVR2pckVGPRuogdJYqerxN0
GEf+SsAUhUe0aZwUTnehevpLcnAThPQuk/AxcHz54JWB4PC6d6nPG9hh1ywGARhN1KLwVym1XBEL
nXE/wQ2027a0jlgMb3xtCdgmnCdUU7cNpPmi9zwU+QR23Qly+9Y+B6QnRZIF+uGtjUzERHKnjBjL
wAPhS8x5/y2abz/ltpfjrxgMfOU/rJS2L8937vOpdOUWQnNeBz58HjqkJIbRqJg10DdZwNLAGYU9
1d7RWB2ucEzYQx643yEjbDTGoxqh3wyWquBpNMQqtTSzk13zYnadlKGuuy0pTzuQb0RWnphsBDcy
LRg8yeUgUKBaUc8DeHA0LNvNr6Nf2WaO7Q3yICoCynXw62viSKm2e75M9f4G2m1fwbLvZXvE8JRL
rnruLo4eXUHwCSHrGrTTDrigXoT84BbzhdB5z+wgf6tE8q3UTjLYWt81pTKXbuOdaHhHEvFX6tNa
KRIDOS7thQzG/ne3e1qnp3+oZJqiCbJRyaQt/8hICvhuIQNKPby3C+MLvrdc2jF0C/9YzyaohNGK
NTDs8p2tjKIa4KttQKZsEIXcms9N+F0tGwimpo7zS0Zbn0BkgZixPBdRakrD1l74I1QDrPc+SfD3
eoptWgAn72F0qoFsDu5o+LIDaB+Rm4YYvog39IdAHmQfOOkGNxxWGkhBvPLpNvy1IlCuDy9afxsT
9EUdjM4fpLsnCJpPBcLtXi9DLh/wgWyn8CYpixnTyxb6BxKd8yltN1UDkQJL8n5VUqITT7tPcwSj
fRWMY4D3/vXZsex7rHERTzDsyhdeHgdpb42CbIA7XcmO4bKDqS8yoSoBY7DWQSDdXqL2fIGNtx/e
TMNeQhz8rLRkXPfza0XJHnN71wDjcx9bNQTh8M3RiWflVk7dLc36lJ2bD/om5fdKvA8dxOLhvZVh
yzD0NQwkuIU1r6STATuSk/QKU6lGBC2dr1heqBpB5tByEnFMTif06nkxo6zWnPSxrh2xg52pI6qL
ICQYOLiM7KiE9pN1ta4UHF1+bDN/IbgB0bnVIUvgbkZrViXDvSaPoMDO/u7D/kX+BpCKepDYSDRJ
ubovoEWj+lTWxkkgH5zDHqKcEsRp1K4DOt0PwCxM91oLhyKIUMtpLvNtFcox4AvnqVQtYoMju5ol
KytcoXEcL8gi0YRxzplytaLQon2BAZCvrMQ10RqaWx8PbljD9MI5BT2bUGf+5RV6nnOKH+JxGWUh
YP6Ljy4fQVRr+WyfClBUnNG01LxXpWSJuJHRtU+UFk135/CvmC2sfmla02uD7fuIvtjXDPXgJlLx
cW7kzQ2E7K9+EJvEMkb58gnAihVyn7zGkTIhKLgKFPRRJP2HONqtf62IARbNi9i2G1uPCFIyTX/d
Qiff9FU3qpwynHfu077ow0jteD/i0NE9qpflt5GoUcVNHL8hhxVWrJeVKZNEv55BrpcgtUgs/9qf
LyuWlUacUIvpVWy8JyGldPe5BdHyRfHI1asTLLsy7Zw/9p2+9+EImpHOglrD7tWMFDpwNzgwRbON
w8f0BrxlfY9C8TwcQpk47tf7HS5beyeaIMq2dJeEaePMwrupHrjMpM/qZSJqAynP07Ise3TulftT
cDeccSLB84z9m7B05mIiv6+6d8BDu+Cg6fbZdjTrCxBuhumeO+w99rcqDilHxr3z6jAtNgFxaE8P
gec58g4PjBNoLOetAHR8FgWkAcVU28at4gc5pJdHGnOPy2MU/omZ98qFU4xRX8WB9tA3VQSeJNZz
5S/KjpneoKjlf3sn/RTgWJwof8cxqGrbTP9GHNPkBns7f+KlIWlS1PsawfN/8Tdx3gnID04UEZ7l
YSX0gZS+BMbDAieUu0D6Wh6Ff8bbsPObsTcTuI6OmMWFxjeSZ3pfi/OBSd93ymo8NwsDR8ngVmQ1
BXZj48z9KgCtTmVDIQyaYOpfODegV+TzHPJQD2C8yPW9eV4JAQ+wd29v695RXI6OnR9F6XU58Gd6
jRWoe74VXnah0ixNkw4sP3Iik0jWFqZaoW+IUCaOAPScVhSeCxzusK2SO+w+dkx9OdUOGLlIdK4r
z4wt3fx88by2iGdXj5PIdB8wc5EzmBOqPwhYjBOQ9ijWwWBVewFXhI4kiyHqQIiw9FPrAyvPRV0L
7ydkd3o1HIviDDX/rfZEpyKhUw5A8YmP9SVtyFbV6JfZpWUlw188tCb/k9JKuYgPyY5ma4CQp6Kw
fZ9AxXPnzehdWZgqfdHrKToqlBOzBWrwkR2t1ryrkKLWDZxzWMB9O4KxLj5cLgVDzXN2kXXoI/tz
N2SR3n5xH0iPXhFA610juVob2tlCtwtL8LlJC8c+ZSmjnCJKlHItXqxeZY7ukkUCX+GSAwYPpy7a
6zdmSGOrVef60ltR3OQC9rbOyZw4++Np4qCtzHaTRfXCO7IqC7y5bwJ0BSLLhdNrOwiwGR0nsLNM
bG595K0jDt7A+GoYJHfSfYjwr/1OzUA0WrIZfFRZrTuM4yXIEzWSp2wlgI2vlTR75o7CyXi8GGGs
V1KZV9eI3LRAjdKi6sRZ33PFGFPuxj0fCpw/DDSvUyMMmHsoE/feRxfPIAoraySO4fK5K3QBdMC3
VWHSXwSj4goiY7GW9T6s3Yo6ccbnsjPWVlBEKQTchAPpoKA/OAwiEdQG/Rpc/U3qilPgsuK72R1h
GrJ7/2hC+I9aqsIfJTsq5kTmOnSfu32qd4ricN1xWuxkE/leTYJ38IBMgmM2b++K16iNpshSkNrq
37ad4BuptwvbpDLLULsDWjl8pgkhq+a89+rgCgaM4fKH+Ug0s0/dtNsGCV2f4kLZ2+eV23jTno/g
rP8umnglzNRakBOaHiA8FmM2Slbujp8iusEA5WeMmkvLG7Lhd/VPfEFMorxoSDnSdz2XgQEOcX3a
EEGMj5pNUCDdGmHr/AOraZeJhheE3RaqWM1U9NKYvvKzTQutD8MI8uAxuglwDsM1F3h7X7O1MEY3
eI/GxlzCc9TpT5pJmYbS4YA7Qfj5ZhfAtjn3PWWZeHyczg8OCvQaRva14DiPxTNSPkps8wMMxVxe
md0tu5916h62EcJZxlP0ils87hxFWoqpoSs64TIwHuOsvvSYy834usDbUhVIuznbsQrNEJ+Geegc
e/oRQ/TKkjerh6ushiJRct1KWz0YOn4XZIQVth8XGJCat/pxhJT3VK11V8g9Wl1eNPsTZ/Fm5o7O
nKUcUZmjMAXdSXHEYiRHKNR5i4Rg6vmL9En3uFhfDpq2kxXtHmB6ESFg+hbWSLNDmhukyvqSvn2H
M2fVaEtZAZrFNaPY6lYMCf42iuQynSZOPGzeTWYerZOl/nqT31DZTBAZU5MxCnnN112r8vO4k3mU
VowP5MLoPSFgMAj550Mhu+xqbi2Axyh6rAyDNqPjccFCpCEWHxqLKWJHHT0CeEjO3Txfi3/sy94p
fpW2U0/TCQRom7jGs8RjjRL1Nhm1yVdYnKSm5uQNXgy7OqHcZh2huKJW/il7oO4Y54xIzbkm92m0
qe1vd8eKl9YT0E82ryBoebXRTiyeSpCj/PAy0DIdFK7AbclUVLzZlRbcykdiuO24+fzADHcBF4MX
UG/5YJXYc/1H3rGvsWAPO9Kkc65TretqkoYgHghJ1/H81nnHkrxI7bBXgXNfqAG22S43jzItJH49
n3L8fRwaRCBzmYTLY4MzgWaPHFrgj1gPCQBsUzHBUdlSu1dfRTDjpfZq5LRP9on52mmzfK4n3SLj
mXcjCHf03oDCVAR2rVLqliNSmN1i8CZwEZBF7v086T3kZYbM7Mz3vdrMFByAXTHfvLzpkHesyJiS
8AzEib2zQsYVpxnM7EsU72GzQCtu5F2+wuKGre3H5Zm9d0DObZ3qg6/25A0zT7nhOmGxanmOnepA
khM8QV19oMoHiEXHz2Sev6EgJi0igln7ljpkJmdSt54waeSWf0hiJWx3ZmoMyTY5zfwyS7qvGf//
7qJVB34xXMLWMJFkOu2eqDAw1V0xOzrZMlyUFOKkZCJjU6HI801eAIGuFmev385Mjfm75WJNMEeZ
B2Ews+R2Eh2WWQ7BdBp4l/O3rZAkiqLnxWc/LyW09TELTtMVtOJSdBswYtXrd8Q9J6tIFcW38nH7
igMnurFtWbf1U4taKaBmfXRes5KX0KEZd6DEYQea393rXrIUen36zzblJAS5ZUAJKDlmdPw+ef6c
D7TgTihRoURjSsoDfJ2Q5lGahF02iMEo1qWLzesQG7HRXkZtI7lAznxT1ygPNy0IIsGJZFW3fgmc
Z8WXwDjJfYLCkktyPF4Ok36pMPfIuL1zhoHLDrmOjjcbvEUXXKwRwjarCx0Tb3kpodXHLmfTeDKU
+CE0IEoccJ3kUuPnsPWdo/SN4sG33v4D7sPNbWTKQAFD8xfZY/gmUIYNoTkTyvgYOhz4/8oREcXL
mN+xhjsZPR3PzHphKeHW1XbV/Yr85vGf7BX3eH+bQcSCotLZkcaxVGVkThxqlmgEKQ2qma6ckTGz
XwKEHQtE3p4s9xzY4kdGMjNGvaVWD4kw/O51qXeopMVbLKFjkUz/S+9vPr6e5S2jzpPcm6Xxfd3a
SqBsPcArar9m/7OBH8y8dk3eYSAcXsM44Doc+3ME+0CTZlqw4q3NlmkloF5+5cOosd5nIdLZ2HW5
yd5j2BICyDr3chT0xQtkpk+NjmOaWQ8dAekGCSFioqJuIc3Jxlk30b+9yPubZb8n65sefmKvFLgJ
lQatUotAdAeG/+zNOSqPrBvQtM/yhad+7zIskWkyOl0gTjZwQh3YWR/AMrvyh3Ea27TVPutXKOQt
S0QTtHIuzR+9mIpQ5NDxBK0YqKEjl8o24YFrCeQMVGGHsvjruHngrb02EDZnXJUWzNYcUxvppgUQ
carIJ06VznkSqtR9ZoQdq/viRLjJ/8HUjBqAgcbj+2zo8ftggjWvHuuxbqrdlvXug1IpdsBMjSqw
Zpw7NjPhy8FEdcsyf8lduDjs8HaZudyR7hDgkyjTHYYKquAdpDRZhwa/1OmvMoLUo4cB9fpBa8Px
UUSqCoT5uX2xU8bcEwzkl9yvxh1F4REG3K4qwzWTcj1mSTEs/XQHn+V9IXvQA1DMlZq+wZcXb5h6
WRxKP1Qa8cUtw6IZTUcsgCeWMA/2xqMBZ+kJ72S4HMoLcBpLVjFvkuskjv3RvmAqimoBynOtMYkH
JaygGPrl181Mia6Ag2MM27ypqNquKyMTagGQIC7dWztHMrcDifpdwebrWHwL+DL3LyG11XuFPWPo
a2OnEm3kUIc6Ccxdgyk2eYIp4ZvivMD9Tz+M7nUKfW20JWZYlCSX1p1NCeJubAnqVCBFolu23BPy
9ou89U/2otxyJRZgDsDOyWczJgLF6fT3mXl7g2uXaeOXEp3m3E/D+1cyKd9797oPu/AE+ZHYTXkC
5JQkuNtFePEbXLiz+804Vx8tHYGF8XpEozl6SE6m/x/E52jiYY6crMfF/8LBiJVWRNSbv9quO3XX
1peTtwn8QizON3vJd4EilAgx2yb3mtDitJ06BdrMqKXtsFHDxTp3+AB1B2OBgjOLvgZdMBoWM9av
s3fioDtogFAQh4LtVQQZIPb8z9aNdQN5BCB88XvYmMA87o1u1S/x3Y682USwZIQtlqRbGKKTLCRG
CdhVBRcBD44SDZg5zruajLn0FclnUSKy+sI+N9hBOZmxx7x6A/yZLz1ODhRqTbK9Ejz7ZEW0z5yg
pKVo/21XpUrQXsdEXXcaUkm1usAp5Su0mK+rsLpOYFnusbPHGqm3Ax2KyfQ+KOFFiRwf3SSU7TNX
lytZ3g1aPT0FVZwny9n7GBQXW6k1vcsmW4PLsXJ8TscK4q75D0eC8CJ33Y5N/4WpeyU+M+2SJrqh
EWVy1N5QJpjUO40cJod8aABTDRll5O6zrVmb4isLQUxcowNZdaiXPoeHErHu1bWDwE5mg8Dn/6yr
yXEYg7OgNJHSL3syErD0qS78gr/sZcKS7BjF3yrPI980PZjCTvoPqR+ggJi1ybCSR0wx0wyAdzMr
o58QWA5cpXYCouKY65SZLcGXjnpECYA88+pV6QGzRnW0rvohuIh1Cf9eenClAkUmkxLp6gZU1EeZ
iMCvifES/AYhjtsY4He+X0ZB5Yb9e2KlxzlTFsvTt9WuOcv6EFUqhUlDzz6uieF49/OIUVdZRXQ/
J56gpUE7HtJlpd7J5U249UcSA1Ci1YLnitT38DZF6PVekpkJIs31olAPiQyiUx8bv5YEVOR2O4lS
f49TkILWBrPTZnpHwkIEwlqcyqlt+slMQ+GegCmhObhwfsnagmM7ynygUXLpoRgMVJ9zBv7qZzX6
VIBfhZ7vzWf/DMQiB8TRHL9DwRKgosr69rhZJ7vvfD0sS18MqPU53NLt1sX9dKf+D425rvfWkUXq
JBsOIi4kEYXdNMhHc7I5Srdho//WWV+0cjvRpJGmEz6uyzfRrleYmLhX/K/RvE6EB+tm3s6WsNew
OtdqgOSl840mIbU3ATnQl8NFpIHAk2mqqHXr6W8UfzXCZuo5NGFpHLmzr1mZjwI4k+/IgTiPQ7hO
eJst5+GVgjtTec8A6nqshrBjQHU23BCcCyOCKGiqNCJwq79CfU4IcjVcUwPcnAl/e0xNzCbfk5R+
/OdD+iLZFE+GKl1QdJ+PUDGI8hmSjEt87tuB5BjClWoHxvSQFrVNwqx3x/NnkAkL+HKmtEWXoE0s
/V/fauPVxMr9wdT8r9YUhdDI9K/T1i49kAFZrb/Z9kn6TubH0XiFv1QxZMmvLU7Letyv5KGdtW9i
b+oGAjDFV8QWGCd4CBTN66KYoT/NZz7HR9GLbpybAL3EARe/GTUKm1Zzz7idiHQuSn3748ByTJSl
FzmNSpcg88vj2pBrsnbGvJyECiV/t4WkN3wzNSHIrxVDLt/T6FAUo9fQH7Y3JQU1JR0qhRv/qaY+
RRczC1XmuG57/GguRVAdKnCN4gGXOvuXlV3jZahSVOHPfVFqWVujWC2zGaeJT+t4SDOaHT7sXkOi
fRoc/xrjd2nmDZ0EtNGoyInOPKKhgfnXO2SiG8KWAGaOSfLa0Xpn86t/06I+INg2SqjB4DdMkokt
uZaHntk02EE623tg+1cADbw2lHnouC2pLBQM2RH1J+aTsIFC1Nq3xzBeSmatkBF2H0sFkmJ1MPy1
h2V4pdsjBT5m0FXoJUqqdYECyF5ktT02YAmRHvkLCrC8rB+19BcVXRUd2ppu5WI/93YxXHDTzSN3
vATh7AI+Qq7WYi7sSTqLM90+KbOblsT1Lftwm+WETekylU009wnNCMl/LO5xt2UWyZ+a4txJEQCh
Cvh6FGNl626AnA10JMI74Tw9QVbbaP1bIYY21vKXtiXwCvGFDSALyQXK3AWHgExMl/ZZH+h1Pt/o
YzmrgSmWYZ5Y9nfe4hHvrQzzEOfj18FQW3uQm0xznutUpTbBhTcWk1n49D4nBSVhM2Dk/103CH3B
A1fZOS5TRca80LUElnsm86pSC8CKdgZ40w/rbB7VF07sNfEEANLZXjV9CuQGZFKZ4jC4rBOR/p4i
lXzlDm5OVVdePSkLitGzyb0WPtZ8uhOl+lFLvMXOTa7OLMbCJzblwWRia/4a3HyaC+C7HEG5LG7y
9zHHDhhu39bTD3c9QbHqeBPr5yuYQkkxvlpj1Yp8+klUgvq3xpjHE2QgWDFCVAGrlPf/ahHtDcCt
xplBNUgFUZYr+bDl/GyoVetkq7yKDeiW0dED1fyyyKEZRej3VaemAUb1REDH3DAPrgix2BbuA+FM
yH0sqlGqj65E/elBp224VUeusoeMtkZC4XsSSn8GHcRRbw8nlGF8jrIFnxXDqYjlomrhHTA2Kng2
mlwAzIOD7RTtYMIvHgwpWNUIzNcrekqruSkcdmQHdOfOB5vWd2a0Ak4x4THzUC6qLPQDQH4AdO44
CnwANpSg+kqDDhDRD9Xws0TuoRHiAKwlbXga2OpjhQ9BpQFcDlPnkvpcHEGIf519YgSUnbFGRm+M
XtrJo0tnrpyE/hvIKFwkCdv4L5qkHKnVXkcZk1PM0Mbehfzqc3komemCyLiSmtdQGyTfmJv/2VLm
vQCH3JhZIw1j5gp9ztKk6FO/NQn7ZdwZXUqAbtAkh06u5fa7pt775APs8SKGXZORp5HrRGhxKkLN
Dk6dMZUmHbO9sFYCQI1zp5U2xTgNA7Ceufs/Qjuh/ey/lw/lhlC/lFzXV1sPLCSCKgGJUJsmFedC
kJFVUb8GbwrQxj7yvNziQjvhSt0IJwZ8vRpTh8r/N/L0LoqGU25OCEwBII9zgm7Ioo9QrqpvDsgE
hobO4Qd/nS6y2NUk6qPUbrP/J1G89srPbTPekgkYR4uSjHVQxBQLzdB2kqjFtwSApptxQ6cZhkqr
51s1YnvRCcjUDTP1ieSU2mF+tXCqI/L4h93ZTr3cZvGNqVi2usRKrkV7KvPoZGXyRt9r71mOqrp7
jo8bj2ZZOnz+FceO/W+0772CktlLXS3zgh1pUhEcvP+3OWxf2Mgcf3dd/AkAa5u4o16V7GiN0se1
8Vfn1gMViOmVFhQKRyH4vG3FgxWlhSNlnl9mW3OsY+xm1RDzYHJrvgFmQPcL6KKICAulhyHKhHZs
zacegUpOWl6y6DEpvHZ2zfr7iuWnzxAQm46i6DnLHWly9pJCCI//aerJrVMCb9KeFGESJ3YoboSc
gAbDjkq28EM23I+hurqxbs/ckBHiXi1PO/scnwor/z+JSmYXDk3gsbbEJA763Gh/D0l0fYgLwXuy
5pC8ZFxsnv83SKd7aa8Cq9zKWDF1oNKSUAp3LYEgjvFV9jVMe2pKIWvljv9Non39LpzPmYvc8YcM
vXCkA2M33+7fEt4LzbF2xUyhZpuNrwOI8L1AxFt7F1+FhO5wtzR3Qbo98AC2luCle/ncFMz0WiDB
syPamTuHtlXGodaieDY36wOTfyPNFF3xExlN77waM7aXQpGl6RNQ59Ntq8Qz9kyWl5mNsV2RmSjp
KhkJvBOyA0PLCUZbVJq2RwHZuDiZ+D3ZwVMkkZr4HxTMlQCOMk2S9k/MO/r/TES6XPXCK2Hv0fZI
1F7m11f2/wPw1ywKjARgddXcLX+T6WxHKkCa5kzh2KfmNo7EgYfYNu6yvCqYO3YBfnRy0tnPTHJG
lB2EF3R7jabv1enK/R1PEPtrhPQY6Bm7fx/zeKw9jbV9EnU23QQZIOVboL+k5igYjBGxLx7lbQHP
QnSa8CIOS7JTwiNno4jHsK2ZsfQnmLNj6Re2786RVz8kEg27tEz5eV2a2uJM+sOJiKaxP0KYk2kf
Rc6dv5q9pXmci1g8XCzV8JodlCKDIBDnsCj9DAAtWV2Rq6J9nwla9OVp9D05kjczGaJbig5SpDfg
z2In0Im1FaecYtEmWmdrfLkG3kOcmpvwpeIX0h0XK4D92JPPEy2DfyBQGymhDWewonMsc1iQ51Xp
XDPun4Le4/wJbR6WdzMadIazjst9GIn0YihneALRLWkjpEYHulXqB4xmF7KNtDh8aCBY0WjychRW
KuE+aK1MARWib3ui5JGqewIgokmDzA5NuaKCiNj2bFfGa5ZnkgD+S0scpYEl/Ss3vEivFpq7BFPH
JAxNHvKboiW/2wEaj2ONkzhoXuNkLwmg1IxCeIwb4UusYavQnl2Vkbo4NMcw1IywQ/EFnOwsq8t/
gA33TA4IRohedAyYH1NvKV5jX0jwXq1v5AJoDUTNDsffhXhosEgEP9kxMSze/pE5G8+CwX4FCkMt
OgolR1T0TRrAWSbhg0n5s9rdtOZXOIYbRMMceZp9nCq9WF/Fvgpmp7XyEFGvuedgrtP/+zoA3+0e
c3QtiHU+Pu6TFZeEXKu+0uVmepIvJlUi9DgdeuPxYM+WcLiVog5OZ/WNu9qlrorGy9HBtkZVcKQA
PekF0I6/MN6ECc1pLPvRZIkeyr5da1DkR1oGYIhQjxErXE1ODJ+iQR8zoCPh6L3mgJ9sqmGWM7cV
MR9z0StZfm5EunwFJI9xlwJAspGuLscJ6kB7zUpGbYxYcQzf+EmzwuX0cttu5puwgPzW8q5j6z0r
gPgq6BDc7w48AboyNLf7l7VnU2ZJkMG7Pi2gT8GrMu5Lj8d8ycIb9cxicJuqw73P+sHtOLUch2IY
5ZcvKOECSwrv+UAW1H1uT5VGMezv7hp5ljMdCXmDtWrQztYZn1BKHQAxk5TF0o3A1VN/NgRl6V9t
xW45y9FyMxAJI6owFxzkKMzogiYOH21bVrq6VaAhtGelgOPMu9nrm2QWI6fPXa7+p5S/5q7lpxbJ
OcZIeLF96XEhs1VjHpC/ZTY8Yef74d11u6vpVYlxssYcLSOfEL4GOnFTKhLaoWPuiWxcJ30zI0od
fRLEdo5nlYsRFuc5a2XgezpJt2rzH85ScnKnDaaUTyxgS0rycTSSVPHvk6JiNaWnQn955fnS1GP0
0BB43kwGt7KLWUDW4WLSShvwM+bohv3YxzM+218whM4m64OMQ6lIEI1cmDv1S7udSCC2/arMkoxD
z6UsTtSZHSlvhVujD1K9uB6GT2KTLVOZLrRxL7j2GnvzycA+kskBs8zuHOtyFhq0tiud62ZMvr5M
I93qQt3/t9HAMAEEDG8xSdr7AELlVa4zdL2if4R85TX1E78Lv9Zb6QJJHAmis/FHfv+d3hclhvrc
JzDWI84CdI0+9S9SzRwp2MTKGniFbHeEAMiNaj8Ap+twn321oQmd6r6048TntaCxYI+f+XJp+13G
GqcPJ54o58x3OuDA7q46y1ZPw9XzwchtkwWpHvjX8lDrnCKwivzb5THdBr1HnZHyHsJ5AjYAiJyo
wHC6wpHSFRVrmWmXBKMUBLWSbLYFbTMjm8+ZCkKexWZ9FAXgd7T0kfq5WA1e5l+UXvcxUbD+aqy5
bkDlLZ3f/6FmaFs3hmgL+FsXfFiFo8WgQUbMpqW/viYzwMtxgmHeLS0xfLh0l8xtKetcpAX89/fL
DmZIksP4Y+XJO9vl7ZHNivqeQWCD9FrYfMZIfmDHE4a/KtKEVvLUhK2UdIZBOmqLq/xFWT5ioCnX
LKOfFHhnn0o5Zgvu8D7I+fZ3m8obkwG3mnphNdQQHVl/BrOYYDDRIn+HJP6fypxUw4u6/GIKRoV7
Xx+FcDJP8NRzfAQCuNA6eJ/mXpiTiQuXSd8UGflAhhG2qJe1IhbGQyhB2D9UHINdM6Y8FVOtQbJW
tSd1uOaMbn3hQI1zTy5FvDGlxG1wrIZ87cVMNay1SzWUF8Gz2e1vDH055lJVHe40LY+eHXvMCpqD
E1UJ8pWT+Qe8oTwuS2iR1spdzlPYNuLO+7iAcxDP3Yz1RxETcb0GM7G58vEN+B1FOBiXQT4IAIqX
BHo0UzVpYfOgfMRFGGg3aP9+mU3orYJg0aokRYo89n4y74LVUHK/sqRs/NQp/mjHoQk29nrnuvrK
Xi4cfX/KJUXHfVltEwZ8DUbVfkel7Zfk8K9/Gp/DG+zZWKgNtCzkqkvu3//lcGLR9v47HkDbg1fd
q7UD/69YO13U9Qb6kChh6Kb7zRjwZNn8gYVduhlCO+qAO8Es9J80KZ3XsxWkQPpD+2mLPJaFvFAd
B7frgeteFXpjyflQaKxEDak2Og+1yEznUOZvTSrvox2T0VIPYFovqmmpCe5GwfqIjr0/6W417Nfn
cBEC2cZWVECYTj4KM62dGfQpqBd/f6pmP2UnAQo7lv8hW3BkcxomDWMMNMC25nYeKXXVEXxY+J4V
BfH8bKABoWiK3DVUXTMbHmJ5zZtL4aGjfU0g2WK0lj/JjnzqorJ5o480WXmwDtzCK4PcllqWa9rj
1T70DVDZ+T0pBfQSEDz8hrNdy/hGFttJgF5dq0dvZm35cIcb6OSXEfuqYUgkIopS+TARGTxSbhwS
RC7+uHwy7yEYSGXw+165FwxK2B3prEaUAgcQ9aeSu/2Ch01ahT7djrDaeYZ/l7yfwqKgA32dQja6
whbCmPgc19H/SxDAAMaq9zK45ktJqv1ikGneHzrjd2K0kGajOPUYc2lbbm6Ok+1NxJjh94wu0ZGb
bXyYEcsLI29+7wDguTa5Z/Y+IUV+FAENHqLcI1HVOpuqXMK+DXXsCyGaUbkMi45EjhyDLTM5prT+
ONeIUTv22uJEBz0dUQn3pwYRjO/CXDgwvMtL3/AFz+ArZwZGv2ecxQHI+44n2ghsEiAxR8X179pH
IksCdi4pYIkwsP/i0zJp9QlPEJBPp9aoOkdegDB/mPATuYIUnfnCTKlSGh8HPjJpVzuTnntg4mEc
COeQrAKZTlf0fjc4weK43dXXiI3KYr4CdHwLFLc7mde0i5MXOECA5ziIkkMh62qXQg1aONs6i0Dx
eV/DKFUmo6vKwPKmF3RDO+LtqN6TWjTaaZZNCGAdphAZBc6WB/ZZZt+yiRqFoe6Ifd1OqOmxDkti
hgOdswEqQA9u6eueA/alyJYDzi+YUfliJm6PRIRe9UdmN1MWYDc7vOml3/RmEu5i8sEL10PPZzpT
QcWCma3HxJZ34BjYT/uZHPwMDPO+Dw0pUJ/YVgGuWv0bgxPUm7sWd6dfXQljDx6LsaGe/MaoVNfC
sAKezp6+QyFCAB9TCLBjaUVZ9ShX3DBZ5PUUwVusMokv3ye2F4kIQZj/OZJI7kHTMYO72PISmf5W
noIvWwhyL74/uRyS+ibWDHNhg5Z7bYMvCN2ODB/zhyMjt5W+HUV+gYAZIn/cqhfZXUkEdvpBNlmW
Rj1TdJk7Ltfwy7KXWxfxoTZx4bYQcfC94uwK9yNOvnWi5s6huk7e+Wm68gJCx673vl2TS1M/otcJ
DcBjYONU9rgHRDQ+hjrP/bp4ZRCF/bx91xYqDez9ca/vClqtCnOTTefjAeXJ8HYPFzYCnkx3tvhV
fY5uRLS/xyabxy7r1dyd4cVIDSatDx7772GhKd0RSC9ebPHqPpBu0MDfPW4iaYdgVIuHoJrD6hZz
LNqXfNNDAr2pOqvjVEixW2q28fmDbJHjnuWF2v9u12aIZYsIwwkwzIhnAIcyRshD+iAhCpbr9+3e
lvrdezFRngSRVNOR4uYcEuaeSeVe33yXgSzjyi2QHUr5tJEgf8GLfEIrehn4ZOxKFG7qHU0OdDsf
4T4xihXHIp9OweFxCs6Boo6O69jFr1ukpKisGUPgt3oUVUHOWoCG0r0RbOHwj4Q+AswQnpt86UkF
m15pV/B02Z9q2ytNsSNdiTdiqw6PhyC2fl33hjMOsJszZ7oD2w9/o0o9W7SNAJvfS4UmLqMBsa56
cgTkXvlgeWHUKfrsHgUWYSN7A8UO+Oz876BeB6HxutT0orEgSfT6F93pGD1D1s4X9ZMGhwP7od/A
5fQSGUHAerlh372l9soY2D0BJYP7lhWSuqfXwwEpjcgJbdQUTGQ52BYx/CTey32VA9Cbi4cItVRv
8IUm92odbhtz5kuLMZ9epZcRS8PAeAz0NChk6qV2fL/ktu9aMQBff3EwlJdgFOph0cPGqJvZyAcd
ei3oPjbcF1Vlm4CiCFAjTK5CPxk5meh5S9YxJ52wXql5PFmrvx7bHgv8CuA3YbuJwZ0kkvWpP41C
2O0IGKTAWhppeV3HnhKoEwQB1Dt7XHLbYS4uAmkcppxrE6v2MTmHR3FxpNkHryGuyPKQHa/wlCEi
tmnP5X0A7uKIXNYv7r72eBXWKQUfpER91Zatuae+OTV9vPy/jW5GN2FI0eHhbzClkjg2wS0xAQcB
6YiKvdhV/VnZ+ssINjqAlmBAU+Xr6cFkGZG00Bg9A4bwc0piuk9aT1MmwmNg3/PJkuPfvk0REXOV
3Pl7ZNJA43CnuJxE8OTth7FrnqknL0vOKg0zCC0sKW89rflmdg1slobnEUKPYCLfP9KIa3WDpDA/
erLOsk44N16+9C54YMlVwZ051dlsgjwaBDoaVJZyBAaqTEKcFhKuN8CG+9LohRVuB5JLhUD/3Ss3
jH3Dh8eC3EbsDE/QM+c5fC1jFKyRhFgsIL1WbN3vtg6xj0Li9Yoqvrvti463WbAbZvAqGYxBwYaK
x1jHRXJ6TNXb+PYjSJhFOeaQ8hFIVOPTlbSzD+1upQBliHZSDGNuht++Do0Y6kd0EZxff+ccIk7W
89xfcNzZgr5vaCi32C3lnRPLbZbzofpXGT1nEGvAfSqy8vYQFg1cniGc8HVhih7YSeG5P5/TZOIk
xPEo2usgF6BSfzfpDzwu6TaPtAihn4HLFR41n987lpOdx2fsxsHVYWi4PusRai77u7qLyO4RzIGo
nvAi5hyUSPcAQv5juq8Gz/uLP/feTAKvb70R8oCSpbljbr4lEFrM1MedLQ3ek1mS8WaJXrxPCaRo
Ldh/NMdd8yN2zRhYpl3tC0L+bxn5C3F82ERPk32w2XLe+IrpcXlwN1WLybWd/NdXa2ZYcpRYFreU
UH3D9xB0xRGCrUDdT0MuOwkS/p8Nk9mwNDoHOJTMC3f/twkaNidJuYePf30XaqGniTnIOmnYfesX
12q2g+o3CXWlckuyvKIsK8J7GYBVCjYJ/0EbYvsQJWKqXHD/vaaDsZAAsmUl0mAaljtlHQKqUj8H
9lBsQusOkeGWldKJNcKVGaezpBMI4qyaxwMQElP0lwdLcWulOqDcXe3DEm3HnHS4L/h5Zc7LfRrB
/i6MZ9EfEAMziPbl+xfTf8CYVVxiyHuwp1bEipr71hUTyeaFVU5r4i5DHCPxWhRshqTzObu+xZCh
uJZw+AW7e4CWn8W+jkq/bLddu+YBBA1GHcLxr+UwbVOIpmmJnmmZhKvR/p1f5MKLO8AeXF6SMTtq
VZKigrU9G0wkqhwTBnIQm5ajyrFTYAHJ8SKrs3/NyEw/4i3eCOPerpCQjr5XnuN1o8LRATtvRXQ3
N9+U6r1p+qcxpD8jUFWOHQKxclkpKWOpBV1UTy20MQK/NOJK02Zdcu03CpfQk9Ameqd3TDpFeH9V
jG1e3YdFy9rXqE+eMTJIcGKVzJMjTEtWsuF+IrxbbgSn9Q/i7pT5POsF4yrwEYdmrnjhCuu9U5Tw
bvcBOsxx+fdRTjRuA2aPXU0gONcc704xYSrkIgwa+kfrP8ErF3btB0eLwBiBR78d/3aQvhLukxur
fzSAv4nUTethRgyTglmJz2DEA2yKa61tqKaqPk00br7iGp5r3vA+LBZCDdEsTZLtLKERQvVWFPHC
p1EsmPWU0LapO/GXkwPXJOjM2K13wLW5ukdgLzA4qr4UOEAOuMOMdkQOlF246Mb0jU6YDFnS0UAQ
esBGJabX2JG0WMj5aPFbpLDLbxmy/+lthCiOQTEr0vsl27u6vSX6f7dNxGdVC6hO5Yi/JtvieWig
jBVlSbYMfbAXuLpGsjbpH1Ds9qZ/GlWrplX23+pvaINBd5lJd5u/0Rgg2MrL0PSWdWV6fG+Ut2nE
ChRPpbMHT+oSoIA+DDDLEe0nMFIbtBniZl+JegFBphnHcNDHRlEbZzo0kQcwFOjS7Fnl+jC2Ntr6
kJptLakqJcoK0uE3JnuDAreUdbfeLmY7KxloZsZHfCIldSSkFRwnvwOT4pUNuwVm3kV4JGNGlBJe
45QiQEfq0yEh6txHJTB0nHJnPL9BUNGtSRnzgtAJdePf7vvfvhxX6vcQpPhmrf/P8x7D53+KkWFq
JR5zw3Az5YrrqF7trijaxXWG/u/bLgMk6HM+UYDb/3LIwJPRtO9m9zWTw6o4cPZXvynSAE+CC47y
vkr4Sr6BcGPn46cnq2P/9ACldWWYJT74p1gP0NNn1p0VsvfQK9Fak+6ISKwxwZA8zq1gp2WMWvWw
kQZmSLB6dejjLvUQ2Usz7jPQPWaZjGWzO6QTlhlCGTGPFTY3SlY7lyXk7Q7zYapMfGF9nkff2wXO
WhIcOjVTRykYCOa5oQrWZfO+hDpqTnSiFTKG5Y5V4YKkxYAFbztHqEc8vvORi0y04zETcDfeVZLC
aa4lSfxJJi33Mc7QWZBxrhDlPPTEV8SV01TyTReyOT/MYeXKMfr08sgfL0WYCySlq+WkCpI73zzj
yedeW34iR7fs3NAGKVkR/0VNAdjAIstv1g1cyx2bSC/tc4EgW3fEBdLzG2cf6TadAyX4hDX8QQ8L
bv2Af3Sjwvx5BnWEHn0JV28tBVG/0d2cTFJMGNHOmIZXJc6ipwaNgJHT7dr5NA7gxIoojFohXmt1
2+W/iLPyr0pWhsmHNAhZlt3MCi2i6oN0osDWMOyrCbmC7hVg6LkwrnKBVLzGGHXvsix5N8oeXMpE
FEOgLaawnn/3YGydvoLtvOzMN16ibCfW1JteeoMXr88B0qGgJC3KLHHobuTLEez0QBt0dYWC6dm6
pB0Os/QJTjcX7dVHvxUZt9CjWV8yomhXDwmXR3L/4dVkR0ElAlLeDG8sUEXh094t8PUB/L0GiJ3h
jloHcCI76TnmURXYl/1X+bf933KY/hj180k/MLrZty2VcB/XcxrPhXldKXKSYl7mEIuYW878njQz
a1KlAeqPlpuK+TJPUnmn9NJaaM+39UJCKYXW4BzSP240ojDzM2pvJU83AKxgwFp45p6u3WQqKSrx
NBObHmZLQpPOx2OSIEE8JLrRQpoVkk1GyYhd2ftDA5V2vEjN9NSDG94fLFwt/MTOcGLF+N+3xunY
mee3idORe00ENTCqVUxABD061TKR+Cr2TH/6rubF5Z/55wiMjk22UKjQHn4xcTovij14rd8JALiy
Ggi2nSVOVk44IeVRp2B8YgA6FjhZkuahbZ6LB6NvTAKXshlfMjwb0YwUWWUDc4mxQBjv+uQwQS21
52MploVByl0HYh2Cj0qztkfX3iZx+MRfXQbJP/1KNKGJ7FliG43ulY95xgdV/jSQpW0PJsIwN8lM
WV0jILzJgU/7fXLur2F/JbijLYfSaFpqCC9dW4T1MF9uTIiz1s8KdVGJDQ3imARaMK4vITG896q0
CyjNESyBTd3jKr61aRoTY/2/gYWZsxv3IMGr7JQ8oauTa5blyJ3UfOiX1Q+IF2kTCCy/6Z75EQ6C
Dp+5y7otYQCFeAb/1OIZTKhK/43q8M0bJJDqTyL5E2D6AqmEagmW19vccVPZgg91bErwoS/O9Jg2
7W5/N7mAtnEZHvEVz3PuyvEqFtMffXgsl+qb8nUraYXf3ByxJI4r/I2B+R+D/ddlqUtEAnENHzVe
G7r+13nIjQ4xzILY4sFWX8x0cyfkG4VNnKaiNL8kr47pOUnyl1Su/EQvmkCrbduWqugeBJxKLsXD
nSoeFqtIKpr3VfW1p1+u32vgMZVqdm0IlMJWSBbfwvpvFyHKojKBDaHoh5V0w6CvEG3UtCg6pkKp
yKfq83IO2lnxVzQFEbsYB/pRhZx41N9nbVZvh0AFKFFn3i3aAY8oZirVIbEMJc3TV4WNpyvncGRZ
klP3FPxbZF0v7ftPtdKh2rDjD22s/o+aaF+v7Pxeeoa+sQdzJaral7SZQVQEZz86H2TLVubW/5bh
PHghe0zGXZWIMskmipwoDy5A/zFnELwGkLnYasHwlWSnuKYWajh4ByEKYm8Q6TWYTINljdtE/v/j
W0C4KtuPp5bBRX0gBl657T43Ry02mecdB5BtLCBF16Im3MbGYMQqHUgPgcoAFePa+lqrNxBt9Sqc
lEX2zdZI+JbP+OUKz7wfmDFkgOhbYSb7klZpV3w+yEh9NxhzX81Y70QL3JwjjRrhrhHRJRWw9f1h
s50aqbgIbYyPyA/zpL1TT+m0h4l6JVBtK7MJ/VcLD6FnKsVu2SLgBImiLGjNz0PSjPP7XnqnOfvj
0v4dy77WuzjLDXlinLnA26ZlEu4TMXQPNw+tqcsC2Wsf4VvjsfAzL2oap3dZBf+5xxa+B/M1ehws
98TBbo0JyIPr4EUUSDwWiMqi0InUAdgmAosNDVc2N+4NTELTR80XjJUAL08C/WCyufC5AiS//NRv
GA4nJRxGPsO2nsX5tEgQHul9jpJ7VooyGqcPEkd75cBMJ5sjpjYvNPTlxkWmDz/ryULz3F1u+10z
InkOLqUc+Jbe+LivaDPHoKUg0nP5EriE0xfJw92We9n5nv4kvzR06XPfi0BZATzGhb1+mFalgDPz
WdxvMgu1zYHtmZcsRNGAX/7gYouuEmuixObTlwCPJo8yu1gW/FNoQWgIyA8y/YB0XGFht3OLQFZg
pi0T6RFtKlC1sAfxiG1ShpUCDmHmtcTF0Ggcam5RJB1jJ6MP2VPqjYl3uw/D7FCgH9/3njCuC6vM
1NezMfvb+ImsBXIjTMbQvusjAjvAAVMR4YwBtjE5IajXaeEewn1jGTATk8BukoMV2tC11Rx0iRgQ
jWTzxXYqNXi941xwrOnVH7rDy+nAvHQ4A3wCtN9knxM/pft2MgPTvJgfznROxB6i/WJMTFYpalh/
RFNoDIDftxEXKVIw4x02phxpUV5mjxI478lMWet6E+xb8D3AI3gyiPrPZGVzHCTBHIU0LZUty5UA
cbEURR0ykVzrBUFvKaYjscfmueYqF2ayYWzKBRK+wd+ZFWaigFqWqyIRPgU4LdtHubKi4pyYsQ/S
rTQHcztiK1BZjNofDttIdoHRHEFmfiu0bnNQi0T2LfWzzI5jDtCa4o6+wVcaIvZ2QfYpByrNocjE
mBDTZD4fnEUG07XYiQC38OxS82PogcDjKANVvxnNQfn69EdCS+E2KKm7H4EbPrw+kkxYuOeKPZ/k
Zn22gWAFgoz4x96Xoq3NNDuF9LYmT1xRuvtILj2zwBoCeJXkN288GiLbeUJhYfEF87uKWexMc9Sk
fLvZ/XtM7eZd8WfVktJZ54CCLWNW2230wp4M6xkvZLgjKdtJbU/05gKjCiwRHMe65stS/6eh+pC+
U65nnufJjjTEi7Sy3yr4C2y3Iq/X7BZX5MYj8hdifm5Jbo/PANY1QxegQV9CUeDcag24TpNuwI6g
r5atlrubTUHIij9zmGXkj/evzF5zvfa4BohDTy2+/ebir5/8TDZqK6m82dFPzU+iPzQkv6jVyNnK
hYoY2E/U2tCk8e1WRYYgyQ/xImxHzEJkWdQ0KNMKZhL4QgIFsG9TlaOLrBi7sjXm7UaDqNqGQx8C
JIraXFqMhmvfB13UgAsVx6clB+uIO+cIH3gnWBhKffu6F3a2vUO28ZxgK5Fl7FRxrSS2SxsNTEaE
BJYydvtpdI4VqPp88dkup+UqxC28GopodaJ9FyXCjGeSGUBdHb9Gk6P66ddF3AmWomv8O2Z4dkWc
3Cf4WqPEefr45TTotSYi/DC9a+0/RqUG4yb4wqJ1TH4sHbyAe9cR3zSJYl76nrajWyPNH5ZXIaLV
v25hLHXJmxf7oVH6t4oao9H+rvVrHE+1RDeVJWSop6elCAwvj1ag6tRl0Xw88fjkgq9Sm/EMd/f/
RUSg8s+vspCs3+Efe8LHRWyMIV7KSOXR8xJ3Bs4AGFIrwP7tlGI2QaelhQuikphdOfmr8GNwNG1m
KlhUNXX6dNT8r3DFQMjPZOvGnJOnpVgv6qHf63Dp98Rp84DqDfFyIeRbMSZc5hVVsZUReIp0KAAV
rhHwrxof8UMK6G6zznE/3PaxcyvuLywnjIWvA09+MpX7E5NSfaROyclrwhgGxDfgw7P3/5+vTKTC
fYahQzJdcyHXieyR2/s7OsnSx7cx8VbJh0g+b7lXW0xOTFeMjXbdPFaa38EZO1h6eEhBgXr72SwR
5o4iXjMJ0ywFsrXAIFmy7FbAOoyV2NM9lqS7qyqvnL564glQsZpzLRw1F3xBE0WrecGwAMLwfu/V
Qbh/ATfRTFx8RP4nzNSAgRjQ5UCQ4KMUEjhDran3OaRm7+S/W6pWl7XDkHTtDKLeleplYfq+Bz4W
ruKVR6NKoSdNeq5ZGfx8aEChY4IquDzcmP0TriNkfSvZfw+ZPVEniwRj/YBtI0OvrMBf+0fWK6yA
HxjbL4p8g5LF6VLzIICsaOLy3yOSOO9iyLaPeYbSdNs3zqnH6UKDHJkM5GZZWKN4XclGkh37suYI
TEd0uJPGy6oTlIv9DStD9i8JCzqG6lnipLnD9PjouQO5CWgti58TXhyTlUJaFT4fDYUXnrl2tRsg
bB6zuRkYfwhYrGs+idjGS/3y8CIC+EiYBLCWz0G1fpqikR6jbLgaM6VliwtZPwliFYGyv+ZhH7yb
01PQSlHUEqJdXIUbEjDuzDb6adJpGSPOBuoVkPJ+dg/K4r7FsHboYoArWnm8nmeczE963MdiTFGS
zVo32L4apfCNbM+/8X/U+3vNm8CqNqd2sz9bqmhAJ+xGp30Zu5N8IxVmr2x+lfRgh4TL3XwwFa7V
mgURMcK06aKWAD8b53OE+XWXKLYLCCuQiMT5U8aRD19r1E5K3y/i1ErfFzmynscDSlCI+ezWGteW
0EfIZxRCYZMkpuIoCx/WHo0NfSYelneWW/rJxgFIz8/BoIhySHvnSbV6JIU8UEwOsBbs8x6eMfUS
pywSLmmHp907K1Iv61AY64cI8+t7oqlCknjZqdBCe+RUHHvzmBUXSP19XP5g7QPlQGRb9nbrju67
XV+6g8ZGhVH4QOQR2Aa3DRhfkMZu5mPXlEupwt0OMJjdRksrpFVXnrjycguOwgajEx1R6XJWaNhw
1+jmQkPECXcs5mNJPRvtSLFKCqUK305cIjJCoAY5vF8CCseTlTTEZZnrtZsl5tTwjf7R2yx/RwdQ
SQFJas+2tg4Ee8d3Du0+RgjId3bsup2nuvC2ZwxIA/W+3UWdZ0ekGCAzwGS/Ycm5cFs+EHEfe7qz
92IhfiwpQ2tugmc7esRj2uNq/zPgP2c7xcEjjK1obFbKLqA3ITjtWwQxeYUjC+huEBNVTA+fwebo
7LW/Z99F6m9WGhvxcu6iFlivA4lzr+1x3D2JVkagYmHL2+wBL5Hz3f2DK/qdV5Lk+ojmMjcVA4zM
2urt79TEmeOfyiGLtLyEF0bQqGnzO+7rCpr7E3S5a7gLRPUWRgX/EC4O4gWfDZ1iL4+VGWWKFoGa
P9gLIxONvPKiQ3iFp/ONZ5Cq6x2x2czdZqsdEwjBREZ9ZIbaImvxEbAaeNMX/Ut0tik/5MbR8hnc
V0WLdDBuzSfxUB7mx9jdkrWxY52NiUsTVi6lCQnMSxU7nEr+zMDaGnyFRdy3hL8mh8PXZQ7La+qy
wnszzkt5VQsf8wpAaRfzC4iJiZY/YkMHq19QWUtdTKP8rKswnetmolROhBGf82X3j6VM1kghhvwV
0ixIJICy+XWA0mdPGMORzOU5DFrlF8FcXfIsHuzdrVBDda4Xq7d3XaVDOgL9spSnluAjnKdJnLWw
lGFCZ4rIAyZ1OjmJzcNsZT1wuncvMbnfr77pweYsvHxu8ohi7ZJQy7ZCPfnl57ErPFL8HcGd/OJI
L9aXuLRGXIJ0rKqETfwWi+b00tN1lySgPepE0KMxwEyf5u4Rtmq7t5BkJoEoGdL6f0dIVwg+dJiM
jQDWIwJhn/QDO8JObHwlUaTilTQujkPWmyTCQ7uXQ00LrSPWqXaUPZn085pEhRTtk2F7H+EM2DjO
Gwka1DO/yIgfiPUWFAJ3IDgkxKJ8nPOiSKIwDxbVEWKSUKjwVSreJBMZY63uWEl/HNTl3u3QzfYG
5/UyI+7vvZGZ3K32rxY3bwpyGFeBoZef+RNQfNS3XO1tBYsCsxXZEkEOchbThP4huBhekoRrjZRz
xbpx8ZphnsVhDBa2VXn4E3KMEQo2e5kYNHZDnX5E7966cmkEzJWbxMsH5agtsids0xAjMrDjeBX2
3EKLboLy9iGms6IQfQP/9JRmDVKqbuUqbXrrHn1bniTPe4+Mz3bm7P+hprUrBemO5i9h/cIbO4GY
S6mx/kZXzLvUfW+jGYkj9agSJME8gMUuz/6tsuDuMREiBHIpTbWGmVW/aMVV+/kt+CxQXXSPLzf2
kJahEKt4FPSTo1JNjzZIPjbpSOW5iiGn82CD7K7RC9mfAw+KJ0ZBuvFYvhrNVpgf2sHb2nVTWnCW
s9nfoaiUpNPacxfLK+WbBq4GyPbx2fDIHWKK5Q85+PVQnmsPMM0FzX+gTgSSQZmMtaye+C5iDynk
XGVK5H6BOwm+Njo3o6pzSF795s3sCL6dj7NstS/3QJYlChLtFQaMLGX7MLyyTDlC+5n3BnhzqRTQ
95RB6jlAiTRk4tNRH0U5TanSHeC+QgGwhpBFa9ccXbNbPZArCpgiECG9MKcnLYKFATwSC2m2zaC6
3/i1RQmgj1Vr26nI2Ee6IT6YI/iWAh1i3lo/pR7j52u6yrWAIsOux+3x8VlnbmAwdtvmV017/LIo
+5ohxjq/g/b+X0KqU/LV9CIYFhPWwqhwjZ4FreMwz7ncUZC9CBzd5kcUD1CAfD8/YAcsFlic+ony
Iv1X+UyFg31E4x/xnEZHCGlhp1O7u1BSMDAY/0bR8Lk7roFxGRxn637udZVcndJWAij1T++/gD/Z
Vyf83oFn7QwZ6miTkRCqP1U0Y5ntMxwrh4TiPAQtS5Eh6njPPScFlWN5XWGASk5Ir2d46+clzJwV
xTjgTzt7lOcaNHt5FbsjeaRsFBs/KZ7iEHrxQHV9+lp28/bUlQErLJ1LbhVcROTaTvazfhNrLs0s
7MTe+O9Lk95CxQIhDwY+W6SQHBU0vV59XRcDmrtdiOtRxU6Qh6Krv40fWSC3LlhN5tfKEK1+gU/k
FY8/Iz0PwoY26HlnCax46t8mJGb82BDgDDAMxRYy6jBSZ+EFAbtYut2564P2AwkjbnUyXGdaLJzX
K1NKskcvACxiJ/VS0JE5sQziP1/T6sV8IlSDXP9S3nlUiBA5MiYDfF/grpbp0gHnqt5Li0dYjHpI
Hf7++GJ7dW4mNWMbYVxvzp0Ko6yM5tR5jo82k9aEAqo1rPQ/5KR4+NzE59aU+F0qsPeddOuFn+Ri
ubKMsKt11/Etl0F0Y/VrfYTjFEhaquU678I4wIQs80eJL8uJlwiSThnw463Rt6M2AkvZr1zdikVA
y4wAhpBwL6ZPT4D+jD5RP/kD9d97kGaFwMMZG3SJX5+SWwM4lmuTZSD1srimFjiyKUF1bJBQZr+5
QUg5uk5tPdiLj47QA8K3Bb8aKxk5Yv1cI6HOpFpSaWuv/3S/0ShtV5mdd/WwlXeJa1rRolxFhmUK
gqrd7Dc4/maxmN0uI4jQDHC90DieJn/gbBhzdwW0Imd4JQIpmnNFgpg/j28X0M9QlCn2iJKOni/k
hd1z20h9WZJ1BJt6yocrusE7svF+vA/T+eVrrT+x4gPjMLolhB/hAQ6m34JzZKivD4SfuOVJhDQ+
EPN3pRIRYTdkHAlsASRPyEHFrpx8bin1hcZbBH+eZ+i6MDnZgtXc2Zt5ugZ0G8MxXSObC4zknFCT
SBZkWQi0FBGKLoF7pVLK9mAHgKLefJncuTJ0hoEUev1T/cw8PxKoAmtuGzu9q9p89ClqTPODsknf
TpwIZkaB6AKD2KDheAxz70P/xvo7ymkc/vG8fQvc4vl1F957e3ngXYymxgR2A1/EFDuYjpGNLzZt
Mcv6fjC3qz98tGDKS4wFMjSNxh7GKv1Kus2/GnoPt0vgRTCQYHploavytVn74nhgqm6nPOEn3aoD
rgizq6ZPNvvMLemhHmDpDjOp4o4tRr4C7N5jSQ8GJNPubiFQ/4g2GSdB1ISIxtUz/EpDcG+sMmDz
uCypUZ/87jykDrjoXTpatw90rI6d5a4JIgCkONHVESv69R0aQYwq40GDcyxI51Eo99i7mWYSgJF4
ippR2fkeTB/sg21L2fYAmZEaV0XqbaxRb9OkwB8LW2H6SeKNi6OIs3tkZykQJSn0CxlsHESMBiGQ
iHFsibjmDqGfAbb5vq6VkWIUdAOXEoY+lE+FiE+IMRIPu6iMnxLjlCqoc8CikOP0mJR/dRf0az/f
o0IFgsuwBe2Sz2c6OlhwraozHjDrNkxaqENQjTvBqLBjkTFi9tY7+KL1PrqqSwtvBfqPSduvW0PI
KpBpZS6/rIkrSgTHar4ck9DJwTLG8RKkphb78Wl9UyDn/IWy6X+fmwBw+dnT8HV23FZhkEaV94lA
k00CPoTVImStt68YN4qQMsfn+LU0wVNQUvYur7bAAcs6EgjXXthnrcC/XR4vq2xdb5eoWmAr4CLV
UKYrCVDAovMPliwu8ruondsXpUqxsdBg6+jCvnVO6TtCZ1PPbEiZHvqrxCjDG6WOZp7g6v6ibwla
cq1qBXMvUf3FxavHDuv6MSXwbJyRHm2eOD2+41psLuyoqGIQroOAjnuxAf8PU/sgZ94Ph29TLutI
Bt5/VbOjmWDWOPeLOw1YqIei7hiHD4QCNoByS3BKuwAwECuizJKcEbobOwFWmfBVCGcm4HAdJn4G
n9odNmOgr8qT6/rFa8jPIGgUfeMUGnF/Uxa87y9OXgBBYsJ+ld3nM0EG7ubkHcz8jDPhIhPtmQ6a
HiuDJX6PayFXREnO8VnywexUhxRkBxR5W88DVBXpSEbYDYfbcEFoBfuykN3SWIUrCMtHranTWWld
FIXf0Kz3EY8V4MXaPdhNRqdXjatk/bQqXA7om5BHvPp+SUx0WbxS/D05LOfWu4sL4tngk9s16HXS
S9IB7Zz2f4t4l6QBVzuHBthEooRHB9MGTeKv9KCxNRP00hC9woMZ5LwwkRQ50MGPRg0vP4PcTx7j
sXFIL1T9qF3R88CvqdOw8XInhQ0mzIbZ+FPeLYqsPINiyH19ZhZm+qRbemKLvoRtNmzTbS0t7h66
0jluKl02wmWP5ubwgpN25BNq2fheWB9zAO1TAQltziFR0AIGm3wJZ+qtCk1JiXtzkmYqOjXPLMo4
25Zrlgbpp4sWXmSQ0mFOqAI0sizTzf/9TbNxjCe1woL7jlG24tw2WBaOJWHZrWFrE0KYDeZbStT4
AAFdAK6tdnF6aFvR1fcNrvcuomoJgaOLf6m7zss636oZ4KDKxgU9pkuaF09oaUtuaHnd5R22G04c
P64NOsE6cyzIckE+8tgtH4AxOgSLcfzb5aommciytF0f7JmVmK0qWOZPWVrCKMm7nYYjm0kipATp
zMr9SfzlNn++ZL4Eq93IIRuNxHm2WshSdRqLFksKSPtSVqo2imB0463gNG2tuVq4ra/W6oe+159G
I/RylXk8UGQBR2Ej3rlUjUOLPMoWWCxHE1+7sIRm3yBKtqWDAuv3D4yH1AfPA4FY2lVX2FvLLxG3
3RHUvqPI+eVINiDBWDT0CstvvJPglcCB8TW8E6zkYHdj+R7g/KZmMBcFgLhNG/suUBy7F2v28Ucg
jkJMpzCBTDU6Ifl7rDP111TyxMwaElFQv6SyjQ7pC19Mq+iOLuBFiOEKqTimQsJqwzQuxcms2tt4
OL7g2t4ex4E/lvlcF90Uqd8aDofoJxW6ABbXBirffpRkplmxRGejd0mvzbXrY8X79tERIyJR4T98
ab6eEfx3czcftlTf/4mZsMPHeppqGSy1s6lhOCZTXD0mPiqizCCtVE2s1D4gFt7GX3nC0paGHEXw
hRKGxjOLBd9H8/5+lzjALe9MOoY57vqZGyKzonyXRjOgpp2I2YM3f1MJyyL4SUkKdQT5b/vWYJie
Ijo9owAtJCv/hZWY5jfK04pn0xrr1PWtM2vLsXYI6gLQeOygPtTLdkKKwFiz7+XcUmicCSB5GLpJ
lrznE2FsLV2R13BIqPHq1XezwxfQCnMTI1gUBLB5SO1A82D/LoapSari71tJKdj2BPy2q1n3az8j
YO/w9nxdXFuKIqj+4WoqX1Q2I/wwKzGDG8Ve5xoFpbiwbgVC5Ok13yTX2n/4SC/hNlhyd8pSrNVN
g3bt5fxugK2DkXJNaPdcVlUU4B801jHh3R9/96ororelBk/ET1n7gNFJe/IKQXBJddBPKL38WPQx
rEzKQ7m2o/tnyP9gbe87JGAcfY+S5FdgTtzxr+hovEDXf1IKa/zwMsSywnPC0fc9RN/cuvg4DGvW
NtczcTIstlIImTLs1OG4zI8X1FGvkxfDVMA6CB8ILn1uqyZrf3wiShceUUHL3xI+3L6+dvtTQtgW
NPZF2FpW5qUId6870sS0/v5KdRrdm0vwwpd6FySVvVEXtIaArVoU/PIV+Gm4d4nMbSQKwT6quT0/
LGBDyP1av7bv0Qv7UrwnYtBU9XEz2zysN23NCIpcQyolkN3eV5F1zQGzjamTkWCG4kUS84tC4NmT
oKPgHdwEfuBJjWKdXEt4pCNmn7C/P2QYKB+b5I3mjbCnOwAbcYEu2PjqUjRkiu0LlFosiNLlUU1Z
giyB1lB9KGIbAqdm6vizH0ojbAVkCRUXJoR3ppq1ZxIEkvrus2vwKkBiB/2joo5ztqpmoRsetdxG
+jSRstqbcZIyrS1rVv9k6VufqwoHAfBuTvgDTBUnWbOP5167dNGMg/szgE+ADSHi1ZxbWXj2vruv
YeWF/Q7B7AbuC03s0vu5MQfCarQ8CAk5mh4nS44nbVwopLQR0KTg66tI+lAf790wDc0S/fWE+1gh
t7ZPnSdNbfnGsAQIfTluv/tqzz0ktqZvsJab4cRDR2TKjLxUpHrI/29QlSLdbrriBedlawUHa0PL
AC4JbUh+y9Hn3eqlJuHI+UOIdap52WjJGUF322wkqK7qAur7vdeoBdliy9/JdnQZ+MSTcEir7WZU
+NzwTFSNnkT5XF36/YtDTTWrvk+L85/+ptYdyIfsE3a5GNdrwjFhm55TxZipjev1afwvJM+rK/Ch
NOKJHrfOcl+m9pQyM2NN9yWy9fXm9fbQqPMAKjJJ0gy4p1LLgQLXgbPHF55yhIHpInZCOIS1B3rC
B7L3uKlSMJ9nzoFcBhe8DtPn3IkEK7jblBkgrLG1TOsW7sdIueh2I/k62QTLBE/20k/s9RNXuBrK
pouY7qPSvTtQi/KsF5AYjK4Fqkf30BJ9mJ94yYPDsfnnmO5cPtYRdLf9wLGv3+EuBYOJrJds56xy
BNcUHk9A7U1vA6d/McieCNOxYjYL5Khgim0wAphYp/EYLXjRQbvyuRZBEGLW5vgofjSXlqgQiVb2
rOTlojGSQZoeEG1t6z8oayWOflnF2bGX/UVblNFsNycrcQPnxu5arHURkEwBeMPFb6CVpby29ASf
sdUgu2WV0Si4OfiCdGGzJD8yEI5PM98m48CWyIcwIMcq6tlsA4ngY2BjFN7X9kvh+crqxak5pom0
pUHI5hYUbErNlgqZPGstzPcscLjIpV1mUXMsn0Tqu4M6n9PbZMrg1xcnFw3V1tdUw2VA0ADxPRHS
zFbzl0FY0UymQwTPTjxZR33MX5H60kNlq3HybVlmGLLwncq0tCKeWfTnysg8D+kzsGiIwn2/e1ES
mQyRV19K6DnjgOvNroP/TmK/gHcp6e2Aw4elr/OuziuA7dv6nkdJo2YPc1yC1HjOVd54pXqcsqdp
esUOQak9rxu87Hb9uBTGrZsHryk0BNypcEJ86rMIYdj29ni8OYlzRdxmmkJECDA2hMJsdv4SRKYX
ScueQz3VTuFla75Wz9I19lyDA9gDdiz9oQ16pe1f5UU/fSJquZU1DJ2g8HK61Ze3hJ1kXxvFOIOV
2UTvooZcMNwSy9DBFN1QROCqpkqds/hr5sLCiWY7WIEMPyuBlUToI2JbGL37UEobzbolNxehE1SC
dyQimY3K5uxaq1Xih25xuDpW+tIB9bqf4jPgnX6QUQNF/TU/o51jUvN6zBdoUsvQBligVCM3XSfE
CEfHgmHvPnUPskCjKSxG2yWCq2AkEoNppaIAJGYiaGDYqRYvMqZkg4RZB7NgfouN/FMJkN3urofy
pC0s5A+XRAGTKV/h8cvbP5fPnMCzdchpDBZ+B5NTR1xkcc7o6W0tSe3g6FtFaUJU4hPveMYqJDOj
fNt8S/y64jmS8atxQtyl59XyB8HkNXe0XB9A9iCPNQMPuY5UvPCpcKLXyPW+utlK9hNu0Du3Rimq
/ZfknGi8XKklJpDVlJISvsYgIq9usVz2k4QanVtSMHgaA1tX5cq7J8nC8r7i6QLnCXHe48aU7uNs
iXtf/YlCJDjbtX0h5d9qdrtugbZ4GTzcUZ48gHGNPm1a84WdTxhjpbdBzMTR/HmWzgNP/u4Pvqd6
VzMBhc4BvyxmyQU4PFLPgR2Z61wamePeFzMhfZ/th6cczTdY2wiY2qmbdMPlEkcGEC7w+lTE8FMR
eNr5mi8JD5YfMNj0918RVNru1Il7zpsMSWGHrM60LzIxSjKjDd6JnX7V09Nxgdu4MFt1Z6mMVkGq
GPi/VXLFqT6i2L0H+eNP0jRf8eZKeSpBwZ7IuVRVUU1Muu/mY4VbbmeXefIH2XcMUugL2eHqIWNB
uwGqY0x73WQCrY30BBK9DR3SI0lrlzEYePQ80TPvtHBJgO0/thbFue3Udov7ZMW0yGuqYEb0/rH+
puNPFqGo7wj8sV/Lz+t4gfGALw0PK76HcMXndQRR44a1pC1nWIn9oywZ7xe4GNzR1+2i28fDoDR5
N564+qGU55L1KCp2JZI7B1dvQFbDfhNd0BosVbUKLbJFLEGx598iANk9oPsyi3Zi+8XjOY7vZdoa
2jvdr9UkIRmafXEPWkJAMh8OXRbIc5IS6G7ezLytT9915+tkbI8N+EvEgLYee5AdQNIIDpUYU8Ml
LUzHWxBacNLtqAPPishQQXWhxHpA/LeYZsutLep9fTIYKq0YFoiblTRMOGLJbKI3vWnvd3uzdB2r
fAM5Tah7rg+7ATaqGcHg7utjkT+alNDfhRED04hhh7ww9B8Xp/h0J7uoJsu5HMUfyEMvZt5fUqs8
wCGZ5Q+maG1aoZE98KDKGYeSUERQ+tnXtG6D4BbgKePOsR4jdUGmLCdo8/MsCTrJwae6teE6+w3C
ePD1ZHpCTyXn7f9kEpU8RQxERaU/zIW2/0LIeDgVCKw24Qsxx0e3q2bSaToQh2wP/Et/7eUWq2on
xOOj3EmM8VUvY2Djas8OnNvAhOgB6QCdIM7/T636oljnh9qnt0eZDfV5yOOnSfU3GY4mDdzss5Ck
SvZWNKDSMkz4MVH70koH9DFmFVQOs6RrzhokMj0AUJ7WIXiUvvz0/XjxLbZ2RhKEwt+2qkllWAqC
f1k6GL1eGkhSHFfdAiKih/9GWu6E50UP6z1JZljNiru6z+Sr0rTABnLZKbfBg7slvawsqEm4KHGf
bT4mlExKOyUI2aD7GQXIiFiHLxdZfHGdpj/Wvt6Eehbh3kro3zr352BEmvMXLCanQCpfNXuCbQXr
ZfthdGORHG25Lsxx4q8tDhGpNAusI1hi43rIfU6uwAX6NxV9Sn0Nxq6mydLXUW9tZW+RbdsQ4FAa
nLw3RnKldO2W0KkY/IRHDRtqG8ptYSbT4G5CU2yDJTg4zuw9uFZ9B45NSUZmh4nDm5u79DgmgJ9w
xjJAB8gQel11ehg6JVueMNYXFo8cEQsgGStu4wyy3UOBoH6XyABV3UI9FmL0sjhpZjG7UCW9yts0
Dq9Q5x5AZbEiojpbZsDN7AfRI/oYyInf0V4Glo+Y1y8/iFGqmE9xmWk/3nl8Rl2eKJiARhEXBr5N
Xmp4ot9aKHAMDzRKUH/GFoCM3PGGm/P63x62FpqghB6sVeq/eHqNLrEzq6wpM+ALWQF8cC+30Vt5
iFe6K0ijRYhSjocRfDrsewYI097w/KITpDktbbuMUpTMUaT3nwCaR4Cu45nq0aSjOlCN1QNZCG6E
SaR2uE+dz42mhWZfsdfdwOB4XsoOElxegRzq3gOPh9YQRBDYUIiLlZHk3uImYO7bUxD+uvaXMpgZ
23nHmavWFUC6yal5ie3xqPaIOYJ2heAjoQ+UCahanhrkSUWyRNjhFZSXi2Fp8VYP8OLV1OY1BhN3
lFrDvpJnaqsCtS5qNjYmjJFBspF2FKBdZWZe/QfiBpSELcMRfSAtP2nnKuHjHzNgEuBI09u7vObH
vXfpOE5E8houl3P5jM5fjTSIWD1S6t9fiHHKzpBorFr658irJfWgicFS9msUUbc9Qgi97PG2EYRe
NighBy8hlrVQcz0WiwZmREezZ3e69Ud/5OclX98Xz3/PxNQBzYaF4bDIXzmz0JacHfpiX+BiduEn
q/1ek14LkBrwObKPbdWLeqpaur01WDI230boGvLS8vvMrm2X2flc/yTG1J9EQQtYB0tWvKVjZPX4
LseHdyyHB6Ool+tFayCYQ9awJjz9Xu0jjeIR+UlgPO8s5s+qpVQOZpQgqT3JEOoU9FQeozcRb75L
JnjlDebWZ+rt7Hocl/LAldWVK6YstZFpV6Tjba7PlV09I3BTYw/mIpLyYqMqfxjpbc5WTI76ovlI
EonMDOIxBQ0npIOCtSp8JbcMrZrn8BEyNyBnUb/E5MPs8eTFAGRw2l4QgxhP7FQHSMxI25UIHD0t
GJMktXMYNO+UIrM2V4l5OKX+oUnbZWZH5T8fb/IoW3Z9w4uTooBoo7S0EGnilFvIAl9epGROc/Iw
tQznJgOd80XyAr7XlSJAW8B0owjrWSC09VekTks+pRR56gtthhkLgfsqOqidiQ715Ex7fv3a5Caq
5d1gUk2F9ubLniepHqBT6lQtSMSrXMOCg+imrxk5WNhyQE3K7HG+KkQogAwAXYJuunRUaZduZfUC
Wir4IkfCuzcAuT0cddcB7pQJm+24t/5A+yjDivWv9q9P/Y17PtqcsIGZKYyXPRZu8L/WlF9pzFIW
EMbteu4j6HlN50FLMytFA5VggjLjpTMjj1HgdytbZAuNSqXZLp/6rm2dg7I90hAYpvVmVGQwC2nu
/X7puPFKr4vV124MyVhrH02Pv4WpdEXAEp72no3bck57YtyErgGf5X8cAJNcU2EdbR4oVyfSOvGh
MiD779/vP5GYJnaG7c+c2skTCD3Q3W/Hirhr3Jnfbhtu/ErE1yk5nYagF7Kc7eVwTYh5KQ1mgPmw
wbSyiEDZrohNh/yBUeKn1h34/TK2vQ8lXh1VaghPvloEM4Pi8q1Ejlz37ExrA10cImncrDmm1eU+
OPSGU3iJZTX30Q2UqOL7ZaBLfDgJlhj6W1SjFTlKkfJwmHqgX+03dcoRzNGhyWziNfBjDs4m5YSy
Z69xIjM9CEwvgkAftB2hokfAYav6EZpemmTgp0pnbCALU/SPVuNm9e/m7OzcQujkw3AqRPWmypIA
qHhA7f9qp2embIfeO5yOLmDiSbLi/e/87Lk33rh4kCekcdQBeHMYq7eLlgumAkSWZ5y8WiWCoAfZ
RXI3ln4VainTvOTDbLmTr9YrFH09/52kUCeFXwZeffrjXRHTjSNKC7PN9wu4AQeGOtpoQuMhSTaK
/SDmOpzwamEMHuUg6CNCrU75bb42IRwgr8av8U2pKO7ib+q4Z2/nAVxvjryxh7vQwhiu1MBRSc/0
76J3ZBFci8R0ORJ5vlYXCVrsachdi9zACUKapEyNTw3kQ4GHQ09Vys8S+NIgRp/RXDcM/owKldiX
ZjW6iiJPYiTN/IsGoWlDs2CqA9vFebdUTL10N/jfZIsqEHZHI9nkzVSIhHDVoim88gtkKczvRc9Z
RC3MuMXTnBPzDZss6a7Sz4eFnpb+4vb0TCkJbKPNEN2NR+EgNRBWiNuls043EOou5Mr6/Sf3sMLt
1h2l3bOUlUSapiZEIFdtFNISWm/z9XZRSkFtaealukvYhOzTwtPJDk/+533Wpb96KriPcDuJFW25
sqMZgCHXv7LkVWlAt3bNE2M8/BRhH8H8VBpGfblWulMmoiVg7Lpa74ta6gYXA+WSV7eRD+N6dsBW
3aNA8Ud9zWdztyI+StWJtr+4JLwkAtyWqQqnAvjMA60XPnLCTOMT3rpl515jdO16KeGNBH0h4mM4
TxXiWIbtlmueyA4zFNShlwevfeVrtAOmLRRt/VOCfTnC+JmNKs5ImjGpxCgWXzI1d2z3GGmiItmm
LQsPtE5GQdtSirG8JMPnpdwzCXp3jLpR2uHTgR1vBWJMdDO03BnIkLYU/J+M+y8EmXtasoKkQSQz
AA/uC7uyhSLORo7iOque3Hz10ArXxWhaZjra4zmiRLusJzOqQq1ZRCGya13OD5o3ABkMGGfby0LG
2iQPjk9ODDy7ysj6bVEFIvoSw0e8WqQPRPcqDhV5ZrzAiSKMOQ6x1pQMGQO4tiFAPjlmgjkbiYCw
ko3mJJE/D8u3ofEt2ipwP54S71LoNuWr9Q8ANQgvLCz/vSRXt2MD4ARII13AsaCzvDQpgj4lVW7C
dmHlf9zjaZhcAd7q+QjKbtZ7V92xf/xrFwA5pPy0eFlMUUqxz5vuY4AEmwJejlVobJ43pnipcWyD
JZ1F7RpHsu9mThhPNpThxPc02dFSs3f3q/6cIuYbuHVG145fVnhN0NdukUMGfre89xfmK0e05Cy1
HoZmPJKvdAsAVgPNiGkFuayLEmRzU0IxLWzcPJGD3MpT/pRCKrMyMrno3DtYSk1jW9RYuAfGauRH
NZuyS2hCv2D9Rs0A3mEaHmwJ/Lynd0QKDfgRum8S/jxB9yOtbWZ+ImS0fvPhO787IaFUn7fmB4BG
BVZ+zYhKk3b35En5WqG0Zzk5nQ3ez5yT6Tmy9RNLHXP/KhOOk0lzDYq8Exx+WUYyCC0cK47T3Os5
DA5RFwY6Pe5mJCA2JagdwMqZ5kALrcG7UfUFzEVnMuDScsmvmCV+dbqn2PGxcIymfvLPy8rdD1T1
+3n2sO0XNulKRDms1fitldLCIa60g+u4jxCTvcV2eUdkiG7unCImp3jbiKmjI8Xfi65IZMS3/3lk
5j6HzEKJx9DVvUybw44XksRIt8mLnzoCkjTfK1PAXR7avHllsf2Gv7+OOpwhdKbmPgHohs855Gh+
1rf58x8Excr32p8EdBE6a7PLiVtwnptSOsbXQRjcIAqQ3ZCyzG9rVfV6UE00KlFJnwaX0YHp/GLQ
oDcnV7opMVWwnu1xJcpwEZIO1web0HQJps/HcFWyhqcRmL85j83jlmgbxjEH5Q9BUzGqy4zKDqdC
elRDPQtmCHfFTxEpaAlKSEwyOmP4F3RDfirAvMTtgWK+liKXueL/QI2W/vklEmBTJ/owzl/6jJJg
Iqv8ZoD57A/omKzNACJg2XVYH4wTHCFohan0rH5FebDXMCYOi8IeWTrwALAx3BpKO8qO6V1BPp4V
Ylh71AH6aEYsYr3G+EkXYOjyxzHn7un71Ra1FMqbpNMLtKDSPrly/oCFsM1mPaIrt5BIsxCkMzmg
pHdbVxZBiUOEECpEV7q7AsBmydIAAkFKniIxZ+38OgiPdDIWUJ9wY6kh0jR1cY8UaaMUHD4/mCtn
OU5HDFKUVvGxdsPhdL24rAZjVt8p8Gy7LwAAaiFgToJFXJ/z61V3691YMBV+3hFjvPhI+YW8Hxc7
xIfrLDDy9pXWbHb/QC9o6D3sdRIm4IoNFFk8spYCG30NhzQoS/HBzxLnCV4WbhubyUvAk5QtTtZS
p80YET0IOfUdJDNnz/KsAzPezZIsBOaob19sE+9/VRQ0NJ9IZIjgBOBI9cJXrgJgHiM7yN77kjHo
+UqzsLTcFxKXUewjCfceeEfng6jc7dBP3tHHw+J3c6kQUvS6+6iiH9gq9T5am+QiewLo+0ls/nJ0
/gfi52OXvjQusoC7hcFUa1/PxMqn84KhAFLVRwvpZfrPxm98/rKRyDtgoHFTwzfCqi8HQC8HfGDh
998z6uzHq2H83EfqLYRmP9se0IyJbZcGZg4xGJcm/YAIS4shPQUYxSEhOzfWI6b2S58Hi+X5MhAp
uab4YcSLAgY5ZPa5uGKhk4GwGn6323/Pc6bSI2u6BmnexpfJC6/6JDc4OhPx6dNgeUGj+3cOn7bV
5TS0UyHKXnUtTqOgtIsTZvxgkNMxxv3WhCozzorPEXgvv16XiO48LHGXvjFFIeANGqa06Idf7HDS
83gnn3Tl4hPbhFMam2lgo77Dlccuhj35R65YUvFnH7XMH9xmcyNxvTJ7RjObQ+t646PR2WlIz5tC
7PoDzmUY5GcMQOeUReFidP+aTQgLn+xHuqVQ2Sdx0NzVPoplPrJKKJzqKPsJXVbDOnarUK3DE28d
jEseGgFxBin0ibJ+/3Sby26xNabloeqjPS+ulpsmHMAbPCCoMRvmKCT4vOOM7n79BIW5PXICAZkJ
wgLd1vv/1NyH4eN7qR5jGR+Mor3ru1LakpQIE7DYDHqGBw+EzT6DGQ5MZspMfsOzugkTycwRxys7
49zWSn5ej0Pk1ksoBjIWoD/+CHYFzKy6jC6gRj6nidv2qALaLNux/7tYRM1VYsmn+O1HLN1RJnTs
/32xYKo7aDjiK0vOO96QC3fI7dwTO1DYGckWbXqizpciiRSn6d/bT93d2tGfT7xscOoor1RDenxS
rZA5OE1J2Q/3x2kNmlos6A6XqyYsgQTwZ3gC4wMmtTvqBQbU+0OrZtYtvMVgK0bWoV1F9OCxt1RE
DlziTeTB2z4v3auk4rLdm77pBE11lsMk5aw0sCI55jpf4itVrSdKY11NfZVIvABe8U4tbxTchU8x
wqyTt8X/+QbDC1my3soE3YgfYJYBYYCj6xRCLB0KfVHDLBtKTsFe08Nr/eu63Go0G/ROMmyyy9sF
siI0qg1s7kwghxwJZEYaaTHhpLflKjpx2hwzHbSmFStQrZq8BqyUGGvbsPQt62W3yqTWSJ6w2qmB
AJbwJ7+vq0Bx/fe9AgXx390wFg15RvrQHIa/Ye4/sMxQMEbckAKwp0LW69QkXiPXKT4lfeavX3KM
DfKhu0ydeBfrgesQ7EQVE2P5qO0CC2DqlGZdNNe7bfWgZSK9FCc4zVCf+eJLxVAzzDjAW4g2XUcW
TsrIRJpQ6GdOIpwJ5bnITBdlGG52cSz6t9yljQAn5mZVgDralcLJJQYHbkrOAvOx00gWyVfHRSBV
WonpfquQTma+ib4hPTjOspkxo2RNpALb43TXYC9rvlyCGukqHhsNNRQIGz9ak5vnTkL2YAqrtswJ
1unz2ptm9QozojzoE+t26kjwRZPb15GgNIiz52RwEWdVVIPsQ9nVVD0xfjFqPXyWYiIK5TtktNhk
oTxjSKxdpfhoKzxI6O+cKjl3RkjQ3pbxiuTQLj9um364NGinOZ5E/5mywUVID39McAjdEf+oFph4
wWjWC39xoCkiu76bFeJ1muC7+ma9k0rnW4TVLe5ZfKtqaA/1pS500c8Qj5+t6+Qjnb7PktVk+1Re
A3/OrMMEdlXzaaF9/Np18lDEU/pQgdNHapHu3WS0UmcWEq/YKBeH0yI0hQLED1fOmQNpfAFNqXwg
BlFIvy2eKLnwIIFWkWQhR1N0F/ka8TeQISH/dNUD1W0h/tT00gUN+3mbK7f11TGnQbsg0eAnViKr
p8RuLqaydH3Ust4ZS9Mr0tpZh7uM4OMIqfcOHrBWe6FScXNjEEKk1kCXHqwG3wlXdSiiQzlFrAWG
5x6QfIKRIIvv5ad/+6q+cZ5cFcjQlMG3zdOe8KPOGzTQBQYjbrySpEcsmAlYSYccjjLzberTj0iT
/d7IjHIffTJmBmLnZxawH97kDEm6TFEKXnunUvSnEBEEQ6C9JRAt39NnKrWPpUh2MDYPKHOpGm6W
bAIxadWj4ZgLJtGL6cLrswzkEdx26+Mwskm0FUFkdLV03Kn+zerSsG5ghR79X3AdPLjpB1hYNVMu
jX3VswV9t2c2by2UCUDssgk0Bvo3U/Hfzn6iyGITg8R+Sxoeb8VzIOuqV/KuoilTqus3UH1lT7QD
3ZL8Gd9F2/CWwCraDVrI/9SdMY3lxNXujXpsw8DLwiEJObQtvHQNbrcKTP37UWgwfxTTPYeQmbsU
TM+q+Rr9fV//WHDxIrLWB/nisE9hLL6e4/nRbUVOpB4R5VIkxe7F4yEHG2/3SOI1I2JPqU4RW/MC
uIGKyI88u1PSild4MaepF740/xuo5JY+Hk2Yc2zs1tfaeJW/i/J4HTcoXmbQpzhGNRnCuBH4DokP
zTXy++yrwKMm9rfBtQlGOCazAUQh+SBSGTQjGRCV+9nDUL36W8fxcEd85JStCVCZnzSnL5Cz7JBT
XkTrIudxFFStO3o9n965bg5OBhLAmZhlGaQRaX7J4UcGIRV81SEj94nJUOSAY7ng8x3VDpjS3s+r
dMvhXfH0pbjiXzb0fwTKJ7iFHywdIJiHTheu2R70wfZWHBSvd4K6+n965l7kH3AC+Q2P98z7gBgt
tUpXsnoX12jsYPcJTPCkVhkqhP1OTk1r01Ug8fyKzOtWUAtyhspWV1hGZXFgjL7keqKda05qBwpo
ArU3Rc3bzBS1G7/KTuGpJmTpTPZCtycBBidwn9+PPC5hGH+cliI5lGAj+TTXjxdeTeQuHkYkMotR
UmkL4cWWtZqIBKWeXNaY3Q7AN4r9QvfFcLzs5k2fDRSE0rPylIRJBiUMBWYv1gza7mjFCCSel/hg
jyZYMSKGzCM14sUkK3BiGeUG5gihvPmBMqat+7JAWpUFbbHmVbJT7FsBvEPnTTSOmWuxGGsP5D17
jDyTuciYbNAx6forF4MV1rNt0u003ec5cynvyKGNRu5SORztUe2dGEHChR8HUW98Rrq80axiNnt8
4ExivymWp75uzTEbBbd9Qj3MKqvi+7Mip41s9hFP8AyMv9BSk0+Hg6JoyUIAii54Bc8d9iBrFFAw
2Jh8duRNKCSMsX/WOgUfzKhMTDLIsqSGPodyxsEDw0IWD5TcWesL/MnTw6bT5hP+ckUNydpbuMoa
v1mUDcMewJ7jtkZ0hBda2yzkJDE3FtbCP8en9d2Mf92y9j2Wc7vMc6lvvwcBTV2dKgfH8W5oDIUL
J4Wxf2ZbsD0ifF95LxJwV+nlLSH98cVaAY4krOj3LyUxQeuPn/8k3VztZ3ExEuXvZib9MufFp6m6
T6PdJEoed67EIAjTX0rJtaEakIWj7Vz4ynKgCCZjbQfTcO1IMPr63+0cEr5Jc7oc/3grXpNgEMx8
0QHMLyJkEskuu21BRP3/LgAyOaCO6ctxGb11sftgseXc7gsXSeoTdRTOyjrUsP2Fjd7GmNuWz7KZ
3oJidWpgLUgczxg5P9bEBq2F5WObT/6OvamfyoQa3ICVO37G6jTKKMRDuco6C7UP48RI8qiNhiqQ
d39k8LDxiHvWll9ua8HuHrGGGd/YlKvuY0sI3amTCv2c9EMcmTtQ1eqo6cjh0713G2JZadkNweMn
YXD5gGnRgIjgPyCxW9OCv9Ue/YYJHOGfzoFm5vVpdwFK/Pg0800EgKxPxlgyEyjuRVAzaTNuZUIf
2g5IcygbmDDLyPsZgq2mQIKY5204IUcAxM3tr5yDLgpHa6E52fanzFIoEY9CVHt4NW5jLmcWv0Cf
XkMepXHuZ8tkPHNrnthl1vl2ZZgAaOz8njNtptUFSA/JT+8+w7cJTExS4SxnDlVnE5m1XeOm2qOD
CRpoHFcTpjl+1FKoK+k31/M1cNogvBF+nrkQ6X6Pl6Y9EB6DFOM3lhXUNI/q/8AFlp8ObMyBvz0N
TT/0ivCidCA/Qcb9uwxty6sku747hazXDJoPudtYfPkbpi9WLMud4TY+K2hk2jSrCdh4jKUO/alM
yh5jhwEFYpIPKgIpnl3cWZlvO6EAk5yrL14gW2dVALCp5T5UcHFQdFGY5P1NMVo/2PHd2SHAjvLH
HB1PtK9992LWA+Dq6nwh7L3yl293g091GSJFTuo4tJqEAFmO2Zb8xdIcNXGjsy2SEJYfO6qvDmmx
NlDAGOsrbzuuG2SK6IEUmjPXYzQJlFUavF1gMwt8R20b6D1/WWSM31KPrNk1LCfJY+d6qCzAKgb3
BkmTl3yDtNJuxqAmmQH5BIDxg06F4NwrrTrySF36Flc0Q7U42dTCoi9bmF+i7rm+ZobiePHBNTIm
NGhOv+49l6Q0wul0fwRFBP94imN57wa0vE6Sj6Qbn9Cs9goL6VpMDel59GKVo+lIBuGatxAvodPN
GZFhblhhkmCEVq3MtxPBt18ur2IfWVZ2GL4IvEIVbeq9NbHhXDXHQPbJLUbmXgXNK8PR5BLngek6
3zU8/UFpWcn4uHg6zlbUmTc6S9RpUESJY94RVZiAK49TZ08KNlN/7I4rT2PqsJniapZe6tZHWUAZ
E6pLudvP4Fy15yBka/823/M04NzFjy44b0v30hhhc+V5LtdLZEJ+LFHPdjOt8l/Am26pVCZLcYe0
jnJbWV47ovIdsLTLakE46OiL01fu5LTczRp5BvooI1bcapZuqhzV9M1tEb+oVHhdFENqCg7vh26t
8zSQd+JdROPgzXqYWfgmuHTn3kAF62KrlmoybFk1Me5CtfoMDEewvGZ8J7hCsyjUC4nRIWgFzufj
omn+k+6tn2TGAn2iZFfhEnops1QGvf4n46WzX/Nd3K7jptcOspR1THdu2MwVa01U2LhxYoioE8Ou
t0NFdydmFd2c9uS12BGwqIiMX1Fp4faKB/Vu/uj6UB/MSnt1+QaSBwS3bUfLMgaiU69VsyJ+J0ec
BGoeWPhG3oasdLtVKdh/oy80cg7gCQwE6DOLC8pzLVfxuSbksNHmGwDCktZMMkpiMQ3+lc9hkrsu
zOw/lh8ezyuMQOALgiS/HaA46hvpV9YNzqokHAe9+7d4KOVH7onFsaoTeH2Ab0SjITchkIg1whB/
0YqewcOt//MGjaWDArDWFqytf1OqN8U1KSIvqQfQOSmI+hx6V89W3TMq4SfwVLYw0JlbFzmUpeSH
wG1k0tF3/J2Xv6Cd/hTUabXtK9MKafR54PWCapevBj0XS+rM4Zqn1/+M2rEJ+XKyT3bqG1VvyX15
3BaulGbJWTyzJmLjU5JC/jqoYWpYR8pYDUM+6AYOmLnwEKG2WjCHt00hA7fBNFgv5F0L1ZWMVUNU
eLeb8TZu30PshsoahMSQNfoWvRyywH503UKsO3EKuCKfkCbsGEPtsjB2wetpscvBJ4rnuZ0OMGNy
kzlULKcm50dZoBM9Fxb/iYs8MsB31uQA20IwXLa8zljVpbQ/OtGGRc4psItkPcslNh4RZrGeACfw
mmEJ1LPBc84JSv0YjjLLtqk3s56CEdlWA6DYNStl7kTBtr9EtI36ezKBdpfOuIArl45wRzScqEu+
+fcsO0spsG/erzLWMMMMo2l0j0awAu+zJhvVqG/ROizNiTerENV8Yp+LgMLQzgv2c8unRAV6ItCU
4JIBaxlorDd8w8bH90Fb8JLYjgILAlAoBzN+RsZR3W/9T/rqo2ytuRWyq5cYMEfxJ+2Y95UtKro4
vkd2qQGh0w0i6mJpy3oiRurTaOt6n2UjZSdxnJ/b4Yj7auY38+UfMkCxhPVlc3/Njjsuta15dBZl
wmt5usIX2oEiNRag7bczT+tNHrRtKSC+rByJUQJOrLz1bV5aRanmuF5wJs+WIZkoEliG8XBtDUKv
tic11g1gxOS+Jr9/sVzOU3WvfxZ5pf//xtxhhXigkhR52yMk2OqrmKmKM72afs2hqUVPvZP6G3Q3
LKOf/npZ1SWOXnuwtsbhNrxhzDm5+OndXapIo4PrPUoz4G7yaTH53LQg+revKrMAuYgFItg3c5md
xo24N9ULWhup59vz1qAHZwEt3sJS9weRdrCOX/z52YWzIXPmfTwVlKLHtSmfvnZaUdgbt9AXtc9o
nDi7sogmAkj28E/VJgDdetrIj6jCZrmj95ZDBVVnV2kIqb9OFwBzyqq40qT7/GFlJwa7VfWx09yA
QFZkCpL4RRiVm8gdViAUpid0NlGqCMO6yli6Cg2C0+aDsnB1+qa0+ds2rfUkuHTzdmzwG/Hft8Ur
yWSv6hXu2dTG3vqwcsnf1cqRclRd89F5LP/Pf+G6eXj1/WXVmZlq+u6DT85nGI3JQJaQJfgwIECw
dhhwoOatSuV45PSqx3gzjCD27aDv39n31QHHalUZm/42tQQ1gHzL1SvLhRnzkvjZ8A89QXbHfAQP
DQS/Ef5xyaIkPUDpm+nZS24BX5y5zgYTnJeY8rZn/Jdzh9x8bgYPe+MaAgP3ulIikyXtOjeRp2Ob
W/KG1NTdaAzR0enfHKU+ZYoZ9KghzUErSOAK6UZbHuDFrxS9iPED5+E5vAItWS772bXoStZ+xkn1
YtUeGFFqerhFoCpuiNt9cGfPLmWd5qnUaeREWt/mfYgjca9kMeotPYh12SENqhc7BLbX0UwOYZmE
EKh29cw8PT31MR/7CnDVzO2/StV6QnIg5D8cz/WbAWUlDplSo0G1hg7UmPzVwJSWehnwZpj0rNRI
bQ/Thum54JVTJ72IgwBZY0nL3snP4BKgiCL/VSCCF48FCpxzK07CX4yMbBTC9xDMLe2Q4cdvgo9Y
vFJVhBwpl8E/4GdDo+OQ4u2R3IR1Vn1jxoAZP3LMCRoJNxjzxRkjNbqrLMoiRck4Qlk/+RN33fVg
P1Bx+QHTTQzkWqAL0kjDDW4zohVDR3O9pimqzukfJdNy5UYKc4g1sLAWKU9t8FHpT7KpqTO4B+vs
BDnAyig3wnRoY+/RbiWRf945SJJ6rSkQZ1THEFFqS0F2TwlkuYm5AwF86tre/NjNvmkYGMT+1dyo
DgxtfzqgAAfWGTcsECtAnQLlZlnjX/Tbs9+9ZTRyskGcI6M94DS6PcobD4vZlmSzH38H0FDbs/qL
/rYiN+LkXYEuPUqR+BGOHrvx4w0DbfbFY9JRXYYyDiPZfXsoQmNqleYgz87zrBQoe+c3AE1ho07S
cBFbrSVmNsQLtmAJVf1d1ysmoiSKtRBikYvpG7B0Po9aZ0O3WPKSngKXM3ehQKx4f2PC/HihmRvP
wZkayJvjbQUGEWaOSBB8E9oXHY9vSRv/nsyHa/lMxu2rfyr7xE6RaXzEn28eWK/dm1pdv7uGkjwF
+VQ/3DaBGrptR7BNcejckjzfLmJRsEPiRY/VECdbw8l8+NGfauu6rzQCdvxak3MEu4+TnrpYte1+
aegp9D5HsXyvojBlpoLoScOk4VjxQj14D/vZiWjjkJaUn9/aGRPOXfVudSYFlwXeINNRv/asZ7VJ
vHHnilnI2xm6dxbHVqTZF9/aGqyo+LCZWFFgbzLgSoiu4T0CDUTw9tl12vPuKUdTAKwwxunbC/zq
tK9LmT3koe+ylFACs8cq9RN+ZVetjdn+o3Bcw4k06KoVIMxmDwIyXKYiXvN1u60VPBF5vIBaZkWO
mui6Papbvv5OC3H9GdHcB4zajH2CQSCr34gTNZ7hlH+QhhFeSSvmT14kn0tgPFrVo1+NDDj7mTt6
/Xgi9EoUkC2V5M9dD9IfbCbOJw62B+jULJxZiflsNA88NmvwezK9Og9DrQJMFqfZHU5vwFlVry7s
ceGnUsQHxzzl95vmfdKGlCaD+/MEhPZ5H08HdGthJjB9HQW2WQyM86I5GioCQFvzj3TgBziwtoiQ
mw5sDXwRukuAWmmkfMpTsLYe9jjYw7iYJoSWwMoch1dylBUdhGmKkBzzphFApreJuGeS8yz5dLdL
sxg/RbVkJ5VqQ8XD7MudEJINKIXPobmb3GCXusqSe8b4ZY2GvA+i4wC+Uk42Ss/rYS6vOlIuvCXZ
tvlmPlQ4w5iHkgGteqigRP72M19q6Vx+jwYRtnoLSIPUaaq0FnmZI8v9rKhgav9R8eMit64PP4bv
T/eE4tQLpC70xWxbOK9BWvu1Hwn7eOa42CKGjKt6GWgZKUgN8T3b2bLmwEX1vu9b7EXYOrn1wbgA
E1VFomZD9iL61GitNejKS41mevPlq5ROm29WQzBXXQ7nAi1pZC/HLU02FfQkoarpLP/FCFggBsk6
sotZeD5puAUM26++5+r91TO522P3S55jtuiQB52xAsp9BGN7ZcL4v1agxeZM96ZPw6CuKqjNMoNZ
jmB4BR3v2EAfCzIHzgd0/EhVXnD+wpSqp8V8zQWVgZdSzw51ZT49YV5nTSSDHFPpcvSTsAmCbwMo
4IKsIkaqDDutzdqkLUk+PsuS97zeBGgAtaPv1xg5E01kh7UJOZRZq415Mt9xB5VPZMH2qXVDILCE
K/OgNx8RTKnvVpaj8f3g/u969kkNxPpLTlwbEGucGfvu3PhNYa9Y3sG7rk5CjSuXnXO8io+rnDSt
dguTEfOVpfOj27fzwDf61I9NWk+dacCOlHCMO4Sm1Vhut6zpFUwwkgfni6sQsT1dkT2UycFygob4
6WWQxWOT/LLvYEig44D2cWesPIJYWBjVOUB/P25n7zGp3XBY6X+vOtC5B9UgUDcvp+MJZ3kCJGtF
btywnqHr9MAQAa4cn0Y3BLw3iSLh/jNgo+79w9MDnsz2ZXBuGnu+rsWf8aQirIcqxW2Az1fYrWoG
AuJQK+7pCVIlKddUnUfAK3POa1yKORVgud1usQN9Y3+7ghXOPSlHMKWo2CzdysOhvzWdPjDBQN8E
hcMXjmaHnBFpDNzSEN0+btiVBm0ncOxGbuzrGi96rxqDJYijVDdYCoH3tOZEtRaCtphk+GFxbKcH
20aOGq3AAMkb5F1AQgOdYXtwsYZV0YeBj8QC0Aj/qPOfWZU191FovMbu80VvnQ5+109IcMwmxvXR
qqrArPm5talPy6mR0M7M/IKqw9vCtlWs7GRcEP59AfpVWQQ5IxisFKVpNH2Ts7ULfS+C4xid5Wri
vhGv+x0HnKUCGBaNURfrW4YQl3k48eCphtJtTSz/enmliC/dntU1Gp8pP8HMyeLaNtg1rEgmO163
vu5lC9RuZASEd9lWK/PQWaHRFPnEuXaPx6+ymr06Ct4R2uWNxrdLeDASlEDNcnXXXfllxv0z1iof
2zDz8jMWICXjFlv5XLOQ8eEhJRDKv9fV9b9fKDOTBINH6HpMcI+6cty7/rFbUnp/2ar4Q2hS9FCt
XMK9Yd3qeUCJW7/iqpdL9kVG+BPPnAvoFxhZfQKK0mYcNFrZUydfEcUgSJu8eLZZOxQNJkRyLmfO
C+ok2HQZbJUVfVS1kYlBlpwAAtLTQ2dBy0nQZkovx3LrNBMx4Ss9Dnq8ITvxuedx97iklUFvWGmL
QtKwLMTiab1FRM/7kEHs6Dgd4K1J7YW9kxeEClnHdvtuPNa3X2rLe4nNCCBVGp0IOkApqvYVgVtD
0XLmGHUonULg2f5GzyGxCT5aCRqeWj72pOnPXmddhcWhd2v4xdLjinShACTi/V/8O+myB3wgW3wl
TdLnfAyCEaWABJ1HGjhIk9VTUa2Ig8j5W36EIvkwYd/x+YmOxCh+oxW5m0dFnx0RTT3r2UGczXO0
Nge4GHa8netV8WYzE4hVtwfibwVLKtsZakq9vGapKm4M4g053ppntLyTTfD8omzbi1o0/bAi1uFj
eMBUC/e3hmmr/ti1lhyLIUoJeHTgPQzHDrdkO+TWGQ+uoyFkOCUTYFrwuK4EZcj9FyXPAyX+HmJK
0PEsk3eP12KNjHQHX1IlWPG44PN9bKL3rAkoidBc8g8skiUifQMNOIEFS1mL2VOjKYVnspUtDGui
otJiZHIu7I0gMymIjty3xr1n5VDI2GPmz7Ld/cVyyMimgSXV4Xc8yg/sA5b0LH3PQY0EANlXG3Nq
+whBz8Sc9VRdawT+dB6Hia8KSFuVBuEDwzv3PoJkDqyLCoX2XVbKBQymLap+el/jd7zIll59e4FG
D8iX7Tl19R7pv+MTTqR3D4wPpiY6CoHIZft0/WmMHTZK9gGvP1aVkerSlBnzqC6lxcFMOa2KIXff
rqpwZtqwGCg7pnWXjRKe7+QLfbAtuQXU7Tn4z2wvewsT6hVxjJN+6PBaQLNkQXjV8UvFkXp17+78
8RMKgNkf42Q4DInlx2Efdwt9ZqlgapfnUo7mFh/poSRfK1k+2yqTsvo47IW9LVsXhdv66H4AkBUh
N76gpz2gw1sbsYwlw23vvEUl29iCShDrUjgEt3KBqnlgJnIWlWAo1glLgAafn8Cum5uQQYDyUl68
ctOfqMmTSVgmy9JhzhyCU6sf0aaSxe0eE+sZbfrbOzskLQdsabNAqk1lsxt/oQIpqmmDn3WVYOfc
W1inTptKURTG2S/evYgeNOYVnHXIPwtpTImrS8xkggrxXH7C3AkEA/1a6CwCzYDhMiBXYTiltoN/
f9PrU5q+RIefrYFZd7u+oS65WpaxYsOkRDE/5oB6ZVQoVa7GmfTcZfvegmFcuWpDqmCzjHJJhNN2
pAxVECbg1pcbntp57L7aHAvEP0zlM3heGLS7CHA3if86W9HztG9or+pGq+ERTMtxPn2KRt+CAPTV
/fDodlf8jaS/Me3w29u6sIt5WIk06nIUAsx5hwzgdIiiZ3b6HVaeBOWLqfLC0B0+2zERzozZc4LK
D/TObUacVRWaG4azPaJx8dDaAFN2D18WSq/sZupRHfuxihiwbj0FocxkN25wgu3+axtyRjKPfEXa
WfL5S3yKJsTiItr4/gsscIdqJypMQbkfds/vDmP2HSqIc6etgiG8durXtCpX8qp1Om2ujEg7/dGX
bops2mI2zPBkQnQaMmuQuq9oz5srf7QldDgzyhYtXmrwdG0YOxPYAnPCJm1z0+A1mvpnRYUyNgRq
50bQCWWmLszwXpHmL6zN/DOlN6oDzt3wuTARYMDi43IL+ZafP/85rE6e3i+x112b7rpdJlSC4VpD
8vOVFM0udAXDTcg2er+pLwsKQWLbx1lpX0WzO+oBLUTCnayHpmmePPVZTFUPXuvzDgLesh+Sp9/D
HxdHMwsKl6V+q2b/5ZNdrcL+qPZE1+OXAXrCO9wkINMJ+2Z1Djgr6y5g7S1LWA/foDofc5fRnDLR
0x94InYoRR4tiE4QJF18KFW77rlbfOCY4msNgsv5laXI7uHT2GvcDO60LQJnUum30VZvWoBY6dxU
MGn0cXqB6O0KI9YzcMijQM6hAwi5grNRP02E+88YgEYZkxpbILQDcw+953l3ZLd2EvdqA28jMzdr
zhJvO5DalvCg/0YwFcZubJ0q1Asv3CHqdLr12o9JfvChmjAl3iIQmvwt8Uk5IuwGs4PcqvzeWsYS
CNKv4GRHFdNLLoTGLi+jUm7gTeVDcLoDai1FVVkt545gxqBUonc+Ii4svDFljuzMaylZzWWMfDw0
y/diCZGuI5pF2iVtlOEAj+O+NuK5iEh6ywsJFJzKgHAKb5uqH9hjDVlJj9tqkpxXisbLamwIkjd5
TxZMK2iAW2sD3Pe2LIWXHR3gMnoCEnabiZV2ttHFNp+y/GlrpXujK07N9oldgBfxHdxZV1UD1256
F7VWL9mnAw75zLcOs5wqY4AHcJcwaYK9EEj0pLLs14DOn7fPGhlsjcME2wEK/wd8Nduy1cU700Rr
T4RlybSImXlGnAATwYLskVlbgmH53IQqGje3QqgghhSKifTChO4heWY6fP455HVkbYHaN5RrQ9aQ
a9qMCsUHe5hA1+/G8X7lrIXg9KSn6oIvGuhdP/6MSVmBsOcyhVj6sdJckS94FIgh/Yna+NyF2sG/
ghVdr8KDXqegVoq37o6nx8sBCY401fnPWeH5Wv4XWBmPlw0TRlFQZILSahPqaUfZi/r8nyGT4f7a
QcLcvWrIDkiub2o4CMH8ObwnmpCDFlmlAtpihYKRx6HybI+hjI0yxzQCA1RpsWD9fOadDC4hf8KL
T1xTRBGrpvId8ZR9pIXUga+1hDoinX0YRGcsmXfviPp6cYDk5KXLT537WvgA5rLtJ957XGHBK+U+
ZtOk5y0x3wjkxa/WF4Tp40juKOeh7BJqkAG119UCOSI4hP2U+Q71JSUl+RXrfUsh7yh7s4L0KHA9
YWT548kIhuz8HQIp66X9PYp5lAm+EtRGJubPUt/zfNc+7kC0yJcXMpI581Pb+QteG0y2MOsxOHwc
ggVCkeZzoQ8g7q/2CYU2mZd/WW+kMX0K/CuAWrO8w/cwBO4AW2doOmmzYNzsquxYGkDmRu4B8eU3
/inIoUip/6CCLpYl8Q15LT0UJxxZrzdYaT38qTdFvX74BDjvdbk2ogcLFy2WhUbWKNixgbCChr1P
veRs52SOngJDsAvqTSY+p8+yFoRR0qY4MdZTjS7HYZnclecZVlmlZtwFfoC12ze7hTc+LJV1cNJo
bHvbT8a9GC5umtxyMn3ZPnoCm8fPsRM0RDkEfmaF6xwLRdy8G41NvLshgsJGE7xNwFM7QUYpaTVA
fetEut7OCPL94gdOXMVUx9dCTcA3MHxidcDvvWzzuCwEDn+Cn960a/P0Z7e9+H7mqMZZufOPQ2e+
msjGZbF/rpnBCQIHf4dL3QKVZqPBGNvoWP0wIFgbqQ1rboGQT0VvRCanYdzBORyW7ua0T87LzkPa
FHQIFsw6tqrxxEWfMHIBnJFbNyQVBKLo4USA2qJn3/y+bZajRykm1ppVoAjl9HzZTL/aAWoJgeZK
nPYoqhYdz6NtI8XzLevoc94iPCR2wVNuuK9YexR7mRCQTPmLrBJq5rPit3gHUcnPb9nOxfOc/tBb
TALVuN98LMsNicxNsg32vRbLtLlxtJfOwOzFiB8dbjY+i8u+ZYbsgsLkETwEA7gSdSOd2G8oiG3j
et9Gp/Mmp63ovKOHXj5mrsz9quTB1hh/B8M0+syWwjGOYhVomTw4WYxTsChzhwniySSB9s+GKIZs
BOtJxUCYMO6EQZPEmRuD/oTGNkQH0lOe0t9xdsGHUC9cqhDtUMEe024VfrIgcFMOWutcXbsGe7kR
5TCIs24/91g3ADj5y0SoT3sJvnUSf8ipWbGzPWOAV1CGr9ShAQGW9Kx2fxEei5LS/IbCFykG3wAq
f3oRg7t7swUhNAyawVFOut+FuH72Q/vL5H/Bgr2KrA2sEsD2pc7pxnrUKXmbhxfS4YUJY4E71oLt
4xvMv8rN0Z4DiHOiZq/Kc+1iC+UztCln1JZHrFjInvtOub+lp1T6MDJlcUpuf5nUNcY3k92ukxr0
DeGjKyvJW3w+R6xcCy04QN+vQZPI8j3+H9k3jLW2QPFZTe7c2rpUx8pRvxeTqvi92RGd2oSOpHyw
9P+/TmsIxHO4YBs//0zwnA3M3VZ4UPgymdFy9q4F7JI28zE+MKCt7OPEit/A4oI/lsVw8Jtn5Dmz
jDR70g7LSXJWfrbS7LzJSKoeaFAsgkwk/khr0HXBOj/csiF6YPsRZnx4da1Jw6Wvk//MFLfpVEDv
a442Y4n110uS67cY8DcCYSrlVt1u2TsA5oulOOIlvt8Jsst0ZDSxd0LDv5Djup8hXYqyupxQkkI8
ILgw+vbxZEdz6wZht2/7nIeubcVBfzgT5VnWn5IXGuHZRMvVdtVesfTOh+KFA6Ix0rktw4osDWzN
oV8/GNwz95QxmvAbis/dcgDFEPiBBHc8GjM3FAFuOBmomJZu4ea9LnlILWHvGgNheI60o7yWLuoy
aq5tFSy/iVhd21ejHmKlzjv4e2zfPTRpsL4qWmzK1Qe4/iPhSPxei1u+NcEj/VL70cHp2aNALtzD
jIJVMnRsUaL2Bh6e0u0GBgZG+8pLb4WJaSQ70+q3ee24ZD+PQMafFUHpJZYe2OamK3xp9shii+OQ
C/vAjjRL71OEOV2v6inpbBrZzv2fw9uiMIzbkw28Bx7Q2gvN8OMgKhDgjxhTOuf5QWp2SXdJICxa
csrEwJkaXRuRySvampc9PBbt5ACP2vngUd163+/Wdv3/TBUS/1Pmx0acEL7DAx768iq5da/hm4Mp
qmrSrULAQYSiryW2C3VT/8aAP/QylYKs0zG0IybGrp9nYPd3ULVeQyqZM9usvVDGUPeI5k0il1TN
OKxJSSAJ6nakxvbZitUlo6o2NtDe5Qgb55q8Ha098aujemx0DmIN01+S4PDQZVtt0LhH5rMzVwj4
KVWEdnhjgfmUjGbLdRic0ayP7upCx8kK+erFPiddstDhMPp9svJjhbrVyVaFeZkVwI5GSquLsuyT
PshPvGWm417MMHwzqx25YadhQc1E5bxksUZaK31vY87RDILEqbp6zlsWApNeVu7JegCZLPqtQvwI
v8tQgWR7fmWyOfIo/7dy+qTepJGsnAaB+QnIvUeqtlWetIxgNk3llo3V3sI5x71k0HtdWAlJcQHE
efw0shyHBh8fUtJm307dZjyGy3tHz1zttcP1LqOMuqvFFA0dQNdRCP7GhjfXhGMtcwbggF9GUY5+
HqqLJOKpsbVWY6V//NOCDzUjyENAEV0TK2+zkmqVCSk9Q4mIZzi6fh+qtqLM4raptDKuVrjNglig
VNoldGK6TfNpTT6tiBDs3LZlcmhS5C7DlgTQ00GT5rK8B1UM0eJ/0PUb1mI8/lcWOKEo5E9tiKPX
twtgDxANum/X8KYOdz5QML+P4qxYTTLqMvObzLy6PyuptvMrvxTF2vzEAe22ox0FyWqhwl6ozeIk
vVTURYdppD3FgsuXjxAcfL853ZaK5sbtRgdrr/BzmVhqLthv6cnHOniFBdIrlCxfcV7F8S234/6D
Qs2vOCdvGIKOrqeXurToGenlw3hxPjwkX9dLZ1R2hTcxrnF5W0dUs2dITG84sRj2I2cln9ci/T0n
8VLaDhxFICyXEOdOkbpEKPz/U4RCAFalKCb9MNU4nMq3edDcRRxjXqLw381cSfqFdgsCKYau8STP
lhtSI/KPbEloF/1lrBIcbcSxfm1mQ1AezWhFCzXsolg4nk4O88DKIlCDou81nfBRdw7rKngySLI2
Y0lWa7+8PV+3cSPB+AJf2BiCoB5j8qqFGKgD1cANhnReze1AJLJVREWYOZABtMt7wbeYUHb58/HO
oWhgpP7mRjgwz+djrB2Ip9ykP07itA5Xnr8T66dEPXY5daF2s0M2rPS6T/RVg+RFvXodcpV966/k
d2FAoXAnOD6RQTdk/qeZDPQY6Gtq9tW8Dm0Ijd8EjpKWqRd0vvZv2anwPrA0G60eQDIrBFhEaGMK
pUO1w3FK2/x8oBbWAsYw0/n6AXyT/pQEBCWk+sSuo45aBQCnRbuD01xRpbOt3Q80FLpt8dZz0ft5
8MPHwnKPXPl6thAoNwRUMdkAcDAubohIfB1hbuVwC2AsxCm0vVsWqeHTwkAE2WnWqRlvth3UvnVV
qcJgZcIs4W5+yoLGTs4wWxts1z18IYWJcqu4g6H4UWR5DTHWpXP6hWqv49dx3wjzWzbN13VQ3bWU
ZUeNTXr+D9wUxjQYj1By5Bl0oVcymRcwNU53OsTzBPMviEKrqKBGZ21XeAb1pKnh6f/lCdg8nlKd
yOtG+SAjhUhUm08VZ3RyFzi7Q6yu2OyH8/TkxjSwtvt+CaPWWQRNj805JpdoVavQVMhrCmNLRogl
tulSpLbxWwmQtHVhVvMKihPvXnY4gNyqHRoahAVNezeZtDxWvzcEs+Da/16gXodE87F3/eqsVT+/
kYBcys1OStXrevZ+Op3pN4Na5lx/FwSWoffMUoi6x3oeQzWpi/UzgRGgItnpNRM30yAoqjsB0S+h
qDvw+JEKstqcAlOdQX4JPnXGp6kdTg1FGuLKFKQBwbwXVxJ5OWeTuY4x2WWCwbziY/14t8YF9wKF
gzD+vh+AqWwrpMYU14TLeJxZqZBpXnVkDegPNGqZFlT4nTo3m/2wScPwC9WB/8l8q2d5zTtBLo6m
5m1Hjef0hSL2EO203pkq03neCGufJtPJ890AHXX+uKqeFr7iaugjQkfePYURqbFNYS2Uq05dfSV8
RlWG7quLcijH+pLB5ym20wVMfS9Ytpvfg4vjbkon42eg+0179Q+MUTbkh7mKnKYifuaV1QWgR+9k
BnNrqQ5LoEsyqrPPnLX/aqCoH+pUVqT+dgnXw8ri0r04CJKvaL+EH0Zh/vNNCEjgGUrk4tY0qZtb
RYYMBJrCRp75WxpbKYgmKfjCpen7sFstLvpn0v+unQW1n+btnoqSyzUrRWpJT2AtvbRhQnQqUjGU
SHxVoFVuw30b1t6B/pFSaWtkUbkVWHtEq2x+Ecl/AobWWp3Ds+56NJJSNA43nLT1Fl6QjMNRABWR
UpWooGLXeyh/vglkeLIt7d/d9hJVdXPVNomfTovJwI6rWydGGn/D287ORhS9NdgEzjdNF3smsFeR
XcBKUPsdoZxAm98u6/vYQVu+JevEeFZsGCYXEvMvtIZTbQqFPFzTmTWI3uiuCt4mRB0BXhhNaMdL
rjiQC5R4tvBe41Z9Asm8jprdCMNJi/HxQLbIbUjFgotSDYZk96g4veTmTHUDkBtEVUHyIMSp05+t
Gowia2cjU/KowPVdxbPtYWBHtYZ9lle3YYHPxXmSRA+gU3cYWsu/I2/NaZ0JY95R0QAqwHxrvBRJ
SnCdU2CssZj+eShfg/oE01uC5/gOUmhUNXO84cSugmvY2pBgFgEEEexfT9TwdGUrv1uH8sWgBXOQ
UB+W6XOoKnnZYgmCsablcp7WXvSAT7Em2qjpwWrIEUWqd4Al49E4xuybmRxsSsaKdL/6uoKsb9FA
aP4jtHZkPoi2YzTmvgI3LXDuJmUjYKqAfj2S0JDAqghos0L3xzignckgiGlNSLRmWRl77APf66of
dGvMFrt8zoWSg5R0pH2dOpPFeb11MemAV7yqInZCn+WuM71PkUnEcnr3eBVPFAphHI7e3SSvLS7r
3Xnkeg6TjCjvD1WRSsu0K7BJOUJdyWseYx0KFP3G2zx6EVd7Ii3TJounMF5h43D68HC7YBmPbS0Q
Wt5iM/DJRAWO5kkOQUNfGLJ/REA27XylyNSrGXBWf8Xh889sON9TGxp53LpKjwfIRLgDrhnq70yw
Lx1EFTcwglJMId+NEwMpr8c2PWmsdTyIe8n0cmF1sCYEnxRZU05otPxt7uz6VE5w9LuMYUH9h4Jw
0sHN64SF99ErR+iFqctZhxJz22tomswG7k9O2fwjo6e5qhUoB623L1tqbRh+3+hn1ZO55vrQXaUm
OOn7RAVX5+j4Ht5TJI0q8DwFP8NEkDQQxgbmRNe6forM2PRdPiZe1kc22D/U/6ErRL3cxNKJyVB3
MLYE2GVdMsTd9v3b8nWYknY6zIA1fnmdSbq+VJffgHh34EqzlynKlADSaBvgq3CoiT9w8ZHaO0PN
rumd+OpjyCz/jL7bWr5mXk805lCw3rtLuGvytx10Ni7EF/kQVTmtitheI8xuKP8w+DoEmyzd3/KT
NxOLkaCpF8AFpjteBvj36Czqav4AH52mZR/ex6VH8Ki/Nxttt+th+bt4yB0q9jAGjDhN86WFNTFx
nFL3GGCh2bIkgZTdRfKaaUOdoTSIDnck53f8yJd7SD6Ts0mJnvMu0qzV1RODdXCfuM751obJu8tj
Fcs82MJezTVkBY9hqd1trUlZqvUzmprNRttSV5Fruh5rfWy8wBGRyX9yExCQHNLfwEwOgnlSiMlM
BoTQBK8zoVO51m1xxUiAXYVENwzmZMcbfETvCIswNQOIrr7GY7b8/XFeCWGDJSlje3wTcG/OgFdX
06JVqsyRPPfCgSHrxtxqxYqxGKORGlw/fEaNJu797bS6+bBcV0ro4lLHZR+8wo/ECnVjaSUT00wj
3UBecuIRJNYco/lt3ZAEwU7NFds731jYpMQvwCCui4XX4vsESznCeDY2Kx8p6GLNEq4YpN7nfX9U
YdLi3O9xNdVm4uph7nfQFmLng3kDylqoxUNJBYv9YBDPXL7opMWKoAb8tVLBHncyx40crkMlBxnA
hdajyjNbzG61DNz/9lpl51LrjgPHAVXPiBdSuXgG1nrmrpJYG1E10F2zBuJKskA1vvf1YflJr57U
1ify23eILDLJNaypyoCCnBkryXg4pJW8OcMrfTOa9v5varImRCQYgDYOYTARmH8bWwdUaHG6qPOH
qxOJ26hOAn6pPFMZZuLf79ap+6YWP8k86B0OEAvxFDVqsKsfWV1Uetg8WHPlAQyxQyK5U2W5LrIg
8NQAekL/Wz72GI1vYh90vF9Mg1aJ3IRWACvT9QCvqbCNn0o4lkDvHAZVwwv204t/XADiIf3nGqwW
/APiqdvoTpQffPSPpi0ZXOVo4L1KYbhZf8i+8t7T+yvfIqS1Jo5l9l3QEWBo6WkCOMvxaWrRsKJ2
GWa8utx4zf9mpj63VgIMiLKH3LV2dcpxC/pJS7kd3fc0tikBB4zxcbYP9PDO6fv9L8LT8YTTwwSp
05td82xxRmT3U8a3HLZ2zgCKMeTg3kttx1Eu2s6cLTk1NZMHm8uEhXO0+BgStq3S81olEwTeVLT9
XSJbSFUH7l40iGZA2Yd5u4ShD70qG/EyCJhwsanXbxIzmqOy9dtvSsDSTSgQOvCfqk3MybTSwsgL
XPzeZ0KE8adBPE4oBQ7MYya4W1BSO3d4aM6oFhFn5LzBr7B3JWUeTGOewTtzUk3tjQRdOynkLfUT
i9WHLFV2SRVJsRcqFunikNEWwb6s7tAJY3kjPZC83TI6oBVBEdMNix/TlEtlTcEkBgo8aI9XbhyU
DxcAWimZCjyJpv/Qx4O2MELnWlPUgCedq+VH7BG9OZcED2BvWOHCy/8+TK7XZPP2+9m/TS2FtISh
BsXyeEJBWZB7FXeYfZIumLT/bEUmVK2G2GZ8FrA5sZFVBC4rFMZFMjAN2XOOzNwMOTnWKCPgC4WK
zVjGD9NohS7cdUB1m/iyKdpk4qNmga4YF6acolH26TVVsZCHyX77/o2Av/gnU74JgEn6Y3WU8Qg1
saIfR3JQrhp789uzVliI94tN6f+HBnbLsZHCFM1LUnL4e4B9AI4LPfn1BCl3gwiMv5hoZQQAuztt
8iP/AZSmrxE7oqbKLp4SUY7zIAchCIMP9YOogdv3wXUPFgHUdGrSVBAydRXtmidbCa+yAvaJuqTZ
d5u1YmmJWtM57qoIJwfSc8g4AZdNrbD+euu4PQxTTfA1KxTSC35z3kVr/hVJ9Eeu/SInHTqXwnoI
KiEAENWPQAPwvwDXUDrzPwgXbjVwlOWqyt2w/iUw7kBxiKqpY4PCLiXV41EH2pbnIY1RjSJIVCgz
MEr0wx22/DiUIkvyK9LrumDE1V4mNnAkkkf+oKYCYlu+beq4yQmeqLjucdVgWdQEA21AJ6lmpn0b
5Cehl2gpkEx5iAY6vEuiTaRShYXLVaMTLVsRD0juRrS/FFNptVUanSJwUTSZkHcWQ6CsT25Z/X+i
3vhdGYYijvwXslaMrvvUvKTfH4Rz4X4+/8tEoJ+7YmpABbxX9llOqYdOZcsGEIc9buDSlujAZXfY
hgSCC6HSCO30XLCbADlhpAi4lgmyJz3WW3lw98syQ1EHzpfjDrqFRNRYNam6HQyXHBThnVlYyKx0
PPyNGTz4fL59at/tQ+O40X0mBHL7bhkpyIQy5UQxraWurf3do27ZpXXowKEr+i1FN4bTZNkyhr+Y
VoVf/2y6uB6Eq542H9ZZDhhIYogb5YpiY4tmnS1WC13WUbLsOUkAmsKunIgn0kRlMMgik1MAgryT
klpi2k86AMtQY2QY5NWVN87KdBHHq86A6+n/aAG8hYV5LvBnii0JqJlKwCFHa9I1yAQvgq55WgOm
gbSLn3RyG38FzRmjzoCLmho+Y4GFszZFH5ho4lTy8wiihuCHTC63byfp4zOMCZmGbJwDLyiy0YdC
6QaQ5GPt+3KPPPZMVJjg4f7RltHVS61SsKTpaX4jdPpotPlzeVa8aWVB/KZWvDk746lwdAHMpPG7
mW6JxyIngaKRpV174h6LNQa3YaMdY8n28KjIVNajE34pcurqL5A6v+xmrr8XfgJpdN2/YqyVp8Gz
LLFy2tcmmBhjHYYaRnIfE4A8TLguQlwAUdN0ntxuWpw4/XgVAY1JJgocw0vUnOyItkeetnrmKzEZ
S9jpdce705SuzmwBoF71aBn+Tu05iaUX1Wx40sKcfpbw4diYuUuS0X7G7J1v/Ib+JGQEb5j2AFUd
Kc62JgzQoVHwZ1RGsx+chtwA4OD/OlRlJGEJ5/Y6CQtqvjrvgBNqHUVlbhswJ2gRH3TAW9iZ/67z
JQ406UtOUdFhxhFbuhAH19edgmW2TUVEUz2Ivf4+nkw4zORipUxnvMLhqU4AT/mvJb6gYnBvErl/
9GNc68DqhX+beH36sTdk7lNwdPlLJ7asKGRu55AzI4xKKOUdxlN46rCySX9KlyZNWLaqgTKQLOmF
5OPkK6vjeLMgRXxg2wRHCgoVhe66lq5PHYs8sBds0h5XqNN6eXFUYDEiLuiQzy56o8pefwK3yhEe
FVj9Ly6mXp7HsD/1+hiEfrsFKshDqBlvhE0tCHkS9MCzDgQQDeuMjbQyF7PaR2WWvMqcK2FcIs1g
wUQikkEkxevJJtD6FqJ0hW9MMetyod12ntPUs1NLOiuaHyykoqVAiJdERXyfo1HJwNw3f2EbLbvB
QpzRdbhxKv1r36zctlqqNPJMOLGQDSkGXuFgTZg3zF+fQ6t3FY8p4xG1uQAWJEkeI5SCe49aib8I
JiQH5A/dQIsNrhYJQYgzmLQ31/Yiog1C5u93tqZfeWK7Pp0mu7hFi9Qtoo/ssldDIGtYz5arkQ+2
jmeBK6g7O5DlQg4gzg6xqWljwzxyodU5xebtfA0cW8pwtvYnVtKhU5efvyIJ4yeYrWeMbA1mP4/c
kC/T+BawaFxCtrs75g8hEaYN7yLGuy7dLiZ1q7U67jqAavo2PDjWP+uhgrqYDa7RVPKfyYlWVPiF
DuRZjD1bA6pJqXltQmXNlngVi7z45XEc1Tc5ZvT0nlepdJ2n5WFnHun8IolXCHpGZwu/Czydr3FI
h2eXo66vvfoCYdWrQzkHOrwlrmKdEgk1FPaO2Xv7inXBjMNsK2EY87fBPyA0OWCR7Sl6idvCSMgY
HXCz5QjSkHUC50v4sqZALtJvelRs6bqyKlGGBzARNvMA09TcpapYTQXX8iPWZL9iUz8exGdE7gfJ
qpk6P5eGBdmrV6o1WFYLqIxqhNpXx4Bmtjh6V4ldtxZFKz9qCzT7bIc27s8cfTJiM8euUIc5vgo2
5oCccwcRWuasglEo8buEvGeKnS/GRgzkvVj3GLw1PITAhup7Vm+IRfKo2VThSjUvUXLDNAitqN/U
q9vPY5BQ1WOtP4q0CHcLTEsI6cnTf+7JTjCsfui/cxL1XSEip58misdnjV+RvAyyPVaBpQF/Jd8Y
CElkIe7uj2xQGxIlY7ObieeNv/IJ7Zm1swpQxP+CjgGsHmm62bv2UhaBX7w+LPMS2r4XcwUIeHwj
pjWLjz0HtYD+ircfoaUSLXoi9lUkO4U3BgUW2dwohA37MFiD87CzfaIkvCF8cmnVtsUuqKr+sm22
BNAoxdPQqHitc0J2M+B56lyBhNmTWDTgT50P8W372g73FlSCECaAnE2N5Ep95Ek3naaGZx0JUWcd
9p7KJZgMIN+aqPbDO3zoHjGwyI5cmJYPI4q1csdlJQ0eqK5y7hKLhqN0RVLiV2IZSFup6WrZjgaG
IeuYp11VOCTPqMAExjk1QnZTBRn3FPumrrhGkre+YoDEPRNb5CE9xBez2Q3rNLd+OPoMadEjt/3w
xnsLf1h3/VxONonM0VvXwQlKwJ+WyVKkvWnNxYZ6YzIQbmoEHnLEKBy79zLUJ3h9uLU8sofondf1
jVprS8LBxSW+XBJaTCAVG8YK32fk9rts940h11aEes18m4v12GDpUISlFr8L5rmkbvrPNfGKm7Dw
VxHDfx2TY3kLPqKP6xttmu7aFuirfh/sVe8C0Fgcb4bJbzNwRusvyiQJrpzSU1w7IFdWh7yY+3yQ
u0elkC1qDPvUbfVqZyBGl+QOGqNaN7i5adC5CD8PTWCKJXCepvAB4z1GPVbrIFMiOdIQM7jRJxth
6L61BoPq7Pu1y6TUW6mJPc9+WxMtEvcjd3jgZHPlF5LRf9H8ZwGDP9ZDSMwth1W59JwSVkRxlWXE
A23oFMaoUHFhBZJ2ouHL+uCIH5qUCqSwcKiJsh1voQBpx65CxAciG0HF+klD64Qp/s749x5lbpGs
yus7W4FKJ7cUcpDztE0sB0I3JCKpQFFYEhBS0VIKC/Xf/aM8X0y2H0s77l3LmMEbQqvewgnMddJQ
M1FBkigsrKjp3PB7DoDL1BGf4tM6VJ5Jx26XR7cx7A1C7VufqTrN1FKh40FWgNWhwXstYHHEXwHb
GujKzl0CUY7H/xVGlFwVEoEF5qzYfLJHYfJQikEwfGSvn/1ItvM7gweowMgnVcldPtmqOUPp9/ky
Swn+OaxY4pYDvCWtCbabxk5utiOlXYyTlwWiblUO3zH2C4EDfA50e6OyGaYw2WlUHFF5yeFwxQt2
60H8DDfEnBHnqK75WzSPu2o5ojjuUaHQJOdwKTwAlHEBoFSDgPMGh5BB+b8Hx6GL75GimQmdsvnh
OIH24dddUcoMwXSIhVtqzEg8yBOQDE2oEPEKaq8qlJxBkuELuGOFmt4HOYuxH7BU+Eq0n0HHvNYJ
nQ6byQRQVprTYo1QW12A/XAAtQufKIoyqvvMQDv4OAS09jTBgXmnYBfBWv7jOUaDkPw1ZimHUA/5
mIUR0egB4ckzlXM+k+C/uY0SMEZxi+J5XHQsWQe+wGgJ5Qps0pSt8zEzwpP8n/9iowziZfIKRu/s
crXNQdu4JTgY8fFE65Ya1TeDXZ9Ta3LSRnDj/pyTEMUoiKTh8fHq/4iRQ5VTTbZ7Km0tq6izHcA+
IJZYrASOGHhOW6t34cDzhuCoZjmtr7lYJpH1XWKsOtxoReMEYS+6+pPZPIfa3uy7+pTnHanew8Tp
beVhy3wR+MwOm+KuKu6ATe7ngLDIZu2dsDsdVT5tDcn0DIiN742ky0V9pnPhkZjhdd14F2bwqTh9
vhPT71uRZrsRub8j5Vb5WOR6rkfA3pCpcpMPUk+JXOODfhvIr2oB2JCfgkoCMCIjlFf7Ddpekrp4
Qz2oYPXQt4glbFnVTmKswYJBjvOJnaL3HOagBzR9d2P+RMaqNRsMyZcUtCUreHT6eHd0G6mgZJt+
wlk9dwjIfV9d5t1fPCHyw/QNYhJqcod2MMF6WF6bw9uf1zmC4FeHTFsfvqDBkw158Za+kgXZL7WI
bClKyv+LOtZPTqu7JxbHNdbg55uhVeozu55M2ZH6/bBo7HqVeUqpxFl6IyPURtkZq13/LRPuCr1G
7Wgdx+72EKY17UeWZuZa3QiVUNLSpjRVOTHE/cSLWwyRq5Dq2VALDj30npll41LIYJViSYP4MOVf
MTJLIbyejIgji5H4hpu89yaGl0cTfJaExT3TwM0iZuEoSxEn92rUZUL53Sb+fKib1xyXZNFag/vb
jj5X6vampkr05ahH+paG92bnJfQi+P7o57GW+tgUeMBEcTlZN4xhK0cVMd4JVxgWYcbZ1ZbWCzZm
CrQ6PVzM8SFW2Wlw5KXbbuQfAutkrxnh+E5S8CALd9s/rGG9OmgMASUINOrpbDSYRaf3Hna5inCm
veeeXu6S6qo+N8UNEgvKLiZj9/b1k14A35dId20AFUucfoflO3zknjOM45nphGxStpoDgUS7kEAg
SZxyd0iuXWPPHUCMBXC21rsKTwlhnH4X0hAHhMp95jybiSwqbxnTM70x2AlYiRlf+/ZCYyPPs+DR
bnxxDmMcA5eVI5Yz17JzmaWNMYEFhEXNGFx+8rGuRw5mRMDBJICV2GK3TZp5AIBwlr+qA8hMZ/lF
k8XtsM4m6x0/2YYh/BWGbQg7ADB5sCwBHxE9IFPiXYtb4xKwIdNIWcUApIdI8th4T3hxWBTaoiqP
FQJcX5e7YF/2hZypUlwdySIaAiYLIAiIX4vVBz4b84UrbHRNzSNhLh4ZwxtKmhAdAZeAfOlT/GjR
D3q8QhNuMrJbl4yxUIvloxgVH98+1sXTgJIW7WHtUHEqiISWYuznYH1humEnsHakhkMMeZm7qfqe
m0855kO84cHZ1doDIQiuz82IlEuG9krotYisZvMuG8ii13/IAG+1bM6mHb83q7x4Mu7qp5Yqs2oc
xkcQkFk8LI5dSjTQ8qJvn9FQ5WF4JXS06ZizarFAXp7oC3QOADq0lrCVq1DZZHBzJGR86xiHe6Ya
tbncEe5UEwbWd/UtIZqe5LAd7UKCAZtIOMVK/stJXxcFuDRDk3YsT9uFAZHwGpi1pz2OK2sploHv
144BuanjVUObNI5GBeQGFW53ey/tqDb2y9b+GQPaKoywp2ZPH31ngXXjGd8W2dHCjQaJqjvBVijr
BDJbqcIZtNU43RRsa2p6ieWl6hBjKC8l6TGBSEoN5mEs7GFFu3WtF+OrQpqPPAA0ZRrQzp/KW8gi
gjnCZEKLSIvb9/27OHYVzqyvwf+681mPFKEuMd/3xigah3VFq0oEVe8MC4EAuOLfP5dqH2gtPorV
bg5S/JbiW7yN5yjXGlKruNRhsvHUcb1w6VM94q7orxJ6Wyv0YhYt+asguFyApFRdahfwe5C6+ZUE
mGUBoO0LkMDCgNi5lILLkvCkSHHCEf1PI2DmF9kQPZ5Bw1LbLdNCb9w/OjpBn1BVPSBSQfVxg7aL
u+hNXkN7TfrWoWGBN8aW6jczux9xk9N0NB/c34O+inVlLIyKy/IuinZWrt02uo0jGjw0dF/uHzG0
hiFo4g6Kf04UwWEZ+5v7dbgE8pL8XitRj8t07W+amfM3qNR042mlVboyZzii/JcDrTjopFZXwbeP
/l9SBacrIMMRHWYN9HCMVq8rj5CkiuLCnYCDgrGrnVWJm+ye/+/uNbbEcS+omgVfWWeEx9mU4yHJ
VB6bkR80AWvpqwf78ygvVc2bLMNH8QUulCO3uXHUIXbPNch0Pj2Mxw1yMCYXNTwwafaIjr+zAYQD
7WNs2iCOGBSwpUyKsOwjMvDB7mkkQHPwlmhujUDd/XXGYG4YO7zodf86p+jPoG9V7s6Oa3aFKIOb
H5RZi2Lzct9E4qrLX6cAfcelY+lT718ek906s/ex1jJB/6jAqOsmCD1bcmCCZdaw/XQulNfu631V
YAPIhZ/PwLJpJ8Q1fK8RlGTtCdQoI/Tn4GVR9JhZcs67apwMAPoXEpaF7UdL5ZM667CJE1KWQUYj
WwVph4JhmC9j2f7qVSePMDmcFUku3X43mEGe4ARwbEYnAYR6HPfQpITot+2k8bOnjIy87L2DKHXF
KYfsGC254PYWmHoXlXNJ2S3xfyxWIwPJEqxiAr/IWvXFQ5tmr8KNF+m0IZlUaQnH7Ke1sUvDjsiA
ikxcROKHZwlOdPaZtpk1l/JBndkYFvz8QGApePhA9MxkAMoBtuGe58sxu54b6AMA8jd1JJIjCeub
LCO2AapAwZzPEKqH6OwojIcpSaD2TdlCGL06eAC2yNH0VOxSWOuvQZbFvCrD6h+/WyQy5Jp5tHnP
fjyiaeiKqC6SQwQQk500L8ynH6Zx0hbXO2ZTYUGScklB3v2ZNbQccyND2ECsL/pXPXjbmSGQd2wn
O8YsJjTlAUCyHpb3oGhantAsTJLTd1yxQJ3lO1cLBowKVF7HcWmQbJmVEN5+SYyUTLZB8jaB7RUt
2XEE8K9PMYGcdT96PtCLtazf/VeSmr6c8URwMKgxN75kTpgxIGfL1u9DWsjMZ5ySs2Jpw8kLW9Qk
3kNdX0YdLuHmZWxW+DR0Mj5scOVUHZUICWukRFRZCeT3d9OzUaq8ADmB8ukYGYqK1LFxDHfgWlw8
3+587UnXT1AIwUZ/ArCdKXP9/j5M41hzTDuhjkE6alsvOQky37ee6ck2aREXBBZMsKRNp6D2SuQw
5yaUGk7D4JQxzcjSWyZa45KYMZF/RPIlpAK/ig6EwZCJeOzPNMT+LDk5cIM3hjLZ5V89iMcdRAto
JLkdrIrLCisShnqhuhpNz2X++25jTHXsZTLzRONsJKw3Vy6XuxcIrb4DtUVrxc3mDMR6jOCopHmF
x9BECZ9Gs59ZnURwaWlVEXmP1daPN+0VHv4jyj/6q8QjI20M1hkFRwmiY125GRvEMYbCbFwP/7az
ergxMDYobVxSjfOFgA9q8zHOji0OpaLHFN8sLhvtf9KHlSl1tNNH+rcb/SAv91XmaZ0N/sq0s3GS
2Rmfc8zkECCobW7c3i9h9tHi9Lzgk09c7xkAfNmTR/5R1MECEDHZUNJRc0egoTa15HKdiZy55PD0
GzuEJ7A1YOCODeSvGewOvePF/KhbYbGtFEaKRbic61SIU2mMgDdzRppqrLiSaE8EElk+69J8OJEc
p4IfJG6hR5iqeycPt097ylEXvQTbOHcisC7GUfpRThGADJufab8Cvw3Zf95FWRPdKr1Jj13fFuHP
ZbT17ddMagu86DJztVjGqs6LiN44gqkgevcLWw+q1NtQBW3kVXiPe+//MHj02yFgalyHFuD2Sn9L
53bt6DaFhH3R9XBguGBYgCySWMNS2Bv7U0WgOxFQYWzf6zxMX65hO6FB36a6+J+eSAUJaW8qWqsi
7fjVtwnmERwYER4A2+Jylt6dJ/CRtIAQAWe9ljJ37sbpk/DYXhTTc20EpcRuILBd+dl4tJzH6c/m
5xfr89d84LKcjO+haA3zGxyxe8fe09xWdR1edipKhF9/Vs9cdGrY+ANJ4qEKcYN1ihg2ci9bSpD4
2I02He2b68NXLH1V+g2q5nctlvgoRRYBYetyEjfJf7EI06f9XY8T6cpnsSK8ha0pLZLraxwexTqu
tyFT43fD0Ra8AUcBDufjMNv8T9pVuytlgUOKnG/T955IEau4G2rgUtzjwp58siSxWYfBiRrwdytU
HArztTpCphYAXHMWd8E23S3oW9bkRc7GTpKRyUSo3gOrcGK52UDCrw4puxP/TUSc41fccv6ItX/L
ONGm3qV8SW+ezwuSdrdyrW9M5l28/tYCwDMzJTmqAgZrBpF3+t7TUG+MZrOcc7bk4O5OO28FNv9u
MHczSGPhqF7sFQE+GBZcTRfBjvSma+/LqbC+FGeArFnuvZV51HjlHGHjrgxPMLenObjWxtCD0Jw9
vVlC6GYBZZbQKqAjGDQkewZMafCg2qsCX7dVCv5YrAPkNIfg4ACkUs5xwCgEF8F/Dju0lpOVgjiE
L04KTHSt0lhwMO55473u5L2SnkVhY3TF1y/KZN17rnubkWNdjNrcVk3hbgnLXqsU3YuvB59dqJFl
dSW+1paOnNEFrFgw+umqYpijiyZALNMkh/vh1spq1eYNDOy2+B0WtP3KSzd25DYnqWrwGDei2qt1
56gn4SrjAt2Otg47i6FO4TKSYCt2yoHpVOoG1Hb1TMx1YNfUnGwRQqNoWsh3n7Hnpw5GTq14khxg
1scWkpycy9Y0FDIZl1reyfJcMHA0zx1jx8gGAQaaYuL9ZqHILDa3Ogh41rkFT56YJ10tvPP7X/N+
3MdO9YpwmGQE1uQcpqeaMBgfsqRyNwb/eMBjOafBl7Ld8dXdWBgJnXD2/MBBQn0TS92BYkmcotX7
/RKcorg4X7JlUOF+bFilR8s4E+qHxzFU6rnLIvBVsJxQ3AckiXdvn7ZgOumiy1dNXk+dWvU1/2R9
H5wYPzYnEr+7UwWO44HblmR0zuz13/rxIaSwyMfS1fG4f+1e3FDrsL01hoMw3zsmc6hTQl8R1+Qk
N+7pDNImO9mL+K7EccQegPvRTYBb5EatirqV4+FmC47YpcDgYKOCrvy7Js5+auQMJfgPeRHhCC2M
zB9fCtS+4CODxpkuznW0QCSwrNviabGSSxAsIIVhn1aySxIn5VQAzUx+PpzJg5cZL+v0zbV2/SCk
7a95CRDSP/AzeywtoaVb412gDxirKXSllGiP//esdWkB4UbMX5GgFrYOJQ0Tnxv8xtlgpITRoHpl
6CvNXj5gJv6aD0ZgPnGCJl1MS6cxxmTKjUZHmD6GHtMA89aeI9WQaWwj88gtwO6sS9FwAAbo4Y4m
U1LNFiBdwsspqjSMU4YLXKN76/fJ+S2PUaryRN5XiO/ffYcdQhCHJHk4hyrRFoNKk3WMLi5m+hDK
qAkMnX60oUfR0sQkmvjCYVzIjIBkYakK03NSPPSwrL2P0EVgf6ER9iZ5zkp/oYmzfCFILfyZe52h
ys79Q7L3JWQT2fdP75w1xnnmr8yDb4fxhME03QORSCDNtSauGtknWOAZj4xZyR/kKpterT3wdWeX
4ajr7b2JL7D0Z6bLmj9HE7Veo2YRwZlRtcErcPHePK3QHm3I2iDOs+INsFRzpKcev3XTsQKvkTFj
5A2PLiKTk6CAFhjMW1Xmr7hvwiET/rHOA/WLoaXITZXjzrXmdEtORs0On7JyzeTxZ+gcRpYVx6v9
BaPP13wFVyubZ2LhVUPvPE1Bo05RUvI+ghk3kvq+w2W78uW86gdr2gUJ5fttSKotR4p1Xy7wrNcg
yqVwoui+aZGXFlkuKXB4o4XuUL3ydk0dWZo3yhhxwgLDUGBXHaTTOiowDg/nKvb5nyAicZLCp10M
TaHqHSRo6UGboiA9XtiOASZWDh8gWRdvnXCZohUNsSy1AeZpvvW4jlMq7BUGB8yvy7uFf6GHi0nC
Bpqek0HSDgyvmqzdztYx0lfdSJrRm1V+00LKRXNgJBETp15nWEgKmsh4Jt4v+mbcDM/hcI8L9F/0
Zinwu1hqGhxHDQkBUeDIk6Bmd+fgsk6hdxabq+GMXufPLBbvUZ3DV/3IJ/GlJcc0lnuPATCkIKod
uB3BGtTNIeuiY2WMCZgQ0Efp/SGuBC95RHx2ajRW/o3yAEAND+XUEr+HES/z+/XxtLgaq6IAs+qr
Ll/idLON+AjtdOF9qqrGa1CRcHwrEyJXf6c7QmxdmX04Lw+RmQ00/VK2qELh/wu6IB8uNpfkFbEI
510BnESvDZRh5Zw1HxOakoEjaWTAvmBZSpN3hk3HiUKiKREIOtSKmoZg0JiCo9joYihlXSoZ3jNB
wGhX4cdZcDLUEN4u1zeBeXXJEgiy3o1pLGkiwUI0+EWPeC4Q1eYJWOlYzh7/m/MMimsMgKSzRDaX
tfmMRcpUngxErtgywBbBnQAPq/zH+x7fEF+6lHidMtaC+atxFBeCk1BgSupi1mVKpXH2haD4gTRL
Xa5FpHnjOTJheMmtn0pqAT0A3+aYHZa+3Ku9WnYgFShWo0fKsP/ksF69WtNX8O539lBS/EJz7gB+
jefCfmRPwXJt6DlWNYJuXq4r0u++zcOLv+Fg2FjCdMgoyREB4TLxKaMsytWSR1MYT49YXUcFr++A
JEFk9l9sl7Eu3yUy5rrMPBOgTmmyPmv8jC7y+13FxFKJIcCqmh/jmd7YRaVN/gHx28EX6fi16Rxp
IHtPrqXCblwsST83h8k06utKWit33Uqkb8O6mc2Bwyg1xYZCKut8Dj7132CeI/usLKauU1DPgBbQ
Wd3BiWRbhMPkJG/8EQLmO7X6CEhdsRoQc1RCdoMSfweoCTf1pu0AfuvLgjEdClO6yJag04nBbLaq
Y2yiujT2TgtPHyFFntNeQszy7FNs5IvMvMzRvrj+16DiZSw5fJPK805oa1rA2/1WiRc3qQG23QVr
CSk5AgnfwT9bm0hmaGiQ9spr2ZUSR1a0E7RNBpJWLsQDrTpCQkYcYPUfjlgx0oHNzD+GoII7Du8J
l8nMjj34YVeOHZaKFrulu3mU3LnbWaj6fxIhZ4z8cXPFT1WFZTxQhf4Cg3VYW+gHMEWuTOfSt3CB
s6QaW6T1ll0+0c03s7nSsgoWmja0rxoM5f7cGwNm4M93YCq0DMQEeeKkOy4BHk5noxxWN1e3PVo/
nMRWWlIwpPXR/J0twhw6PO2tYTjkbcaZyv9y6zJQM6NNoVblHIv+2M8+VbUE+TGjAi4SbP+TZDs/
kP8oG1dj2+Hb22YN3IhalULRtQ7gtV/dtRPQVqWoG3j1cDHZvY8ayHLDgqmLzKr7zk3pLdXePk62
pM8Y4EdrGsvtcp5W4x/Jpe1++gM8T3Yyff4ulVIuuG/jU7L7PYW7PRaBKoWCeXn3esBFe8xJ/9IG
JbT6Qd+gwLvhHBllHBa7nqRS200/J4tg4tFO0iAlgYRa9Rikm7lyVwJLl+eL5qjOby6gQRnEHuFl
+ozbfBur9Fzt2fCmoA8QsLFVjErV7t+mVoD0JulPxylEAqb5DIav6yLg/8OdeUARzZVuGeQDNHMI
esyM+lJNx3IWFP8mSGV4ujKZkJAV3VxXR9No8saR0HmFS6U9sH3ONNKTVFFo/WGZWV8PvMzyMPNK
/UAfg1x2gT3JFSs+Y/6RWXdW8Vvi6I6oZCAcoGYypbcPYGl4Y7YzfyfwW+gQrigSRm+srM80JqSN
Zun4QVEpETuIdv0PP0vmYUVnhOII7C3E8ct4ujnptrZCjHMeS+s0jpVMi7+6TZLM3r6uM0GzDcEi
FflcoDwm1CEZC+p8drknbd1EXq7glo4Rvaxm+QWvx01Uh2dgKATSu44Q9L8kOaPK231Hp1cAq7Ae
8tZ7f2M8AqWKyEMFz8KgmN8j00h+Uf3DhZe+reFYrg/c85UQLN98OAH6j7Ko0pdW349lEr3ldeWm
6XEhlqKoY51omfjfOi3MQYwn9/thoAjpWdATy2JMssJa6MQR2H5Ul41O/9F79WYogeisGWF1w+hY
7PSMnxlfVDjxufHa9UuvRswBKx0y+LIUSkL+gU07CoyyGWMzVeDWIpPJIqOIaLSCQ5q4Pp2Vliz5
MM5p4JMWS5sAGmML3i+TiQKZacdo/7vtONjq+5njjVpUbkP8Vrr9aAR0seGO+PeYVmJHidQ2/mIZ
rbLPc9dPxw3U8WFbLU50hvZ2TdTOri7n6gMPNicIoY4mDOqOM0j0ILo4OqOANTayXJkgAkHr0K/m
77oTnPR2EujxIDRBV+fovzo1dgJLmvupR161ccc3M4B5++gRx/whemO0ThE22lMwigyhaLOMjriR
I2zP16OvaOTp2unDp0hDe/cQnSGP90uKwzQ78xu+wIm2W5YOTKwA7kz7631bCjgX913MAEsEQBVT
KeojLYjuwKAdSHFLDUw2ek6c4QDgBOJhI9P5W2cidpytpMBTmjvz7762t1N5+fvEVZEzjwcIB2bK
3qTqaxfxqoRDIX6EnDynpn96VwNoYxukC+DNVYEjn2nBoB4BOj2N25oILvf1N9yA45m8Y9X1SieG
NKkcDDFwihF8sAYciAJLtHi8sTx7KhtSt0fqE6802IW/Z0ffiFZ/l65pNVuPzgeKJe1S2IlskpAs
z9XaBCdZTzO+mABjIqKNATfgkOVuhLRcbsnG7OxYZEjFuorZ0ZeOF3EpFytp4zg75Ofo1l73DHYu
Xew92BYxHl7c/NOzDR5CLnl+FqrsdDlFKXK3At3ab9d6sGsnD5rv4DC0fKa9FUVyuI0GfL0T6SBv
rovdrcO3FO+bmy/gINiHssI/UJslJyfIRgYYUsRJukd4EHMkS5E0WtiFOBzKt9ZzZIGjRRvGcIFy
7ZU9debZgMgIlVF8kPpPz/4ex/NuyE1CgNIGsWptYGkFOu4lGfoj/ffj8UR2JQDrCXA4VILHNoAG
Tey6G6wIDhAoxt4GDTgtZ3bPNvcRXg0Bd7ovv4KD7DL1lLRZvW52I6X/0dbX+nLMeytUSYxnr/c/
3UfkNaBGJY7vpNLN+Ylxowg9O4nk6HK03YtclptIm80DulykrT6PPd/3C2sgPgmWVs8+LFCUJ6FV
6BT0V4c6vMI6fXS/0WYj2o8KKpJi47NukSrNZ2NWayYW7EGFMAJoY5+JmwfzDlNbA0zJYPinEOIl
Asf/Mpn1tk9lL+5EE1nH/P2sGvL0DXpHLUi11zAJPVSuzZG/XGeZJwIq29NyAbsEHsaxxspmJBis
5n+eSfwcM6P1aq9Ok3q9/emTctdjxdJukyrm/btBDVSSlDLJ9bxPAw6Btqg200gflrXvSRYzPr/d
nTJccB3/HmJGDFcDZgECyX78bNgGKyIajMGCBtqGsmcVb1YSCgNowbk42iLJlq7KWg0ZqAdrbP02
c0UERnff6mEhJbCKXMsun0qIbQL5nLP62/j05AJGQ2ivmi96pkrSzNsZ8x800RFX4069ga3x7249
+/jXBVTZNQwkacRm6PXEtLQ0ft9XPNekeoISLu+5PyYtF7UDqVN9ZaNnOs9I3c+bzi88ggMRxPGB
/XLi1AAeIdmKQTbo5ovbzbqn/o2B2v9mbdZPEGqBcWT5NM9OZioNTn40YFEUqe5opTGzMCSGqELo
nADaoGrNz9WdZJAerDRcPahuXKFqNLXyDlW/UV6pnHYhst6SzVzAxNyhRa0s2lpOdKTgidctSdiu
qNCv949uGTPzMjpQi+aKcDu6YFY59HtGNBb0t+PX/Dtr5Rok/+Sf/CNvPgy8N5MsqVLgkGORLnXA
c2rqd7msyPfwzLWhMbePYlTsW1sBaR4Ruh9DkjAJMwVlvNF2oLah1BUvxR/WqYhNMJDgRAhO3bbA
O7AVHk1AL5xNK9V3MkDzXoc1SQf0XsKWkwa7Sa1w/ou+9jjO0ddlFoW9DubkI/zLt8u9VY/OMFqW
ozn8u4Vn/jfD8X9U2UyvW7VXx+YAsB+/Whczdc4lHVIHQtpmPpU8D7/KGrqLi3xdYKu1pJ3GnQYE
GYl3iN+TlOPBPg4w7yxJtA1u4eKEzVv11l6j5w8oEFqUzDqb5keLyopWb+c2WDeSe/750ojCef5I
kDbz8H0BSJZUYaI6dCx/szYesYCEM3nos4MlhOGlgWXXYWMB3STRRCvduNFXY5YkFqFzh5WSBniB
POzTus9yMiS0J9xyFZBDAF3bJLBthh+b04/ULCfNy7Exr3Z676LMsVunFvO5LvNvsYWw3L9PBCHB
BRa2Ev3AYLjzUxO6mF0XtxHo7/gUX/EyGoP+QzWeM8xEfUWJYO5K5rDkq6m2nnmPs/uTTQBJuLBR
wsYkEQYk1qopay3rwyJO7jJdi8cvauDzOtVgg9xHUQrQGnQLvmQ/KZsFv5bzSkIW3xPUR3O7PE4W
McY9hb/NS+8ixb/63yHmw0STFwnlHKzGZF0K52CrOP4Ut/iJ+nFtmKU4P1xdk1QxLjxwbQQ43v7k
W8cvY0H723e43GQ6xv9zaGJcjhLDcw3I6TRl2VSj1P4QllzVWPrjzSavA4PRQ69HlrmO63npxQt8
q5VTqXI8c5a5bQqY1MfOqAYfvthmarAK6HBPS12ClsBW5LT26CteohR6T9ZgWuZCSnmbd1GroWnL
BzOpsO2YzXa+Y/add9yCrU+CHQz1F+V1ghhfh47rpI1G8UTcANvP6j/Un2VsI+unYBahEP7lCPNa
qgT9cBjYNR8raEmoaXHUCq5rYD6REcmOFmwO8ldraZM05LtYLcGk/JSc/HpI21Vb22Zj8eTNM6ED
QV8yDNfEvkaLDvSpte/eMUCWHik4ot4ACbSOR/rZt3ycBPUFkQfdUe1TGxLt8JyM/03UFS0eolmc
xz3SAqF3KV6SQOAmVnq9hfHV7eZ+YVk1Q9AGpHB4LwpPsS0GIzHrRgqwRSegRG2H5dfP2txciPxM
6N6gExws3cjlB0TOOo0fndS9EBRbwWYgr5g/I3W0XRxGDlRYGftk1ChZOtcX8nnkYU03luGWJZ5q
vD+q7IL7kJ1lgk5yZ7Rng58f9mxdAYUAeHx8690sK9Kj2zoJcNrtJlPLH1Wd3cuI3pdDsUyiJxYe
41BNRzN1rUJblUj3qvwbIDlvjfwEmN59kxS3ncrgZg1zBecPIcRnKW1nRxp0NYb+6HnC5Jei8taz
vPG4K1Tnp8VN5PDGn6JcCuZUYYXzxpELELEPLbqNK4QTQ4Zm7rMxW1ZX+qWOP9Q+V6z/EzTbEKPy
DGc+EsIxOakF+o1YZ9PvdfzeQ1wq51p/crl2FyzqTz+blhmULo8V1ICHhtKF7rd2Q6XyinepEGfV
20QVvOC8zqE+2OovSTektjfbvqBq51CWsa5WtsGgiRl5r4WYgpTYm1A44YUJP1FEp5RcILxR8BC7
S5OjwM/Ljro7VcXa1YsPBNPgQ47iVqasWx2wYClI/ZXSk8cAkOroc+disdWjmV8T6hkdgCfBJDOy
+2gFjdEfrReDjFnoVMJr08nF9SMWrsgWKC2bLBQUWGPkX019F9NtsBXH155/99qTtDY+RL5wC7mK
vTKQoyi2jPbiP5JVdT+0vW81XZtKXhJPJNU4/J7WbR7ay6N7tOfiaHl5lRTx5anVWkE2dHPuFRcK
pzFWFbDVbwoNYpQVrmU8TW7qrui+b1H0oIJ13EHCjQvu2Cr0UJfs0G3xeVtF3LbKJy5Yh9HHTjCs
nrZSqcTZj3WqGZAehxqQMNCPiaC6m+kr22dG3RzjzWnGTwXcxmbbJJUI9nWCTk8vlczgqjC0F30F
3naL4CjfMXhFwhTdUZHKjlLZq6oNeaXi0zIFjo963nh9Y1HUryUaGTpplI7uLrz2IDFuaDGXhHzC
LcviE25JpI8gGsfgXQEcJp1EY/J3mh2SDyhmTRimGTP87NiTWghlZfUOiAG2n6pcESOr+HzrmBOd
VbZ56KShlU0yndD5fvp4trWcdaDIAtAMRwFdj/EkBjeW6QTXnJ95Te5RM5JnyP06tLsA/m8rC38K
ibIN+ltHZDhE7ijHuhpS97Yr57+XvgeKlB5bYsyF5nka5sgpGfincDEU5A5DnOAIxDKKefeKhLHJ
WOCMtNE4BaKE7ari30kI+FZDHCChiUK4KutDrM2VoMHMrntdkhSPn8S+6OXezWcZ5D5TThoROirc
w1cGOLMHmGZehjExJ+379AVncoR/sC1en7BhAoYmyc8tie6Ivt4BeW70sChZDd1XT1Zo6aWGnqvL
VwZMSpntRQ0XYKROwLyPuno+YReWqZra8Swiy0mfhIBRpD35z3a17/G8FEAYG04vrWUvZswymGNW
JIuKUD05RzOL299xSFljf/Xk/TPaIJkd2x/pygm5DhMpgCK8iE1dUN8tHsEBpCkNjI6T2wo9mqnd
6pfJzJ63FwSgNj6ie/BFx5ujS4lh/K7vye2o96VnGyiFvOodxy/oZi9y7oRLdv6oQCi1Msxvw1Qb
bRgbQy7vHGZi8wbnExQ0WeMjXKjCzemUeKAavu1U0vQv1pNasm2KE7tfeFFLDm9YvZsnfbLuzwsy
52ahJ9O5OstRrJT/fZTizTIVojwY91tBbqdSZ/naqeSU94s1JEeo8e+pCSalxb3POmXKJj/c6m+W
y/BqePh2ToGGTR07ZinVCNR35dmVhflN+r6OnEtNj4leDeVdat+UgMIYPVxF3NHE/bwCKbnA+JuH
qxS24r5iltdwgpOX/rsPbVGNkhOrY2bccGcwGLFPAk8A9NQZfAPKRgiQ7rOkFFLC71jherWMuDDF
oYI+uM7L6KpN9vJYe5wzAUEwy0ccoKvLx9cbx7BqF+Ip4l4cxLaOYSucziW+T4jq2QakPqlwRMqQ
FkRMFSGdaWCxKCUqtzTj/v98izAYj7Ip75wLGBY53JXoCk3tVcgCNw0LLZzQyzvYvTx+Gy+MFtd2
4VYuCYHLskpA40zjPAQzUvjws5+38XHzagBaigFVTo+n1ALE6AHv4HsI+TYSG2kFxjfcwqTCSwSS
k8LwJidU4fEPuF7OR2pNPn9MfxlG61zmlmGorUhUIQtXPpUbsGck5TSj+JTIiFByuzN5COoCbYxD
9OU2UnzJCxRnIOdtBTmQLK9XkM1e6A7EivTwL6pk477tSOFAzmGkJO4rvo6aKO9PNqNBSlX4Y4Ef
1fv2eocZWZDmFqOaD/3izTO1tp4R0+GUnCm9D3qdoocIExcXxD2884ZrFUl6Pjew4rc7f8Xayhzz
CuOW3aIOtlSYiXnce/lY4FYeoqAHyXwV2oKCeOH2116S5b6k/MKOgF7N6pWFfo0RwzjvQVNlFd/n
p1WsZstR685ViOte3kyPoBhpb75oI7hu3Us3YGBK4Im3+Zw9kzmN67eX5G/khscp9/zWrwGeSCLP
yR6jQ+P3fuNVTD9kufm6TPyv2+HIr9PaU07Ox+pZpwL31OzeMbWWchy3swSVOiiNz6K67jzOFpXf
w0El6yP+afvYG1m4NBxR6jlYuwsu4Akqkoor03uuhN0HbcHjBc3LwsswMgeq4G4t+nEw3z9GfcCQ
bBvQ289LUeHKX8wvVTyExNE8mYNQgIpUiFoRmRIbL8/rjfAgwCalTbCFvF7/qjx+4DLqcjtTVO6D
J73MSaaYyTY752ZXGm6tumTn2dut4WUSg8D9J5B63lxMiHoTpwioIlXMrAZ64A5m55jP9Z4pbeyg
qI4aELTKpq0lnWgBfsAZCrThp3bA15fH7oUGTjohpovd3EkNtSKT/xmBBxTu3RXANArs6yyFECbK
VbXIpVmsoIQqq2MpG0DSQWRph6i+UPxGX5ls+1wOzeTS9N4MP9vZdURiP6dV9CbIDOEhutZudsPG
OSB4MjVzlBFifepWRSyOaBg50Lc1qH2XovDuLhBk1qcwR67xm5c2Ma61yyVHBS6jWkTPIf9XD1yY
gP8zUvqxEHSR7ut+KjLXg72FNHajAYKWp2GPO1PdKXnqVskf6XTDsIEhyv6ivXHOgPEXo5czAVhc
qn9U0PwbtewLXbnBSwgNH7VJ0f/8Qr0ri/JIo8Tcl6JM4NkscLyA6ynIZeXM163AzX4yuGh2AVbJ
9Lo1PSHGW+lCIl5fMFgaraNeTKzs2cIZS+pH69hj5v8YHfeKnop1ysiO1y2lpcD/l2/SKW0JQDw3
VOlfkh5GL0yhOTRxrsEzZVZ6TJTWwgdMzjXSOFHopUACn8YaBOnwkcoAYF96ZxtNSnEraFb2+Djs
NDvES+iM/b1jetMc+Gc9HdMsiC7vPPUDf1KgyEIJCM9llcHihwkhg1iZSxibQl/OxcyiSkGRpvgE
xJdC/9wLfVXZdGvHueUoasy42B2RkcqpUssCE+KufZVhwx2FS30VTeCSRkb/eWai4Wn40f/kqTMq
ZWhwVGHK2Md4UPhCYC1/hyIFOJu1bxC/ObW5STt2B95tRGACjVSmQDsMvXgUutISbXb3e3hrbf9d
L3fZ/SBXQudWIqh5ydQiLARe0N4qeKWnhq9g4vXjkUY8ggiLhvTPlBAhy9Gjbk86VsHFZQ8h53x8
4GpQsC8TrLP1k7DcrFhz36SGNgPZFViBUjAHo0/dhWl5mFoElO26AlVbzWssRIXEaZB5MiwaiqDT
nRYOwag7erwr4q0DVXh4vjXmZ7yVlwFCVuHHB6sbuaQplzC+SVRbwcINCRhH8lKiaWHDq7bW543P
U/k3P1KTvMIaA3gRZlX5d/TZROvVSPLfeE+losUk64GXRYI8pLqWAomww7RGQD1/Jm4JQYa+DytS
W8nB9n8pg/ldyVyXXZvKQPzazKfl7JtAgWab2tgHoz5qn/QTnq2dJcEIxjIxtTuKkE0mYI6F9/iB
Ohju6qHrmUo0knwK5TUOW265NFWG0IQXKoSOCcTL/e1s83ak8DCNcIv/3ctX1PUDxvzHRJbwYNb+
08yjcCs+pBtcSGP6vFc8kUQUJf+CC7OuY7VHyG5SYYD9beIWJIG34hOuVsK3X7QjaeLSHlY36LM0
/3bP+1vSrNt7vYCKHWLLD3oH+KDRB7LTJgBMGQvuk2ZznAkIQbai05UjAORhIJQ3jz6Fwbm+rT0p
2ka9wFzLjIVVgZd/B+TYaXxo1i0Ryvdf9TX698RF4Ipyz4Av9q+q2DFfHEQP0BsWj1j321aYHM0a
6Kipm0Xjg8X3I1pIA8OeXvyK54Y5SNYi7wzZ5S/9qRQykmPgNguJpPA+1w52ZdW0F388u2K/vAzk
prR0UFhxGs54n58dMF2deF4E0ofmWacVh5I2Mx/Dk9se92hA/oT5+DiLVlxaO8wlkcx8oVWtP67l
mMG6QcqrKv7J/ofCUl1716gS0tt1zgtStYfpXkNA4zb18xUQTOk5Hh3LDkN4Krw/sPCRNg0M9KnF
hHViucEOJzc+FwnDG0hR0gOnP6WCEDS3Bvlh/GBdmAOTB24KJDDyJIttIfNk1tEvX4CJB2AwVYmi
tr2A+VOmoRauxmy+cJLrkgiH0CoHWsU52vzANAgq7h3lRJnpl+fUQ7XfVKJCWOSxFR08/cvQwkBf
3xwqqOxK32tIjUL00/voOWONce5d+1SoBX9dQhjnuYXKJBu8tS1BHsudXqBPX45nsssrtxxjRyzC
1++0mePsXu0HTQahxhNWixGv4nAdioz+7AbcKB3ISkqGmPoZHKql3aGIXa2m40G3mLg7fXLWViUG
c6zYpiX7yQMviB3q9IobwROeS5ZknGVy+Kk/Rl2MxFKSFeN2A0VlJDfo48RPwoa+JTckso1Hy5uT
b8AaZwB4gFWSBWtCiiLvB94DaLgkEFLC9fzNSOwmub18Lw6sjCf1B9Z9HnXiUiVJ84JMEOyMZppn
5EmSJTVGB12uX5cRsswm6pPY2ViRJiob/0wCuGdzxcXBc5XWI+iYC+lQ5LrJOp+uDjoaaZftaGJJ
sPm97eFi7uToki1Qv3U+oc/mO6VptRleGR3kiFLuIP+IIgvMGubqDvLyDbXXW4pmpY25fwbH/F4a
aStANjjeeqGaine1zdA2iL0YVoTwLuv4rFp33hZRwiiamSfw+Qg51OvLoLWyJ5J/m7Z7oxHJJS4u
+2cE9nv8lB7n1/78yAsu0guniiRB/EhlorHLrm0p/afydYCVTAYuiecUlMY3Mp7m2q0aasK3rE/1
ZuUEAFujiOywYel2Q6vaoUTzjlRbKIvDmhw3FNeA2Sx+Q8T4juGkryZA7lTFG0/TIg7OJKXJvamh
nZdhR6Q/TrnbQR+A5JWe3XXM+nE+gCn4DKxzknCGc0uxN3SNyETs9w1jPobT3V5QVNxcjBPq/mSG
BDfWhvzu4BdSKYJgm0pp+IVEG8XxrTL2giLRqpB84nRxRGdJepYKIyC7J35WTPjevrHrLaxB6r3c
PO8izesVod2E3zHaLiIiDAYseElYRiGhTfdwJC4iYu3rJ0QNGbwhfr7W8cDZxqqMPS3no/vapFGu
6m+peiT1EJJqU/IdhpHQDzxF2YYD5jtsNaeECrI1/A3MagmmkYJl25eNRc0NKpH+MsEelo/cIZgv
m/J/uZSSi4yUvf0EJvgfK1PoN2/EDyMya9BFh3dJTwykdcAcnT31SiM3fXyfo8NaWHx2jeC7+KB5
fXXeJ3OZKw6L1rVyB8mUXPM5GNapO0dv++0taqYM9bcxNEa096+76jRHdbwBYxg0opGKbvlGhFOL
3bpa0kpHkpqmhBxatHFu3qe+3om7bK7JAuRZ0g6taoqyLpuK6VP44HRgTdQj3ahZ8by6or6X6cOB
MwvdB1/p9eUs/ir2DFufg1sMvqFAKQWsFHxEbgFxX05yNEz7UpBwieGQHsM0g8UvufGnWDwbWLvy
AvLWJNKSyDISV510zLIFZvmo9tXdY0z58TNASDjdR4g0Mvxr/a8HT+ifh8kSR8+n+anFRanKEX74
YV0GqaHoSKOP45x+LO9bSq1QMpriEPxMm3zZ8Zd0jBKSq/4vH51oyGO6K4zMI9ZeKS16W5nwGk40
cNiuPBHNGn7RG1MD8/Vt1uKhSr4+qV+xPBJTikfbl5HIw1kPmgUF/HH9P8JB3hiP5/bwiQK0mCMH
9f9sll9d0Y5sfy2XqUO4F5Fr/ndjwleI2/PcGRYv2gRjf/x/XZcaBTzu2BWxudiaXdVtkmDwH2+c
aUn9DYHcqOFDTcKucWuqiOMaLCinVQSConC5NGyOd1aehVF/zMS8VFYxTQWqXv2IknNNDUumIpaJ
01m9M47llIdosfvB8FaqA55XI/Zs2Lh4clSmaIEqfNp1PoHCjfsSbKM/6RKds9n3cfKywHsVR85y
lxMp5vBeoaS6wn0FNqPQ6YR2mGxkMjimJVxAhBksOQNC29/DhEhOMpvz56/Ux5yl30msks1tJLYE
bAdc7HQJu4Be2l9WujCuFTpVeVtVJlGL8yj1dtTHAhlWqSnYJnN6mSpGCPeobIRbO/nklZoTpL1U
+j9nci4MGG7Rr2P9qJwKjwnJtQ5SpduosuIyJ7IYvpPuhLOibOYccNEZ7WKBROKsPDgqSTBD7Pgw
0rpsqfN0gU+9QTYT19MBZmJlogtff9XLA7Xv84QJPyKDgu+XcOv6Ec9Ax3IE4OHN1vfSN0LTLd3D
34RapZeM7nUxfxRV3P18eiJBDz7ICX+FR5Vz/sgis75xvoPN5Sgo5TjiwkvCJx36mwKEEgMzmMCQ
SOaWoq5rC2ShUqp3YGyxnO5xXIQoW4Bmdg1em7v3br02oODmVDGFuw8Z0n7UWOot2uf/P5ihJBAr
WWmFAJOGmW8RY7dvKJyn9GZQaCSSnioD4/Wnyy1ZWYy1uEnY1/rqAiza5fGbhdEpCCJfWcDFvlWK
S0QQyhW9M56UXsF+2O7R0VaDRHGkO0DkAeQakmq1GdbKbrrZcpadAkMPUJNsWH6sFysF327xdd7O
5BpFgZ69arfeDa7E41hZSD9fj9bgoy2aR25TMWubIbwJieTzaeFFBHlf4iOK7VPMfVgGRIx/i8gP
020BCqjZaufL8GvhwTCBa1sBi1scXQL+ve9hhhp864UCACWeStr7pXJnfJaM2eixCfzcewt5rlnu
EBkgouiJGjTbJ3WP3QUixMPZ1PEgmewFrlpZ/BWfthNZc39M31MoH/hFsMEx8s8XopZR1rHtx8yC
MMYFQG8Oq1dDjmYsu/nNS9salmOVE2gp5EXiUwjHaWWm5DV8ip6q6so7uIU9xhc8uzp0OcDqnQDB
nPIzw70lXsTuZ9nJuii23NfOgzfYdD+1hlKTl4nevQqTF68Rx0QViFCbnq9hseUw6zzBP/FL99jp
kwquouPuAUacF5gxq2+ABq5DnhpJvZLRbCWFJc0clRitP/nXroCsjzmK8Il/7HMUsmH3hPwjQoJq
LtqZl8lBawUzRMxou/ARKM8ZsLYtAZv/WNGCzl6eT8E6NsLf77YzJXsyz/7aYZwrDLkBA2c6+7ST
ZjZGEXqNEVGZt83EHmFPPLS+bOR7npv9r6+DCXaHg6gYEGeOEPtpJV3wxQi5T0vsR0E1AhFIQyJE
0cAZ+wm/GAl4BQTsyoea7+Q0UZ126/DhW1rgPGS38CTRbqOmYsLrRp2PPZFVPDKjaacAOA6vy6xF
FKRth8wZ/UiDmmZhUVo1Sk4TaZoR7IHmX9qk5UKnCKJuUavuRxNmhAkQPloZ/mampX5NtzSs/bwL
pm0yBNLlJof6ttGxOmTZXY4Srx8fDiVAR9h9eRle7URdjG3F5xH/cODvXkrvW5tQ8nzrkni3dWnq
hePCqPx+6l92+OVRyVr7o4NG4j2EyYz9t3DpgsDvRoCesAHebZo72HGg+2njUqXTxlM9M3WHQ77K
yFLt1kXPXsrA2Oo4AfwRqNHlN4dLwX/QVxO4wUTgwkO52Y4/ZzpfYATaMYsHJVw+DXRr30FL/WM0
DRkF88OppnoaHuy59KvVAO7KUr0hrIOaSLlHfpJAE9eJYq7KpWXn28Ggid1gitHcAoynDvIqR3Lp
uo/Pq2CUUcaB+TMmUTSFQoYXg06t3DIf07Kwf7juUjC63UucNF1maXvcoRNfD9b0L/ohiQAjEaZq
KVempszfMttx7L+ij2v+Huqdtk6c0GOxNIGpsuOo38Qw1a6VEphvQl04r/MxsfnYtyO+uwIwfhuN
N9fk1sPjJnPT05kZQ1YgGs+o8K+EBQ8GnsWY2n4npe6U3qYb+IKGMD9fE6QVmTWCZco9ZM1krPFy
spMEB8gbP7nEuYuqkF5EsXDnUUxlmehlTQ+mNM/iSLgR/J/Vv5s5LqHeguLGmB3J1vAvjJXQAkcD
Uu5mrqxmgWiUNEGMfvuwtDUPhuSLSqetoeo/jkDVyO4albLBpxa541mqzUvRCYEVtxRzNPeHH+5A
ok9w51paw8UG31Nk1N4d6e89+tkBuoVmnBvG67zOQB8YMhjfvMlM5mhh9QQceQy9W+SS8YB5+VVj
MC2CA5ajUaVXrVzhS6PKazVrxPcvr7ejydXkiw1GW2m8qJeWt4SMVS1uzG8cW0JS0raljoqbkQPn
hdXyXS7v0m9Y7fCVglKDHD28GIg8uRXofPCCDeczGRZ4MeOnKWW2HbEd0RnKH91SWCg34y58Q7IW
hxUSWvClljPGc7KqR6P//dg+qH6IGNQhrC5pr9OkWbkpddILpK7Jli34KSGJxdmUO2zURDkt9d7R
9nbolJjVVM/osOqDtfMX4YE1oFDvluSkIMgLJFkphYjBn6uymaemMPi4kfENd6oaro8Q6mlEgXx8
U1I8G6okcdupBjyowAdHBiSkrrEtjoLSfmLV8EVBWXP/DSw6zbUgqxya5kPup+pkGKFYf4zaHhIO
wZRcmL0AxKc9ry0caFOYL1AUgfZLIx00Qa8/AYFq52KhW52HSKAhXo3Si3rLYViFdpQ2wgxa6FL8
8MCApJ4nw9FrdxfvAlHdtkpX2KMIsXEIgj0KwC/lv1eotpDuIa9PMFn318Rt45C7x2/QqFYSgN/Z
eUHQ+IblCXA/7VsJ0HyAmh/Cph5iqFUl4utVlJ/NEA6bc9xLI1x96TDbJI0NyZtDUrDjcMTSGOJh
nd/S+hLWwgpzuKsmzFdqm5PNf/fcqC1KZPIbTAPdf3MHS41en1MQRj9wirAMjCkypapHHY8SFSZT
crpIDh2qq6MmD0YyFb2RSImsYqTlVbBC+6w/1paYwXJJRj2thQFXJs9X7qLinXjVkMb2eOW7TKst
7GQQxNLp7NVDhiGWam2SJpf+PoWpiAk+7UzEnr//G4TUjuBWjUbP6jlzmzTRSF8abzmIYzHKuR3i
8kP5Bl87lhOH9voRaKcOTXMQZgCPIQsNO8RsGbciVhLd+9X5ks/kSQh5LaAosnJEagAs30gQVkyJ
WtgjZhcaA/rPekelTHmlOZUreE+QFw1F8AGmmN6gUwe+/S0Csxx/i2LC88VBJfUj7VX6ROqCPrMT
ix6nUstIjkcTv5WJGp9I0Xl1z+Rcv/qYEG4r5/zqpAcfmSdzwTzlepsFIrHy+G/AWUtklx7rTjs+
7Ij/+p3nZiWw+HwfdjxzQp0xl3xfW/3js7jN/Nfaz3qgHkrJdB+eRjub9yqh6wjUvCnqAQJgoD2v
Qs+UqTaauomsXwbBZBPW/+v5set3J1OscxnrhCsi83170mtlvC8MG0z0dCPLitpsf3oRJwolHx3U
iarsCP3qEsYr5vZ5YRYik48/S6k0mVnPsX7BAKIrMxt/H5QA7tUcAYDvZ5fYrR01dYE1hBJUEZ08
UwHXUcK2eEt9WmqKmn6QHQDAaCGk8lHsYl8d/mU+RJjjozaf+JMsMrNDUj6WUf/mKL7HcjmfHuIq
Jll/GEAqnRUYL7netO0pe3xd9ivj7KI8jakU+vadU5BdgSGGLX4e8vSIFTePEvKojh94NY+3vtcu
6Fz5wwhVlB2peFFI5EoP1yjmzfmqDm4jD5kfuh9RyaWyVQj5d8yOMrf8e+dVPONqAOKDmT2VpQYE
XlyeRxJ9XgALpf0H0WNBbc9LLlsmpbgGZ4kqF2PTCCwmf/lAFmJwP5YCMbZ7I5BXkllNUqVqu1PQ
xsenUgykNH8vIeKqiD2Buii4LFSnnyzLKDngmoSwXCjkUcqqdgvJkXLvoSGqAdxfckYs6+uD1OIz
aUzKOg/Ri09vdm5Cbw2NS9XBca0x9IRZ25yV+nFGzGpR6Rrjj+1gaBym9Gb5Nh95scvhLhPe5NvV
pgo9hI38szNC8y4kNVtRQXwlv0L6o2ZvYepr4Xyoacdo0s9kO4KosjpfgzG7/Q0MZNl11HrzaZNO
czqYbdOvM3gfQbDOO9BoOfp63ErROF7mSHgMHAprdc/kZhQwCwmxvmlmE/HmsjoBQJzHRMe81ZUD
jaAcQjJ1FI5ILD38l+S+No3nDmd3LgkM/wV0/vmSjZhk47nDDMDa9okX1pkFPUit9p4cjSh/deE3
Ox/t8Z5pqJCIw1EQLGY+cJ/OrIGfNR1O1Z4DFa9Gw0/dTiluIeqZ+/IL4skHuZM26T66rWQKZtNU
Xlu1vQ975PeuAE0Z2oL7Dm4c6htoiDUrtO5J4d+weJk5XgjTPRIOn65dqekIPo7oe3H+tJA9i5OU
bQiyRZtNXuBxVApdtJ9zx9XS6VwCkVcI8Y8P8wYmiItYS5oyt3GjpFPegGvTRJmVbI1euUcJelet
Ho5GukaXlFFNEX/DyHrcS1f/I9tQNs5ZBcpRY3/rC542hLfu/s9jFAJJIj4OFZrxmAmSKU9GOQ2L
92bjGLGGEH1o+xcnA7OjsVW6856PrIR8Y0S3xy1+xepa8Niy93sbAZ2La0+agz3VF/OL6AThBuHX
S8NEW+02gVtVBPcu8wSFEA1AqVWBPBYPu65WN0/HJ52HH+ILbfsg3vOeY9oCSetkcl8w2YHVDFN4
Zj3l/+K/V8tkrfo5I+jvSy6KDDbklVvsE+tmPj0UhV867gmkbNUNBgd3TizgOumnyebcFtH692wC
gq+hWtF5gPHMTh4BAAvD7AfSM17tXrmfrD51z2+dhorkyc8pDuc9IT1eVLH4CadrUFyqvAioLtmN
OhPkmJQ+TUxZkqYMl2rNqwPkmHDAZ4h4QBuUN45VPe+53W1CDv1R+FHzedhj3mnGdIZuVDIYq12B
7OHzI2Q+Rp8G/0nwM8FMhxJaA2B7oSb/jjnl7H5wsCKryjPVwzdPVXJ1uNZlsAINarym4jF/MdTZ
KM7rrO5ibsm23tl2XhsqTmnj/qGEtt/HKfG80gXKuGMPiDKXD8qUT1yMen2BjRAAqDxI/hlEAyPE
p85PT2DMiF5q7NHPuWUSHkYDJi/Ag3bp+g7lKXnAJAvtByJZsTrte2NiA2+PRtSpqkO92rLFFKrP
SK3pvMBo53vyzND7facrEE1hBlfrefNFM19HlOvy73xOOYp+o7UASia+MfFUmRiCo8Bs4mfC0Fob
o3JOfPikIMhH72Tu3OH3L0fqKM+FjVcYDo5IroEoB8zeCUd9yR+vo/ZO63oV1ZxAKekdPoYxHkao
dlAa0GWZx4vcvHge4asn9YPc6uGCJv/PqTSji0VCEPr24VBqZOBYYkyE9IKpFdnrnZwwr9wuWI85
z/DA2LrgKMidvt83jV10Vw+w2pELf8SxXdJR8DWSHyfloefvdY3s9JWeVb2woDvwn24QKTIysheJ
TdeCLNiiXZ/8GOAwZXXb21ALbTnpfQM7luOB61C61ai1CBL5FssUgP5ZiMQDNXyo4o6d5w4c9Kcv
2szxq4i6JPZz4cVp5hDWcORmSjtbjlwwz577km5Kd4F0upKB9R8ziFv6J+l+BapQhtbffo9cZyL0
PS3iTtKHr3D55UvhyDbXldgR7pHryZKpQZ/9UQ85D17BaQPPcW2FWX0baGhHyVpQ8DtqVdC+Z7FH
FDjTF2II+q9bblwg79qANP3S0WXIw9bStoLSoKqnp48QfJJhmIVY1naqmGiA1sg3mD5riz8SFhkX
pFbI2ZWJep2uLlBUY/8EufkE1u3iyn9cilTjkWIAfVk/Ltchro05ohzCF4/+gqE6hyszJuFU10uW
AoIKEv4AgExvQLa6mh2kJWIxQBybhidsAPXWh7/rNCNjxbH3w4CPrKw6Rfgwa80vs7hFBOC2Selx
ocOY/7E4NrxUS8d3vofF1sDKcqs2s79uQjHzowHb3swcUH5yAoXyubqWaj040Qmvdh91iy+HWv/h
bD0P+doYox51AHRy5k0BxIyr8abB9N2PXm/t1g56RRwaDP5WylIG6jE23JMa53kaKhyweva73LTk
XgVeSZVHuxhD1Gzu7a9CyQlJdYpppFtTYx0nH3oJQA2E/W5wDJCSu7Lyekrq1mMo47MZQvC4WGmz
6j1mIXHoW6EWwIJnwGyTKRY3tqeqUI+tjaPHJFHWkDAw8DDlobhu4z4z55ChkOeSax0iGnQWh/cu
U1j6TUPKHwYB0PWu+Jzn/uUaYdUtq3S3aezMXqGP0JgpnbuAVlINj/gdk9AofRVeU13R5c1vAz7E
6rpHH8VqjIncvyKMpb1XaCg7+q4HRBQoG0+vwrRf3ll63IRu7d/2vHf8onozx3XIJs8sfLnb5j1v
98naEEnIW7h45JUztFwR98la6XfEktj6h5cFRmI9c2f7rnT5TlGgUwMbbzqME2o36nLVjDuKEufz
0cS5roeNX1q2Fc6ElzfF9U/2HtIs4ccfPQAaXjPzrbDRbEDL4vi8Fc7o06QlmfKizx6GczT64tfg
zWlwhTW1q6/FKpciPx9JdbKsIQAQAbhLJ4mRnPPxMJLurjhKmmW6DH7SHi3OOL7WmQImr2auxrA7
ZPzDaT5gKGe11TezB0a9QtqQ14XswjK1YVrot47aZwopTycT2KFFyURZ26755YbjMhsADyE//uof
+GscdPOvQ75fMF2nFVxXcBZ3X0YbaBjkiC1rsPgBCCIXs0hvIhQbZmARfC9PgMrLSjOprjCBAOnH
6WCX21V1pAZVLNhdL1abA+8z1en0l9klsM2qQA1DxtsL90z/as1/DZ0cktErJ3akcPNKmsGItquZ
s+RgSLTk9v/isMExmmy6TVpFmfpW+UnC6I1UiAiiAUK23pCefkMA2qMCXjM9LnPme5WUkdDMw9Bx
+r1fRpZ/8bvBMAh7vG4hFOK9lA0OPlTl2CAXEkPCrxFgIE6h7Wj063oghlWP0ePoH8sm6y10h1h2
5d4qeVb37k1kCRcWmnm+A17RCaEdi46QK7/D83iB5a0Dp4bEUgQwYh6Vif0/avYnPIPtvE40NWUl
S9zLSccoRfeVSrhdugwYFFs5dukfNOw5pYf2Vti6oj8dUYQABBbUCfTNH77TfDGLnWpwpIPG7yIn
vpvdbqwSbZ68o+aLi9q28wa//oPHULQxwSRikG0930zaOCMMc2PwreCtzZ0kDQLzzpPeOSxG+vub
gZtgZ6qvWhSf834ivnZ2B4XApS2WPc2DI/Gc3xLsMlxyhDW/UEaGRtQKEoIJy+U5cdQD8q0DlkjL
vZebypxkhMHES50NeFHa872ET7BO1eangWCnGyoPY9UKO8Xesh+IIcv0InRTtqcXAot01VTXPOOm
J7lIwrHAKVCEcCSkwXsAdHD04sfSvkNUpAQteJsBh28xMIUs55FKFk5EKo5XIn918adrmufklFNy
FBZiRCC6cHljQgoxIMsayUlx0rdEzloPse4aMeP6WTMBl4KWGtI94VEliTebys3m9YKimVH69Ija
7xXQnZvQDI+VFJGBOINONzHZcUVvSliANcc42A3QQFAGpZBa3zMMTxx7m2pMplh6yctjDdc2pJk0
U+hU8283xunQy+eQQj6887WWKBV51gp854SNUiNXtq9yEABySK4sGRbD8z7MmCfOzow2tEYphchV
liwe4fIG2qMaHgqkCTks5XpEgYmJVNKWgPTKAj3HpJtVHai6ICHEo+65fK1LGxjorBv+Jcgoqjcf
wMUY2sjctE4J4GvmSVEhfcYgQq/neChyZQ6UDKOpmyp7OFLbXLMnMz+76SVe4ZaxPWPeNkTIYrsu
dWkYBqrm1UbhL/fxCm0ktvsYQUagMT+reoekdD3UXQIjBC+HMQ+AikIyKf2adJ0PN8im2qPG7Kbs
pkT/yQwVIT5sd7jMCxUk6pr99HjVlm/LIFfhBkPfD0+z+9QuEgRbuVI2FcoA06oPbEDP6BfrEyVe
jMDCBub8vvoNIoavzIYjnexgtgiU2jVQz5icS72S3ibI7mn2c6iDUyYnglENkGnksAANV4iWGptL
Pr/Xrl1O7FyHf9NvRvz/TeNr3GBeZ9mldebQDQGekRvHa585yjC0sLuzxm61bsAEBnyRhc82XMOE
t/uOph3CuQVOOa95XcS//iNW3YzNyAW8dUJnxdAMNqrZxgWDTsVNhhK+/kTEmsWY9UQ4UqXDzRNL
nAmdcaRD+fw98HALLLEd9vyrh2gfM+SB8HCUQP+mGQ4b669aBGtGngrE0aAdWyl/+Dvh9w1D2l3M
Wu4e9ia/Ggq13SNncMJchGQyu479Vdkg2noz37fzhImE33IL1F/qjp3KaCSoTrQfnbjPX6CALYhR
EkZgs5fFxVpQ/mveVAHMeR63gdSQn0W25IafJQ7NFWozTBxumzB3H/lZdggsuqEVuUZJqZCmXqFx
+IfpX5bVARaU6glVoFsDIiktLMuFrjppfZ4/U55NKAcHXNUHY9+T3Xu+9jl9K6K/Qn06VYZjY4Ar
do4qcOxD5qpSdJ/3HBcxr7J0aUrpfdU1HNNuskO0L8ilAHFdUMw7HlHgVDd93koWQ01tEe8vxyaf
d2gfDQfzJpcGPr6ENVypTXmm+qrK2QU9poRPaBGvC5Z+RUoz8sgHEp091FofJKuCK66KmAgGIUKo
JlBFPub1ygjSSkfQBH8v7qjC3ApNYj+lK1+EjA7juLx5oKFZG5YiBQulkmXk3wgqqgtOGtI4ug8Z
ckous6qLcNlZLU+WHNiV3f21TozL6/u2pLk5LwYr3jA4KBkb6yWXMZW2lhmmNugXdqxeI8t96Nm/
JFQLknOpDhxBt22Q0SSvfcEk7cDHZ8Yy2IK7jmC7Kxo0m2znDfV96Or29jLEwB+oG264mwnlTYo7
I+6wCQEU24Gd+WwLvXVzCwObo6ceSUEeFELVDg/SBQbXtGWRiPlIK4VW1SdEzkCF7etYZ2/dT8OT
TpzVTmN7NOBVjK8EyxGdD5fElRo9XEg9xgaNeeWBGG2pf055HxsXF+XNY89loiK2IOVNy3ha8CTy
vcxZ82tnpl3lLj4n9oWjRhJDyJqEiZrJrHoKpwSqkD5sYYhCTU8if41y25eEnLIqIyQSgqVCv39Y
3p+QTbezfv2Kw5pJzSPRkg0MqvfuU3wd3zzRmBKv5KuTQufbkKHyvjqP4DwDvrCWjclpxcvdoQMu
swJi7fXY1eKpPnzzcIROlXzPuJVC4Xoqmddm5K9qG0gREAyTInQY2oGrP1dFbA54QUDiF/slXR+W
ejwaYOKfPKuCf7cVAusr83Rt5ndBndgfWYO/GCyKAFflVnVEJNmb7KencLh7REnu68gWXRhYH8X2
D66QhqMY4/CBLnvcyJK6KwcLeE9WnrKqSTUOYr06uh0U8sU6GKduSxxLr8JDtAfo4Aagx6MAwD2i
6eo7trjYp4jfxNV3C4eYTQwQwn3lwO9zDAsH37pXobRA0OvSKU99zHRwCsF3STbS9398g1VS6Ftd
5K5ni15rJP64CK7GuI/PPcN1oW5ws1q3/cgzdhiCiNnD5Os6QaLxVPvCXCs1XwjdsObYIV0mnseP
x1rCOm+mPdRSZTDLq+mMwAzFmLZKBQQLLq7vUQNljRVZXcYIfEEuEBcpWpqfL1L71vmbNJmxPufP
4CZl9dMR59HyHHIeARrZj67n2U3yC5gCIXCb+4ziIzoDfMG5ZoiIkYlM1CKrb1DsRVRq9ouA0lM4
WkLz1ol2CZUYvOrw8+mc3zoUlWMoyaKkwolaCO0Dp0rzxi4TtQX+4NPffJJzkyEYKVge444PJd23
AjAovoI2oBZ7NOH6RpIkQ+TICYdmwoQ3BokPqJJ8bbMixllweJVc2BUCsDO/WWrCefgoRxkbAipZ
rsa/LhNZ7h2wJRlt6Lj9NfAnflyfacMPBg1Wibq4amHkoIZp6ZKIN8xK9jif6QO4wrbYrqqzysrR
mTfNjKRYL41rw62i/45xE5/dFzI2hReiYQYzjZSiLi0IrCcEPNDL8sXHpmuuaHuv0jvG0GjXSsno
a/AEIqkK6ee20Zni4S85eyaj/lG3n8Xi1OuWxu1cgN1pnPW1EkdTiktddJywAYm/3VYidrgu4Lvx
mbgXk0CIfhagSpEicsewZHDbJR0Mio3vePlgpd9Lv+w/kV03L1pXq3pYSkRrRJo3E7WtEtRJGKhU
92cbxj3vMdOw5qR83D7oAeqxcH5BBsTrsgGyes9wkqq/IqxBv6f2iNNeT/PevQjl1BhlGUHhokl2
/nE66O0EL7VJUJbRVfZk4kNJjwSv5u3O14mo32f3ngavN619QHCCp6h4J36W9Y2FGTEmoxGoX6dm
SZpig2EreGI2v3GUZZ5OKov92F+drHqP1e7uBtiK6fJbaNSjOj3Ic7/hn/AI3WhAEgPollcfEXkD
X6yfe4MHjK/LKrMnw+dxRzS0ZRHbWYlyG47NALqlDPvSOm59pc/R9buAfl07rbso0PdXvtVDStjH
iomaJ9eKhT/QfQPJzpNDTziRzVGpBDRJTOIzT9mY98PNoSpi/kAwiiLrgMIUa290B4AEvbHuxz38
O9pQKz+blfSheKVLYcxbRLIOIdtF0pXzkSFM3bkgbegKY1P9X/TBrboibM5YoceMIkEzuKYmZjhZ
Q24rXzoDc4rI9doSotgbejHfVsso9jgMFpfBVkLurQCOzBmvP6kuNY+xfSiQbYTBVMZ9P41XpFJL
z3eKC8dc2JpnKxAMscGOWkTyxPETsabvwRA+mGYO10p+os83y9gUz8Y6i9iADF3geBeHIScRNwSK
5VMhqr0PPWM/c3fRNQqdpmM+FFtD1Bdr5l+5G/YG4UIY76TnM6mm4+DLqj0m1RZ9Vz2V2SAae5+J
02A/ZI0VnnsOinO9E8AMNF4rCFqw7BdMQ0jGc5jgSdXi7N8oTrZZXMPG4J9GI2JHTN8mNSFcdY4E
5H8ev+BOAeBkiO+3hv5UizrqA0vlctkQvBOS9/wBwz+NWpyJcaoJtcfvQGAc5CvpKj8Y2QIyPDqS
Z+cLrVMbLpbNfkrMAJpDwfOQqNZq7+XsEcQGiP+m7wb+1aE0R3P02tExp+7SMLYhgndhyQeXCq47
PUk8tzPAp5Fy2m7YImrKfcr8Y4kBWjQiIDbRkLInfMjRopxWx/Mh6eNyTitCC/SJkgtGDJemDLVu
NDpDXRhCOCTnb7419NWyYDw/phqhicoVQ56jSzxOQ/OLmaKqkm3Br3lXKzsFkJax2VguobxagDl7
HT0MpSruHCYCmvdtxBm3twYjwOvG6/0V5rn9KdOKeA4cj2cdkZihe0RxQS7DRs3rrBXSyi54S/09
10KXhS8L3xlU5O5AJC46JKPXURQhFnZlwuMkHCYhSAnEpu0LdAfCKE33ISnwTShHX058zlNYHich
cMyRZs6/NuJwC0djkCVikJbf+Fxl5Kj1FPbiQZuIPNEBUHNOaolArDOYuMwNVDx0BXY1iW/MEQet
FvoPi2OWSqjyH/dQHgQRTvN1IkqIRUpaqSCfFHaED8JqE7SUDHGC2FK0Z1Re08NiAMokmYljwbYA
48KwgiXP/CZHowrlett14NR6WCb+/8zX6BzxxfPAU2dILGIDucx8l+IcxDexyVT/4+mqBgr/Hzi1
Lib963fQIs1eLClpJhUvGn9RmVZq0ggCT0viGPVncNJKgjcoA6graifKkbw6Tf/F3EY2F7fXqUsV
idiPdaPPPihYuYinBw00Avmz1dvZWkVfv3sR1vxzVo4NqE6skL8HlLlbM+WYN/FxnlhKBTo9Hn75
0n/h2Bg9uYgdu3/WsXM1NTScwBMfd6Ex+YWd0TGmamXgcnH6KAjoszq3L2v5KJ4cjah4GbPT/vbx
A2xp8p5/HhjQgx+OPHezunu3pGrN73s3U4WfQJdeSkdUbtKUHr2IWuC+JnpXVj1+oHJ8sbmGYroq
QN4OQcAmAtBDiehMTz1eFh9Vp/JO5wOq5vptWTgXzUmUOBBR8Doyxs7LH6fMOVIV+lxtfYNobfMI
NiYknnmynk+XFdd+xX8sCGGBW+1nN2g6k54PM5aAJjaCYSj2WClg3RLywrUoZUpDK3CeIhpexyfF
BRob2QfqX90Z1YbMcSu98Z6VkDWrcittsL/PUAMlLFlNM1NHKX9gMryHexaakrQQH6E4+U0NSA8b
baKssN1l6SYtx487aUVdVcFXYmHbks8D73WUb5ZRbvFQzJiwuDAhZYZulXOihP7Q2j5XDTzB7Thf
vBb/8YFtgZIRtwjM3EWdpkbNLpN37NXY2tG1JiD3qoh/B1thVR121LDi5E1bp/xnMvgtE03rbl04
eqpkGHSUrSlbyZuYh7ga06iVetBaMeHtV1l2A9YExG4UyjxqS4zQfZI4vfwwGeiSJW1wMnBMuC+X
VMYS38Zg9tPeVyeWO2LHbiNQmiD16IQ0VS7Agjtbk3jPw3zYE7tG8DMT3L1JY19PnE1Xq2DvJC72
oySffj5pv7heQPkM+M7nismMTxiXomdx5ueu6nY+mlfiOQ3Zu7vDpDd58UAl+CSbWhPVRJk5iBVb
TOfAiAWGiUxrx2HcWV8hpzUiWiSY0zRp6ake2AQNns2+zuqYZt7Sv5Ux8Ck3HDn2AJeBl3BNCzns
D0D8UOQScfFw4H3Kf2UYQ3u6z0/NED2kxzmmrZm3Ye7Vg4Z8iXWF9Oz/REbhwvpL/krIFIK4iA8o
euJ3TUMkHM1cPE9TwV+dwwck/HeKJibAyVxmhDpCvmPQA/UB5LLLCaqM7GsAAmBS3RytPg5IXaWk
7XFBKUZC+sSTXP/Z2E4C9/cPu3Aj9d5G6tlTBlbbAR0bwXqFh5Bff3eb4CxFGx3ac2m/Kx+XZWUd
JUR+VIJXptCcf/X7eVuzUSgm6katB9BwUVlaC1fh8pnFBgEt4Yto85RrOw+qLC8f0Vmb9F7V/K5v
eMmIcOPQGar/neSHqPcIBY37XmqzsRx3YnrK2CfVZY8NuOZySHXgOfm7Iw/ylfs52nA8ePmrEBbz
ejKIR7eTUxyd61qMSQ2vzbYIV/GRNMDFS9nF5PGoCbW2n6qv1f7r9Mv9fAQ/TchCdcDFP2V28wfT
lHJpUJjuD3aTOdu8a1+g8z4BXMCpcRm61m0SUIzFbQG6/WLiM6prlXQWrz8ZqmFI0wQW7NhyRYZC
faHGOXHmg643cAotV3rIxg/GnCSda1JSiJghY/pwnJ+UAvlj+dZvKXyKq/CjZXdB/K+m1/tStW30
TcK1LL/PfFFS8PVl8f5FiJH9WV+dD5h/+F/rj1yWBGjYcAddflqKmVGO7xT0CUPQT6/lU/N9w6h6
HOaaT1QJiJgWe0ebyZXjC4gdZvbSoBjdpKtqu1f4J7mRuhbnu87owyq0k6rn9PTg03g/DDMurXNM
XHZQo2bI6j8cngKAKaFNLU26NghDNMnhc+XmCapXkBdQoyqquTk7/K+tW2Fa1tYhMOchvdcBgTqf
jD1Ot2KE0dVkTxBASyJ29+TIgW3ZfAZGEe4XxZcbOgniky89Jj7G7U9qUzmJZ+6/gAxL2yDL7yEF
BZndavAn65yggxcWO2wJ79MbIqp1P20ceWDLaKRuJ3MJOvCyUhxku5gZmlNj95Ip6R6dQvbG0Ukg
ysvqKBLSOFgL+exZXwznsAHehehBEzqCgoorI4xudkI0zfHOTC8DhR3kvT+BhUVK7sEt3gnvD448
yBnIyCST7MS1vI4gl1fIBViyJookhBZPQ0JW/glt5Fj9TXqgHykJeTsDNQyquXy8uyDW0fxI+03m
FfvtGj44m0hzqZwV3sRRkrfw9LRuAKG6Ufb4Txs3iVgRYNnY5ikt0Ab/XvzcVs1wox3BpHmpdJGV
2uU2s78Rh3XzXm+RM+oX6ckAr7jUPMzq+InEACHOSdwOesK8Dg3YHDTBD7MTcIPY/whalaCBKu5M
PB1Q5jCD0dL36t4WxyEhK0iSF1iNdxchVVPIkBBsa6BJFXSo6qNBk6ipxUUvb0Tg2LqBd7a/QKKS
8TSi6PZEfYRRZqiuO9kBms8UuC44xja8ujBTWduLPgMBNEZ1RKJpf5sNJ5XQgWPkjqMpwmejItH5
dl5UCsgRxdKAEudWMcUSoqDpen0qA6XpwuKgr8+OemAqfE8TEEmmYPt2mUxy2NFa10zLxfKMkfmc
KB6wYucoQwUwcpQgtCId8wgmPgqoRxgDV4gc2L7J4q4CRfutq61/tq12jrXTDs6mAWDPzoTAB9hY
U1trMRfnytUlyRj3bu1ISz6rqEHWKpCBrp3S6ZAYkNsyYc06q8Rrl8J9k3XlcSu6/8k7yBFaSZWv
BnBv10ExDg56LOZSoqOUnTLmaFkkyKlnSHjlZft7BVoq37SS6KNw6qh0oHo+ynxMxJjyMGk3HDxy
ENDWm52FvX9XmvEdvbekBp8eMu/QmYB3LiZM88ZUVJ254gX7Z59686+a9G5h6zgFbZFaOJAhB25G
GQEU/pe4vsOUTcifjT1nge3LwWqFn3ZEfJvto+h4RaL61eAjZZNqORBAawwUrSkQoh8N7bYL/3Dd
76CxRvrMHEk1ZwnojkkselIClRej4I140c+mSS1HoXyrBX8/+W1/WkBWjwot+JuAQr6sDSMFvkre
BpP5blbt5D+mnrKJciRqLEtCOOqFkgdD7NSgh4lxB6PisMqFHiibfFX14bDai73oW/WtsmxGYdyF
eYkbcIxWdLDtZPUPYTGBJyiHN+hf8VQ+2lKyW9K+/OubyfrrqZKQd5WDmWodCGkEbovKUdpKotu1
sDQxsRS3zVog7QbCUV4uFYv6xt4dmw5THeNkAJ/bkPmxjNDMzdayiz7+HFgDR1J+CRekvfvelXPX
rMZhZ9/PcH9Jugn2/VbaVoI7/pePHsp06TaP0zxpQ9g06bzPguxlZfL5RXJqnlmdZUvOBLwL7Mg3
xSIH5E7dFSK0L7jgPVyP/zjP1RUcRLMGhn5s5A9OzkNDU7GaYJqSCN1UJSChhQ+0jdg+gmj49f90
Y98ViO2ncQsiGOfrdo4iE0QRBVVBWf/xy/eBOZ30gzeDaS8kjv9O0rMs3aLp5x+JcNJPrkrfB3bF
Lou1X90+svVRfZXLgeP11maE/PTgDqRarA/whAo8zQw1wOYiRyCZKwEQBpZyr1CbUOMSgqTUNm2c
GPQAV8HeOildGt6752r6sx1+G7yVoqIcPA0ig9q4+qF51MBwtOL/F1GEe4lnRvw04P2T6T8B2r80
mGUwahu8rIkkdbnWI1YhwXLaJdir1vEcc1UIPkSet+HntbPOSZ+rZIwGnooMS2NyS4t2UpGlaIld
XSEs8G6g7NsM5EOmTRayM6tncGNyL8jcWH0ThjliflhEKWPxez271sl5jy5nZEKMtMKogtA3/YS+
O0s24DrACs+e7RXq8pzaiobO7EC7b7Tfqm4ohQ5nwCJ9R4sxaHbn3O3f5MwGr1u2LDiHOWwQEDey
bT82oFqwtwtwwh/yn+BJreyyKejRldH/GnKrUc45mg8ULkHGsTA6I7f+RLTUXGJ1SEBCvgnMGHtc
K/5lP9tyPPgKuhVkzx+iXf5DaPUX6+EOU52bNH80uuF0+NnPctl8vEzX2uP4+pK5MOFUeb9SKWGE
NcehzntKkJ8aFY6m3IYOq8lRrydbXYos9spV34hD3ZUqdgJtP/A/RW52ZWXmM0F5rDgwce/eIuOL
ikfvBH5G+2n4eypTHgRRq3cCv1HXOq3EpWaoRjGP3YJV+gWKowmsMJ5IgxuIMXfDeDeDq9ETk2br
WFJz8z2gHGSQIfDw8kGjkYLx8ddc9CuzBhNO77MqZonVxJ8CjJpTkpBjqW9JvuR/n16Ltjed+UZ7
6/DvNunVO47CbKbe70q4n5MRhISIxZgwUlFLcB9zC2R6tJ5zQ40PHJSQbrZof/pSWCkGf5xjSGCD
FLZpFPe81xmBfDm07Q4jrmgu+ZqZZbvKJGl0XUKVBmdyd3RWtsFUEYwjf2Vk/OhN7V0XPlWFirIm
O74Jjw+WjN1e3GAj0OZyWLxqJWl+VE5lZ2EvmuRglpnXs6J4QbEQVZ0gg2LmWMDAzvNPfr5PKRUD
pN0WyfdBNOkoj4klWbJBKLpDtb+uRTUEbzVIsyVILxln7cbuZ3/Ik2b0JBwJD9S2ECHAmXul4c/n
N3p7sj82Ulrm9m/5T+QO1n43mLB2WbDMNGnPwenSuGXYX9tPwPJT9FSTMYppTdHxWTbdhpjCGr1j
XVHL5L2n1T9oq0rVTp0+30ntL5f48SIgkJN4YGvd2tc4qThO7q25gPErit8wEBJFgw2WoOI3UugH
lAoEJkjHZmGUX3CPCbHoQSl2HjOPGcAXnON1V8L8kPP8yQa4qXaDUbFVGT8XrrZ6+OdMH7BzaNjU
AMTEFfg0KztRwo7eKlHhaF/5Ri6QJtZNEnzqqDcAaBkymEEiB5ouwHy4SLj1ViylZlndG9tfvF/I
9Xi8CWVWwzynorIb+PVBes/j2LP506l0Ev9LeeJynw8+EmDjyzM1n6cSi88sl1tHIww349vEbYyO
878ZvQP9W2i246Wmu5PtnDuxNnRE1FTxBXYfhvKqIDCKZTF5a1uDXFMKx1dLNXfftb42yGXky90b
3eoYqFt79BAOrbmBNiHZAyeOFWZ9IXQE+3IkQppzOx4fr1hZ22NwN1XUyV1v/Owtepd4rdcXcgbl
XIrFSgfFbKxdCwFnD0eVAzsxTry8ccDOaLcLQplHWma6y5UnPPQZDz9sbvri0A0t8/trHccR4Hc4
uTJSGleg0w7NZaxfUaks+75bQ1x4kJwSm7WCX5PKr8vcIMrma/XkeTQLxA2RsZWQMvAG+9Fr3POq
JVQJqbC42N1IEkl2bzSqJeM/5L9LwoKwc53R9u2/4M09ME4vjtN1W8WhpxmUPqx+0hiwRCuNxbs6
mTUiTt9kNj86MNsSeZzam8fmX3ddhpst0QGeJ7oQUDRwn6xMz9AS3fD8r6gU8PWhCRKEwEXlBF7h
uYRWuQqXs8BZSoksr4zuTMmLchdm5MxKCOIJxWhVx4ZKt7YXbHGLxfiq8aDSbywKZlwNHmKrrTPs
e7cY3LgPv3EnIiLx3eza29RaOTN8gq+ww6DdWdcMKOhz/AHHACBgu4TGd2GDFHX+hTKAT9OcW0+4
qHcTbYpcsWR9rp1jZSylP/dhgvhFbw+WLtzdMvxNJO+veanEEUk29NI6OfRMKzpfV47CeHw8h9IK
iKt5rtk+uGx/AEY6conJNRng2K/gtiO0gGbcvuur+7kf+ap+J2XYEIoE+U517ihzKDzi4HTuypY3
4OK8NwagVVhSvOd7MnJo0YgER4D5kw47vW3YV5dOT9QqstirUaZJkc9PWAKX/HG9ifFX5Xm1MhZG
u+FB12qHasQSlNSYlhLCGPUq+kN0fEJ4WnwxQz9dFIeJ6tDIAtf1nZGm1dzoq7fdZaJJE5cIAuYA
5/eR1HV6I+FvLSeMRloHs9F5U5VthB5q1VB7yxbZS6Q4guD/hCOF8lb9/IuwN2Guq7fdAHMXmYO0
y7lMvItOVIZTh2avQsFlc/aCsaMWZGTph1vC09eDIe4Z5jUVWUoDFNuvv4STgHu8Znp4cDeCvAMK
+vGU77xo0doiO2DYUcFKOLf0lwekYntvkBzqGhJ/npekvcmFCwkU+GjS/v6TYmVugICL4OWRgkWO
Hl8i0huhw+tiOAw/4607IIwuLrJC0dpzKF8jWeoK0Dkez+SOcyvvqFqsJl4Pg3MYxfkrrNitGAnS
DIBVQluoi3wCBXTzU96qAnEgxbXlIv6wjiZiFkyC4lGmUKKFSWeXQmXMxbTplrgp4GV5XtpQgXEF
sxUtWT8fcnKa5CGa1V7V0U0thcWjIo6egccvUseHio5rf95ce3rJsnClt0oe4EBAzsWGS+HU1AXV
phW2bDw/XWtT9hW5/QdsZswgVmSSjMs2TTbbL97GZx7FY/GVaMj4hZcw4aFR82V/Clb1ZM+P2YcO
AjdyRmMAzCpl0LBVK7J6qVGS/VX7aCrv/TI6kKZN+kZ1n/g9JjwtN95/+KnCkHd+mTc+08GyHQ6X
mrIpXQNromcoMRO/FzyalCRlrpF13Q4anUooTdRXNfcnKlUrCRRtcABUwJemKLfmMGqlRXqizhsg
mz7BRetXcx1ELLsnPig/ycaP1y+kIUc9cslnnbaUwj/uR6GVnJHFl+3LHaGlsjI8u0W3ZgaSnNdE
p1i7ykATaBjv999eh7Cl7/NpbE4Ar94JG09NtarodK+2YDYBfT7phuoptJJPcmDMpjiYQFEDbwRY
rK6nhsUlE3IvlSQXQwe9e8JmF9HwqE0TNvjSpgeQ0iSaF6ET4YNAtSxqjBs2KVfrZlR196UFyND9
37w0hlHtx38fQM5minLC4A0Ad0aHqiNq262RHDmjSOXG47iR2qfTZjGjTVYYkuOY8oz6HbMBEpy1
wMfBH/Nimk8F9afCHkaViz+5SETzOm7pNBn7NSMjM779Z8i63UYy9len2fog5KF/Ng1goRqpnNiB
LVv53XTrk6ebjensBCkbAE58F27aa0OQN3BV5EtLVIdTAgdgMBmoUERlst3bP1aBySouBWxGclfK
m4o3p1nkQbxV5ej/QEBU0QWE5KEoAsO6xv3zUIYNZAR0Hp2O6UF1cDEo8jMlgAfNsQ6eJRUu34/g
Qea57qyisTtdeBeeKZRc7T2BVJqn+I61UwNkjQd886NdrfQU8+A3yoVRuDl9oG3CAG8x2segTUya
VTYdSF+FeG2r0z14Rswk8tKZctkC68wS5zvc6YyZlIksIZHbYuAMaTnTIx6rn8250Hbj03+obDRj
eIr7V0W8XxCUWnmb3LNK3H4V7vBndgwAFCRRKCHPPd/9L5q6C26hTNcge4bhObQP7Ex8XCcoQq5z
lUDGV06uEXsliFyfkXQzM0itw4EBM9LM+lc+z3lgoW/I0psGJ/Kkh3/u6W0i3FlcVMD8K0sBfwWH
WO85T/ceOyY57EE6LzG5OY1/oDo9MXFU2DaKecXpsGmEGafFPPorI3j2uteC9oCyMR66LFrmIjJQ
SxgL69KiDe0mdi0QBsbeCF2TdndjL6oRQSNVYuuaQVlmT7c9zb6g8VEfkcBsRDCt3TjepON2Nf26
FcGz9shBRXOVu9pVjXFE9wIXkvsTSmkQgyDFF4bgJ2IFhFQbiQpGrCAIbGESiW3TXTNwoQpMuNHs
BJzmuhq/8uafgBkKDRFRzRANx0XsdX/LNQz9X2cW6fGKrxN2pVIDGBFudou+5tLrUr+EAf6pUmIU
/O9G/eM2EK+Loq4qYMwqKhcoWyOV2533n5TFU20fRtKBqt/ehwvOIFWclXkVcEBwiaFSJARW+XxN
92pJfmAw028C/jjgtlS7GHg6mgg5Q8VfLHu92e4hCLQmuwPUR5nnOhjuRZ9FHM+AJviXXzGn21p5
/QYOUBromq5+bifVvQw+WVO0s1JzH+amw0T7bNLstDwRieMg8GiqNHi73hxwSJQEtfPQBq25+iIB
a6jca88vEna0queTW8HA1AN1LvD9Y2O2m7GZXdNtL9n3UiucXD3oOxzKuzBgx3o9PmzJ1RgmxTdD
ChT165VXhn19lfJEjYqwt/nj0uddIUfbTVR+PUzjZF4W0Eusjt74AyeYDgxSFINvKMkEsfXormeS
aPVzzezdAGl8SrhMFWXC0FD64Rilqy3fCSZKD/sQuoeu8eyVokByUmLQFlcuYkZ6HImDmq+y96PF
bleI17oFDw3MluQ/darC9ndEK8K2lyMaS5UzGo2xYZQzRtVfFfr4yxUjN2T/zDzOyADlYFs23yVH
5DPzraM3w1Vyr5qJw46agoA+10INPvigzzhWhJLQYEVkgiG9H7PDAQOXKw6q4QLpLSrGu2mQ3Pki
+3B6QROXRyYO8okzrVIzWGtZkW5L0bhkHMCqGEn8dORPfjAc7jQ0ieIBnjLN8K+D9A1RH6NeDiQS
BPX0mwXM3Y70Yu7FP9qRGDb+g+ZExvO5JOrfnA7eauniqQcgwIqah+FQXpF4LxA/ieBPZYJ5iahU
rO4cY4+AVOeogp89DvXHr9SxWuVjdxxORTTQ5ppOpACtwHsI4O+DM2JDb+8KYNpaVeKyfI7DQh6F
iNaOP6TrmRNTKFhCyb/lKlrYTmd8OxMHAigusE88f7Jzj6D/oZsdQggi+HsVSDg/lEZHlgcgh7dN
5673AezAG1ZCSpWIngUK2U5kodJqp3BO1JHLAFpqA1oAoUGT2NqCEAksghYmasNkb82x3ukI85CN
QjCMixY1O24YgAKpBPlVWnTMu/eHsviGfGvwE6j3teSuo06ngvcusRUDdpBcOmKMiPm+cj+Nyxzy
WllkXQAb4DIYvb4qz080dhwYVezzEKOWzZJB7aahHYVnMG0kZmu3Wm/nxoPI3Hjm8bAVY8A1G27U
/3VK26GfIBX+G/mKhSKDQAIKmXXAWpwOkKoGMDug3KAsxNwqxrchBqFwKxBhIzZjJl5128L3SDs/
uZ3ZPCH0w+hJPamDG9rfhcccWwkoy8DCJvZnLn+SihJ0lAL80/s4mooCtkk+R1xILwWTTsH52q2Q
eqp5YVDVR/suUhUVIwgQofU6yTlLxSWMeV00sPcwlro90w8c2UNhTGCeYDyMY09Q0o8cGcAzhZAP
mkdZYxDF+4VHkAolwOSCj8CDTVAADe/MqROe4OWQjX+dqSrVGtGC7jC3UUBC1eu0seMThNmjyQWl
+LBJnfY/PLBBI6EevkO7JaQA9AS3bWRWBLAmzYExYiHMU/W3Tvwctoga2QEV5DcRpH/qQ0hCmOL8
DYJpbHmZxPv/Kb2cIBBpNX/bG7Z5ThNzzH+FFLMd+eZ/dy4YBIFoghWwxPZv/+XuasLxBEDtkfdm
FXd990Mv5ibp86AGHqfBdFj3a3ZaQXSRRTT0TI7170Qa4/W3qTWG5Fs7MYe9Mmo7ReMVtZYTFCcN
3E8Q+XgNij60GSKx3e7kD2GHP+FrEKRbhneuOWPTH6CZUqDIKF3oZSTpruDhCqlYeQoiYc/bJ2Bg
Sd1ePdtUCgEjyjf/DIs5lbQ8OStfIA9Y0jGQRwDQANnraaXnNeAN0ExEA2TuJdAjo8cD4dYP5ef+
z+OrIVsN+LoZfJkGBMb+8/g9ID5oxuvszeKDmEPUPg5P8ug2U8Qjw+gOQ6NPtULTAxORDwhOybHk
iUrwmwK8Cl7Eztw82JuVZbNpKGuIGC3S7oh3l9VWLbEU4GMZqhAJw+0rE1ceV0TWshai40+PW63A
5w99uW8c/VIv2QiTVwgiaNsM9aIGIhec0VkLtZstKQJPnumYT4V3Vn69VgMqnhxUtD5aDu2Fk3yS
o5m3Z3GrpIZLDqUoLpgafSy1AE4d06+mLPDK8qBkN8A8iqfeYZF3QxK00Db5DqgbXltiv08z3PFQ
hDBLr3SmZloKONBlD+IdksHGKp9y6ybfR9aekY0jmzWXkGKRjf1B3sTnl/AiEPCgHutxVXOzMEaV
qgl9wQsyu2T98JzVh1TKb95QRC3iYPelCi0V7MviqWrRKgN4nh/7vyeajemcBWrG3oxXRXyBlw4g
M/4VXLXgYDJLDYT+hLpnKKRoBsnd/1CgPBJtdQH0kjjKbVvYtU2g1HKXcVbPP4IugW3gGqbG/Anz
GoaYnQNVB/JDqwjVxF3xNLsv5dgw+TNSyv4oVRtxB3bc2YUge56zv6nQjNsKDJW5KH8JRC8hj3et
N1aRESphfRTsGPMUyJq3/+1xSiNMmBdjokOqzcnhTfcrYoY9/3Ao/oLP4Z8501Byhu0GiXq+Aez/
214xZa0LjsB3aA6pgJeYoc81W4jU7YDoiEQdWCzShpXNYwV0YeITpfJ1vaQk7RuIAK5pqelD9dDB
WRnrj4RJY2tIY+OJDaQalYjBdJevY28cgePM2vQF4UGEuwiJ5CwUIgDB1+IjqX+uEJYwUwvYexPV
09OHt7tTTIqAdJYf/pM5pXD5vdmi51yWTkqFZnJvQJQYxx4NFrN6hfNoVLZxD0V2TXj4/Sw09aCh
mwo4eoG1tF9GrJbvnJFalmIscDBfQUPjyCwCYPxLAlHje3R1GDBneYvlDMjizRJWecTegcW7Hev+
RVU9AHXrf0Ujo+Tk74cVf12DplfjiMfOgZgCygmsQARBQGXt/xKSI8LKi8rKjG/8PUKOhz1YmA9v
leP6JHxmDRIPM2RqX0J2WPfwXtT7cK81uhiEF1sESmvcDSgKOCBELYT//SFjwB071n71oH62CDT3
q1e6xLWzqeWKCllIgmodKIVxS4H5swrJMeD54gmG83fuMQgCE3/RWIRROzx5iNGb1Kq/2h9+zjml
tb/dwOHlsFmOxJ6FQ7tWuoTSQWOQz2PZuECHGEQy7gR9fMn8I+gAcUJfyIqyft3tk9YcJNGdSbKN
Jpbncu/a4j5c91gQvvdeTQTWZmwDV0sXltnoR4tsRUtjX+OSsSvnbYqjwuYHA0cH3IbhP/DJhVg2
fmV/rEdR+vZPZkj0KQ0v9VZj9rGIMJr1Q55xV6PlgC0/ZYlJBZm6DWQlHQQjyBIvJxeGYkP+FO7h
0uXH9p4QiD50TZdnMpdXNnViA9l1RcA5UcdnZfyvOBEPFGeROxjNTxR0CYIOpLCbgJejRZ+aDoAz
1SrNoxZW7y9drW5p6UXrzKEKlzd3EPAY3c6xKugKISfU4nygh8H0TRIE+g5vWqqmfkmBnEiK7Xl7
2EWSz9aHXeX9Y+1Mr5Jj99JY8xPyCumEiYgbQDst4DivehfK57eDB5qCc2uAUr8IV4zc3QmpE9/q
FvEMv17/h6KZk9wlY/bcHGUZx7YYfkRrCMhuyhxAHK754gDP5DFsBfPxtH0P7qJidqwlMh9fnMyd
C+b3jjllTzH1r7BJ0NaJLzVP883HXehdf8RwCiFxAXaXM9EJoSng7rj7CETv1tg85jc8e+mtjowd
4M5ANLCn2nj88hYE67TgX0yQYGk5U/rpzU53gkWUlbwpE7JuBICA1TYnTGo8wx7gLtpeMBEXhOEo
HbzePNRdqavXQ81IdQhC8HEY0iQX9SaBg7E1z3CbA8JyNJxPWh32801FncTOZMhx7PrgOe0m3Xvq
fetsW1gdslc0pJRERWnDe8sjAsqEhs2fN8W0n0lWBI4892dHJVfEEyBStz79H3F1YLnH5zOisiTP
mLPF7FVUUZaXC1TSXvIY4ibaSKdogwsInqGjEu/6/h0HsWX+PcFQfNI75O5CzGGdoQRmrQZwDTwC
9JUkRsDkYou0UkL+YOcUBjKfl6BAxZI1pQNGwr/AMbXExqyGAxAARubznI9VnKzc0gD4cZK6dN6Z
b9gQxsOcvdYrCMuXKvohIZ83jAUKOfJdSOQ3HK/o3yQ+JHnJM7eWzFWjzazjtLRZ4OYksaZRJZ1Q
RGTy2Df3BN7aEjwNQZ7UBYbbWhDn8+gsukDwT/GOfNzmzkRacdJuFIShWRgF/w3AV0ncsBU9Kb9j
eFv7jkOIFAvptvf+qL2Fh7E1LnxslhTukcTt4phehnIDVQcy5w8xrFsptd9R2d8VSL3L13XpT/iQ
3fscyTV+oR1UpCd8Ghco8pyk3dvudME1OBfVmC1YoFzjiWnotFHXRW71xd7psy01sl29iW5g99it
7mXUNaYndb4VMExl2MEfyrBAL9HT6yQXYDeOMg/44MYkIpTMmy44fgQv0vcfcVgoakd2gU8S3MPw
Ten48ftLhBnUY2C4BbE0+igUsSfxj1aFvgcIXpdeJPcMW9yb1hxO1SoshtRDMeQfftyIf6LLQDAo
N//uhs7vHFcZ/PBG0R/umr7d1G3XFmWhl/f4jL1i8YQo6ONykpUtb0uvYkr3MpxKtErE/d4Irkt5
lqKV3WVHsgPfNdngJyzUvAoZuZqm+4etb/v9x/8+LVhpz7DKvxfhrOBO3AGu7Go8vxvqsGOk/ot5
Bm/LZL1oyB2VjxpoeghdZb3Z2t9gvt/2ZyYUuHbyr+UfEx2YO2YnTxDmpaICpraEJ7h27k/QMITi
05+62uabRqsu61UNNPo75VPq7ZyvLpFF3wneHKeVN5TjBQ2VhVhB1jwxqeSrGexBAmhGeZ1RLtci
ON+W6mfP9DeTeJrvBC1uEcLMVuTGoN98gMlPr+1wWLM5/JP2e4vOwXIRaChwxTqVa5a9XEL4TUmZ
bM+u7dBIQr+yxBApytlUQVxy/EUkP/qy8qZdLpfnrdbVxBe0nqj1wFHi6NDt8BIv7axFt6jhw+mA
2sxFXvvtivIiC1MAid2v33x5u9sLLRk5OW6LQzbRvGO4I98q7NGDw0/aEodome7g9+QLXfT8o+S5
UwhuZVQ+8W0558evfR1L5+n3LczQVxH4CA99GCeKdic2XEPOCx0zmrayMdZiDlDVDcsSA11s5BIS
Q9wYhOJRia4KCBb4uBA93jYhT3sMksl9US9Aqt9uMQzVQpt42QPpPbdRP77hYv2K2RJ7GwnLOXP4
p9359G7LUd61h6AiePi+tq7T5iTPsmX/aMl9ditDyVYNxrwqy04O1X+3UTwNNf6AzdeMcdKNFGGS
A/R9CZYe2HWez7wVYBhyQ91xcE1Vl29Zjfn0ytX+DQOypGWyCPc8cykJrnmGMZ74+Zvsgp3qmkeW
ZRkwjpTM0EoQK5tV0D0LGEjsn3JgI3uNQCcXGbFUINDqEPf34vXVOkbAxr+E6Vy8j9VBrSEL96ND
D5d7UPtSfT4WUafqrvAu8EFHBG2w2lk1NCDC5W5ioi8KhYzI56sQJrUG2ytSyT64N55nebzPIx6K
SY64O1hGuym7cnrm7IqS1VStzLO2/Q4lHDWjRo4XnCOSvuoV1es2dVvYsb8K4qAHxduQF5tjP5uU
8Npk5CBTzP8yXSpH2FZRXRR0A+yUUZvsgA48B4vwvj5TPWMFEpNc2aa7mP+FlO/tqqJ92qE9dgJk
ze8UD9M9T0vDGIfMTKln/onfME/loKKwXCeSi5lfDLczhQzzS4/kIM7pMW51e2uWB2Sge03Mg2LT
tGm9RC+NSa/tX3vzff2IlWUpx3hj9JF28ooxvlMiBsr9l5YwWF2JQPGAWun8WtAb+OvYDkulJGgt
wunNevededN2WRvk+zAzeK3fZRHhI1yUEkc0AyT7/CAlcoaJavPCpuhOmZMK2KFXmnJ5tXiyRbzS
McY4LYwsAq0vQjyxYTwCctbDa3pcAoMRYkpG301w/nblM6CQ8YZk2tb2QAei48GiYni7wRqyymns
UMyL/0+QsKtK/mi9Jf2pruZGF+mkTmn/kW0ERWZGVE+LA0XyqzHPt05k4j74BLdBNwC6NQpMuqtE
2hBORXE5TcokNMeEPGKxCUIquWm+GoulVJt6X8U5Lf8zUf1ht0yJ5pA9M5z4I/vytMGAeb5dBCKo
BgwFO43+Ske+YfLOuVxAS9uTZxVokn2j79wbh4d+0RwqUrCU+ZtX3G6wRM3ZbtDDn1/cwqqXlQ8M
iLwOZY4mqLxF6qpxIo05yG8yju3fUaCgfDE1mgj25u9g5+EY7Q69VF01HIEJ49vSZ79ynjPCE3sd
DOk3W0YDUId5gZBsIX9KAK3kZhWGSFsolBE3ffVqkyniJy61gr8PBHW8uwnrPBSDVOTIaXQkViZo
AYuZvKYzNoIDKprfTfTuxQ7Cl4ygZMoCFu16Q2RBkLJefvhaK8IXgJ2a9aHxaGB0qD6WXFMEctc3
PPZ01cIfgtylUyBR3Hf7CrjijoJ5IWpzcahLPucp167en0jmhaG+9cy6OiQK/vTpE7Mjr8rK2cDS
myfjo+zYGvzsd1Anf2RVykWS8N+ssWqJbGAN63qcOae5avw62R42JMlU4oGBz+u0P8QlkIcRc3fr
KbQ9c7iUJoy14UUg4LYD9MhIyKUBC2fJ2MukdaG7yloaCCHA/NCJbsPAJ35ZKsLDVaqYze6DZtQZ
T9Isv2fPErKwX9e4y2HgdwLi+wHXYQR3C/ddis1ucSMJb3BxcM3Vqma2tv1O2zTx5ezOd1Kl4H5d
cMX+sDJpoB05kRb+DfAkMyJFizmDbbEfG2f3XQ9GX/rZoT1oTLIEXqg1uK90Qctg1tUyBox9FHFh
Xt/IdgJZNsnvxAkOcJaxYkxdZGG30bv5Bq/wIzhm3+Ceg972aO76ow/pB1pwzuyk7m6Nv76EHZhg
tJlAA6iZOgPg6GCkqZUsLVCbcUL/jqRl6htw+bbFHFT4fc2/RwZWNOfOERaUD7NksCdJ+v77s7ZA
qyvclPXl17761izvr0n/dGAaw37fVScNffPvplhvDDgwetvVKIw4U3bzJ3VVVarBDNh468yObcdg
gHKJUInekdo0OSky5iDdrgNKGFIh3MUARY0uLjnAv+ZJv/qv4xBrVWYrt9FSs5T7EHAPEHNjuSrR
rAJbNqBOGUk2EhNrsolqFjQl+utQuaCvHJfvDfB8lv0gt+lWIZobueOIxuPmFNO/Y1RXEzowI2D5
Wy9MzQS8kioGoILNWgrNWpNUY2Yxd3qJd7RGPZySM3TP22oR5/NHbIA9K7SZj1tZDbI3zkUb5RoR
w8Aithde5tycGM2w5t5pDHV4piEx1fR8Xo+HKZsrjySKJzPMwLChfZcmfsMKb+nn/GegRlbWs43c
w0b3G3v4QaDdCH2jMy0mdr/mNpno8/LesWn4CVL/e0E3GRObjkcISMOnlBeo6c6ITt7ps2Gs+z5t
teCofzo77EHjeGZ/bbiSKXQIP4PAlHy5m9waSsKqN6fcYatCl8HH9vy1rJuA2vpgIsBAk4pJDm8F
30QEwXMTOWiT9Jrxc2e1IIbxlqjjS+rhgJxZSjeorye8KBPJ3D9yb/ogHALLG/rJ2/k05fyGaoPr
0njlerMF2vuelvorIyKz/WXLy3XJ1kJiYzdSaQvnJBZDMFgkP1472w0SUtNxNFherABii4PoSUaV
GcVwLU+Hlm2mWJ8L6Hp0OV+TGs6qzyD3teR6qPqbIjC+wacz+6ZsKTdg/F0HOs6KpXf8E8nPUXcO
CIluW7CkKZ+QilHZgiI0RH1bWg6i5MiJyqAAJZQwXyKxSZ3O95enu8sS6Jf/fvtvRnUShUmsmhg3
DXKAfju+zHgjD2GxZi89qDnmnTsk9DG11a21s9iuaZzgk3CYZJwaO/txdSo2aMw0/mqfW++hq9At
tVUpIdR6tNx33dihU0hAw1lQoYgwgCOZHdkDiu/isknozzItRMogVsRvDuBy/cORud6Oc6UiFomh
+qtKftU1JEh6hBpbr9CWKFxIDyXPvE0Gab0oDLqzEJV/VbcMw75mVbSicbO/RQ5M9mzD7zjGBFHu
tslLNRI1p7oqE+G12/XSKdBNhIqiWIy3PFE1Q3afR4uJ4fe+jL/IB7x5b88Eh31UXw61GbAYKKcW
DGv74Rc0q65z85Wgvw3RaMBxcdYaum7EG4WO/PX2c8ehKt3i/GOCjSqhJofg703HbkPUDFiuJGbD
YDpbeEqejSC6HJ9YJIx6iY6kedX7eWj7CwOvhLV+zqJHZUZCdp6QrHGlxslKIDMgMB4es9Bxw4fY
jH1nqtIKNf9FOW9K1uAHzyCvKEL2k6kSM8I/L0wH06aCinP1RxW4mQQbl3NeKq7JP0fzQoa0/isa
UbHJZJQVQuVIJBjw3kcra3qOKLPeNGFetZUiEWsDj6PeY3CBvwtS6liHJ7x3p9znBY5qcCb6KFcA
OxxAuKo6dZvvqwQUwHNwotpXsi6OkvFGIERCbf9Y6tidGVriZDOKndfmot+dohLX/87ASdX0Q/Ew
+Ty1w7zeVtPKFEobIax2txIdZScGryZL73NxMVdAkPd+uyLgRRZr1i2H4kQZN8MdAUAMqx3eBsAx
blQM/umoAickRQMJsYtzyy2NxeoXi3WurmGDSN+YzJD+48iv0ORwteIrAQkLoePC2DM4VK33Kbp4
nv955G/MOouTkXgtDHT5vQaCZrC3OGKZnkSoUDm7yjc8Xf0cyXhIlMYTAMBF/UWBsKYkTLHIeHG7
Iylra1PuArA6q0wWYWr8HtJPsFh5QIeXKUmHIpn9zV3KKMDBwNW2KiL+Fh7GiF7mXcyBG/iav1WV
lEGWftue5JtxSUqxREZ5wzLk6yLnKu+jC6RZ6DQOnrjxpnN9dolnVDpmlg7A7gyrYHLSGq/DYq2Y
49fT+BxlEuvagOPkt6g2bzT6B8Aq9hKMuoBuY/ID8v0nZq59cBr88YT1qISuDOOkTWltEop1ckET
MLfQpy9EAEINvBCixGpJolIPa7tw3k6zKSZKN46sfvOUJt3QTkS2YAIr5+o9z7RTPJAeCTEmZqQC
8MCBH5/nGZE65um5QuXasRNvwfqBb1dkVkVZppy5mn8EVM9kFpsTBv9vlL+oVglrFB8Q/dX/MJR8
87Db/eHiKvZwyaeu13rZs7OFfP6Axap/AfFtlZ/1BwumZwFR/4MbPJihNiRGkmqHSX+70RgGwAqd
9p1Y8MDQRdD7HixcAvGIm3vTAJNhog7QZ2A+xqjzGKb4emOPbCcPN3JXW2AAxzmOwRR9CUGbCiG7
TkRKoAxIhduJocQgpgAMuMrgMay4yvL5jOmE3UEDF3XdLV11mgaas8yoWeV0Z/KSEPszvuO6SaDU
PeD4T2AxFuu1CZ3a/CZmpwl5JsTQZHckEU7nJQ17Cz2q6RYApT8XvXJ8HtMUC0qK0S+I5mfNxpKe
7HOb8oY5HaVIIusvYlskQ+avHvJLpJk68ni4SjtXUzHT+sH0F5/XE9rASVr4T3mJvtP+ETK5gbH1
ktdsktdTvpbNsvbu6my+hnnAq/bjQqYJ2FDrqTdmXh/iwaU6EVFRg8FRN8jUxghU9Gypcu5oiUwA
VrgO4nM0vpGM8v1PTd5Dk1+AsR0kAzueQq7/ljPEodZX1aR8cUuc7BqOGZ9EEArxBSn/rb1OxunC
JNvooZ1pNQ/ZAPWhGAVwdpnrjC2UzaEriwCwOvhuXyQrTrh1FrcrHHiXdoFHXuS/L0+WUaVxjZ4d
X0G1ut/YbsKuY0tnpCYg2IAmgHPMHKCsTAzXTJJoNG0aVSZaLSzw3F6fLEErOfuHqwq+BMYE39Gr
pHFpJ7zgjipE0Q5Mf8mfgrynrvVCa/dtznWty5/E3lmdrPLQpMxbfRyDdHai7MsBd0pzrDjqxJvX
aLReyhxTTiFVWF+5/uiAMwvZzxY0RdLSxkbzX2nIihC2wQ6Zqze9THsv7+uYLViR99BhZzBlXpsW
bO42LhtwCg8Kphl3mI+5S7Tq1BQmBW4wcUe6j0wTMKGkcfNWdQ1F2ipN9cMvW1IFVKGvIVo8Ujqq
3tOUB1zagtDu+sFvOU7UEzsv6uARd3MpXqj6cW5KAsV4OpUYmqYkfb9esUAmPWUwKt1KrFM/c4PN
N0mYIxhtaeTO1CzsUdomlkXZ8XsHjFgqS8qCQAaNNlfII/hMPcF2MXAhk58YDpprsM/S7B5doc5X
3SIJU08H0Y6TJpabXHf23Sd8vTFwYyYb0brn5y0pX+aU0rwnSL9z61R8Ls0nxzLkw6k6SYCLY0e7
dlTcvVRTInK7TAVYvSuXfa4lNfkg/J4HheXedGsmkZSKxo3LV6NZE/NzDzEDx2gufpFyK1hCaLVO
YaiZvpow3GsrRulAP0LlJuw0Ej6nJKnQE18Ml34OyfnidMF6tvTUv3bOtLPrRb9GvmBIXPVIF8f5
pQvNrtG8ipQHllb8jUVW4HkBKEY+jdbQ4Ao9KWwgXbIt3v2RoMtjOIwtv8XqMuVM58YWPszfuTgy
4OrFnNf7/cENh/3acHQuhkkRGKJsnTbZZ2AlhJZuwLrYUDVllDeJSPFbhNab78Doxfto3O+JFEXL
8Eg4h+oQrGa22/6jdtpgDxi5BWD9P0hDd5DvFJBCX3O6TKE+xy5vN1uXnXZIhIA6gx6vBZRVjZUq
xuZ2udW63ABpfWxHL6oQSEBlepFlORCTH+nwYQfP8wfAJYn+B2tz9BlvzyhOBILZhOgISLHNNJe2
gQIA5/mCXZbBzz7pl4DF0G6t7a2kjlwTJXppfVI0Ngq1urKUy+8cy9XwLbQ1e2kOkeAO5+HFcory
dcTiIcadlq0zNTPNUYxY+Ssl0sLZ/ivmzb9MKe59z/aZey13rr0RFEOAsmKUNHXLpMycDZxSX5Du
57QfzZubW+nF+SUsXeAOl2jH+/h509SctTEGyAqy4yXDJp+vDszquyrKQ7y9g65kT9YLp+8oKhBL
FMnZ8fz0kWN/t0Mvx2Wquek3cH2hnDLuMFrQEVIW6a6x7YssB/HZMzNPnE3qJdYnITdOqA3BefCq
6Eiy6bt2Zsl9cTFE1xdeoReuE7LgVKER4p/WwPA00joWrNTFAJQcWKWJss5vfYHhrvGuQW3+VWp+
z0bYlBbZVc7US3Xq5K0ZfXndpKWn7G74ZGCcBx7s0YAnCsIWZXyFNAX3/42sOmRW983dv9rntUcT
emyhGy3gGH8A9kdDBMHUB5KY3Ys+EcUgjcssWDAgKNmn3Siv5+o/Hsj20n5PNK02qqdIX181FP9h
WTOJKmup6qspRTaxlazejxNvCXKvfnerCjMqUkekQuuMvVMJJbrbVMef21PqLqKv6PkoAxi3DtTM
fri0N052gOqa6FGrTCLbtgPzc/n73UQmxC1J0UyNkoE/VczBB/L2zEEGVs4NemLfE5HvD5bepwhV
uHAn0s19UI6mVHJT7aeDZRJpzauxYscBkddMKd/FHn9nzwP8rJeTaHgmp7GKW+SMLoAhtqRIOXNL
+TRf7VtpD1fXVgLvYCWwJ5Jx3KK9gL5FYVjdBkMUiCYFyheFDvRhMr/euxy7/15zoJSmz2WYUgtw
AXd3EWnoVAIWPz76pVvEfPBR5bhVp1KMpNzrLxZ/Z0vPsUyCmIb9gdYwOtq7arEgUOjZIXxvFihi
ajR3wpeb3V5AGlR816TojnvmhmjabWu7CnSsyC9+WC7oWtrjJMtu7U3F77GhuG9Ytm/JFZcxR5iV
+rjWbABAjGbHYbCOAM9sOrnr3ZbaPUA/fQ0v1IMcERAJ1H5iM//ujYRwmcAbpdmot6U2OoYwKbqa
4tWPQsExtypB/lGvbPsMuaOujenOefRoo8WuIQDciTYZi1/SgnPpVVE9nsRZpHOsJOUeWaUav8Vh
3Vr7HMJRhOOt4+vxnly0nfoe3MEMz++TO9cBzxpAaSO/MO8UX+uqj6SlH92KVYAlJ/+uDtUmYafB
GGNUrDw9vB6Y7IFW9ST4o/S4+mj13NIY0l2gbVbPk50omlUyvfJn4bCY/k435xPVWHGuKiCeVm9N
q1oQsRZ9KR4u/6NITQTs5PtuvVoUpktPg71+JIZC+L3Yq+R7bDeyW/cpGT3LlU19lGU+TLNUeByR
ltqXV7icBcpUDHn9uBBgEm9V0OcGKLIMi5LnWS1egLNb9Lq4EEttCQhHhUvzKvPZzIfylmm2USGu
9zFNp770j/ke/F3jBF5CXdp3jI6xNiRfy13ZnUskZPXzXXZ6Tae+SqyzgmraBKB3y7GGWlKG6dMn
pz5YkefQ2I9uzTB/Y4jjbSeu3Wb7XY0aUhyceJ09yulUEX9ZCc5Sk3gFKOm2ukrY2OQjsPGHifVf
UEyx5C8EBkJW2SopJNaCtJXpRBnJ1pfHi+0ADQs46xfSTNGWxDx1lxfAERUfGuIokC0ypVDSi5mU
OdKzpitaXRRVz9myhbbNzsW30zNYGGfkDnOePrzhG7JSEzwD/AEsLOm6kVH46EarmhGTg2Zz0spy
gQBVS5ANM802jSKEZtnXsw91bKTNsd3900JaCifIJO1DnEXPa2jP/fBmnfw8tdwnkaBVlZ4RogtU
cHFmDTVfDjdL5D0MYbGmIBP8yNaw4xEVXGuznIgN+3yDwYt22LPEsF7C47v37XGXfKErbfGzccxS
IfRoYndcJdLWFzuSYKDhIeBjEADr6X0OiL3Z3+yo9cbVHC0NVO2uzWavek5iua7wMCTJsxcpN5QI
8uVknbh5oCSVWbOEkwhLU0glMjD9yC45fb1iIeiWTyKAGXkSbjX2Ij37zQqRM+acl8U7ETg2zcAp
0KbUa9owkwIIFXrRatMJ5PaFeXA9FFmnMk9sWpQQIr9kT+fGjKrVaduWRoRS+1WNG0SxOIDz+vr7
4lJoTBMZwid4V4Rn847G/lm372AbeThMgXL3AkdMsRpu0kdc28Bq3nkr4W6BjfZmfVS59i68d2AB
UzmPz/tAw4nnouqWEkwH6u4gJdjkBIMeUcg3D5GC1XyVfd4xH+qDQsxH/rfgGGLgZ0Sub4QT6ewc
Y7KF+8MR6ob54VkG8O6gUjQ0ywZahi6TQf4fjG+p9Ah946mPKLh8SVwmcPeCDNyRF4mnHI3LSPj2
EIkpxkwcIOmAzVT2bCDmWuiyiTrZyAJfwJHVHi1ieRezgHcK18UNjvdEIxaSihR47T8WkPaK+4lL
r/DclhBFxvrCq8FMTLdtVsGBX8USdLpRxq13IzIIIZey2ZZuXrrkOpdEF/Z2o73cXIkwoj2aYdzH
hTyUIMaUY3RdY61ALNlnKIOKw7fM924uGki/SK9Pz1Re1HV17l9ssfvM2+pYtIgK81SrJtUsGBR/
tqj2/9W1fozjcYN1a9oqjib6ZyaQ4e6trIeSRHIFoly9IK+rbjx/StPbpph1nlkrVRzdOzZxlbrn
7tOuHHLN3lGYcU2iNkoSwvlUd78j62Wb4XjgxHEHjGnUOyaB8knOooh+bUD7xDpD5jeVIRdRMEkC
7Z5PenVdzUODUHPlC1bZVhhf5+lgsM7GZn8w6kbj3rAveRz1ybvFUDP/H2kb7fQBYmuBhQIHjxDn
NdN+efctF/OuMzhpaT0Yrkh80SUGPU8jDxZlZrPuFDsXFo1uXJT7hLNNplCRtttrnwPpczvYYjhr
A2GLMbc2kUDsgqFKgOFntGzkMyaOUPhrZhrhaIn3m7LNGrnB7H6w9mWazgZYgDr/rycaz8TFxtC6
zNGNG3bWqzAl5YicrQIspszeOIWtGMUCnYm1pufdsR3JW4SrO9e/RJwvihQMqGnWS6QTgNPygOsW
Y07OMs2YmVT/Yel7DU0G7Qwy2cJusup5mzRcJZgKsP9MJlApS09xE2+itSyHR/2VcImFLb/fcIdi
lyd6aTUY9ONGt0xXAIcIdCUjLUF8lTjxS7bsdVQxOHrf2a9gz7UH7d/PVdvkFYPOpYcyhOlfMFWG
6XFftapqel/iEwdgX9QyozkYwwUbo7WN/6v63/hh4j6hVuEmpajmFeJ9SdezzHuLUlndNwFALDY3
beyLnb8hJh43gP9yXWBPMHCU/3pUmDSo68EKBGUYGTmFKatopnPjJ6bV1Dytn9jEaj4lO9VJixr1
47cBh662bGxv5PLjkKkmCM3vq6JjKBT4sm4qm3o325Ad4ydyxHdnTzNgdTC6/7/Q8MObT218/6vK
3sL7spZmEzKolw8j71CCHKXW3ynW9ssKDUmZHnAYS4EaYOKaXQgHh4nfd9nH2ggm23/0RlVmYhzs
rueQxz9kqmIqwO1Z1M24iCYghffBC1yGfr+tEOyIT4jX7rDHVKT3GvfqweWdzcrB2lPbSHvAHyfU
PPoT1j0X0NX73LnRr5skQjgHbFMFLLESpgyoyLJmOrgWbaQpPaAc7nZYoSbtGGWnioRmXSV6v08d
fp1AGLNOcEmKQvrVgX1XAAIeUr/nuikSE5XAtYgQrOSwkae5KqLC72yVA+p1TRZjKjr1p6Ihg5AW
ZczJcONrVRdLlFUEVlcrAJAwUy7nCLzOGBGTJg6KEbn+TrUpyyknHqDCKww8haCVRabHX7bUnBe7
fLovlwdPlP6ezal3Mzz1u1f0ebfgrArB0FEzYjoswAzEPK9eiSSgUHPu+jlKgOHOgXEqHFjbCXOn
MRhh1ZIHS9BdL329RuRo6wnVWpGaVnvCzSi9H/dHLT8LVJX8mdw3BX+n6l8EYFUrbkmuLWyRnkcQ
fuXrQPKqqZiThRkgU7oKwvpMlqrb8l9vU00xAzN4jbV6bU3DB5eTb/LKlrZFxkrrht9qvFHs9VT5
C74zKGD/VhQ9JIXCLnE97rMi1aN2PnwebEdRWW8SPX1uiDIhjV0+fmNYg7Qr2bRvX7MCJyO2Dm0g
OHp+MtRZncsWJ1z1VecWxmCZvbftopREZWyRiwXmU2vtsFNcWTgwnK2ASNslpnpmJm99T5Z0t5T9
YrV0YzlGGzgQSaQ5p+pnI/vp35vetKn2cnr5w+zk9mJaXDsLpZEnWXJgS2xPpvkveHO2c70hHPmj
nU7wPivWh/jqEHEhwTC72M2B0qNkeK2MZuK0dPAHtmBSEJUumPkDAry+4xU5RmPP+4I9TDwSpOun
fAaO6njFK41DZ9W51+1zYHkjff579SuT29eBSYkCYNw/JTcTbOlzzk82kZWOuo3y/cmjlp5zofRf
QaiuEO2u+ASvAo2c/70LS4t0e51M5mo2XFGmBu0PG0TBOhSCPxJ7K1qtJOc0nVxcB6e7fxp1Ubf+
V8hBIOqnCWe/byw+YAqBCdJSS4G29nyDgcOHsUnKIOgALrxva5N4wMnw3HZa25HUHgOLMzVUa94R
nHdHuoUoJ1G+XKom5C1sZeWGPmGRHL/7ye1MHbY+sIkqTVvkxjnN7o8zW/nq0MEqr5WsQKn8N7C8
jGssF7sF3G0M0LqtMsBNrSOOQTRntlTcFn1Lrw22wd7TIJU30Sw+g6emLzfOTIG7bdkkpFI2Ne2D
Pbvmv9kystjwhhQSpEVdXyu94tkrZWR4Gt+3uSxzoa2GD3V7Zm4y3Yf4kByh3wFszTfTZJx6Tf/M
O/DSWpe7RKUAmmlEjdTurGvIB0VnU+yq5tsC4QHq/9y7IAinS2Gi1ScpCdk0+joa7ncrysvSHHpt
qBc59NZ+nV2WSAmzumLRkXRRfwbsS2WRPiEPtYU7SQkbt1LW5GtBpskCt6pWWhkFo9F1kRuL2uc/
TeuSSLQkT2cicHlD0iPl3vIA5yqCM/EcxlDd74WoMBa0KPTTNqtghS+8USK9grh38tTR5ksLF7Ld
pzErLSKiFwuUOpoK0kqTtYZ5UQCtvr4QcqywlZ4mhMRx41lurk/3GRRgMtl51JMHyvbtg7wlxnXk
1Vm3dku2ATgHcNz94ccfF5n0Jk5fqZrxXK/BJAgJqDWf4TpWoMO23bmY17yztFeEk+HzwuIPUb+d
4Z8sZxfd600c8sAyNw3Ifp6+5WA/xxP8AzIaVqa4fvHT/rdoMUn+m/MKgq6iF44daYXkER8lGx1T
WCOWa9RhCGSK5mMmTS0JnhaeG0PuhuGrJaY0r666N0DGlF8Gf39y6T6HiFhZL/SdbXeCKoxHGW34
otpwPaNll5r32TvnTdGjCjDioHA0yFXd495syctIs0tyJqcN4Rc5oR2HahFxV5wmcig4qOnxucTi
Qc7dCY9/Ey6cSGYeWdmJaCPwJQMpSJtDkwEtbcEc33VluLURFjEcul1cm2yidc4CSwAH0wbugV7k
XO39kbQVfloQ8gpelZ507TH8EaADhdg05R/rM1XdHxjVV3pHcDxvVL7ntXD4VVo5Kxe3Z1zP1HEn
C983pSNIM4VilWWXHYfmF4ZgZpZB5UKNV29wd4sLn1s0iitVNpwY51d43qyI7MSG+i1AxpTHEqOS
/wC0MNIIl3RHcB5KhjSR7n2VZdX2BGX3cri76xqp8WoCF0pa6koUBYno1ISXaLTH0j+Iw+Y8d9aT
x3BEPM8JEKRBF90aggg7+sxvQEEzqDQATB+hXUp3FhO5/ElNVMC0a9XqDQ+E06kT5lGvFTQsI7+n
bRk3DdwRUJF4Y9nAfDOvC7FeeHLcQ/hxbNVmaougRPr1GgTTWKFNOd01ooooP3DrKLSHh2nLRhi0
vRW6pAw4r7/NB58qYk3PUy0/XcmADv/urmbSHQrmvAqraGIlPxYfkWb8liop0Q4fP2Y75uKezZx3
fzh3IotmmaT89I2aFbs+BLeWtkvd7UGaQbfzUmeKRu6EcR8mBhZRFGpKy/mSjDgXg7gBc2bR+M6j
QcrVWu3gm3RcLfAp+L1J8kdN2J1lacm4SflkQ726EhAK2bYQF3z7zH1RSFUIrs2MWxE3JT0MCwsF
7BZT5XaH8abTCE8oD6dMZ4TtUiZskD+2s5xbwjVDM6ZBy7dQp4iz0x/8mNx+SG+Im9kDDXqoTzTd
Ttgio2iipGDGRkyWG0I0NXEik/8y65IsLLPXbtuN8X6/o8bQy7ZgUC5cJzLa/qAGy6+POU29V4f3
XAMNshUQdDTCQicRmZhQ224vmyEqvoqeRs1nNHbJYfpeQbrfxS5NRbU85Kdy2cLOWQdP51Tv05ey
djRPRKv6QFCj944lw0OTiGYX78RVPHNkFhQruLLCWvNoERk4YZQqHhKNv7DRyR7ITdlURPq5WIYo
rsB2gQYdVeQutfwlhr1J/Rq+hGVV6NGxoHDs4bbA+UvehvOTPpKEkqFDnUfGRG7lSD762rtjdCA4
dyFGrxRSM7KagmKfyzpNDujCEmWvUI9U9hasNNQvLymdGK8ktVM/29NdBsMpAxFtKea0CUw43+0v
YKOPxr+1H4C61c77VPVxORFW6jDmSBVEZwcpQURqW6oapkQhmga/fSPwLY2YJvj5CqMZeyLEFD9j
KumtwGqZW0FT+Y3kDd9ig2nJkICVRGsMqZpJdQ1a2ZNQhVEC5QZ53Tx1BZHvJVNZeBYMifaYvuBR
/apVmYumDo0U95n7C2G0PxL5vYU0Tqe4IG1Xs/Us/ADuTBcog7LV9GoDuqRMoNTaM3kstpyyT4d9
BqscJ2EjpXGjSY1z3CqY0VCcyrxkAIaGHD5jaRq8J3pvWMooclhJ14Ev1YN7YOz1u9O9aaRwKk/i
wiZumxvMZbPBCjk9xC384TRh1v7H1V5ZVLNoETyVd0MGr3tZCyW0QTLHAgmPthKmkzdTTCiRGH4z
lPHLWgipU0ETP7wiLUOI3q0w2mJ2WtuZDsC8F3l3zXsMO2m5puxK3ziUo19MtjmVsiSiSXBgZVDF
6P1fOeWaMmlSzEns2aeUOVl1va8ipM8x5tqugHNz10vit07v0OcIaxvhdmC0biOmw1pSSyo+5Uk5
ZlLmbg9gd6MktfncKKglahQHkuKJbFITkPrzH34ohknh5sDUz3QxfHg913sU+dXiIJRBp6wSc/pK
T37rZxqB0iOZq/uvA/bI2gs44TQ1LI/FgaclIu91gpvEceXtzdI1FB4JwyNan9fgVF84Zk71IRNr
oHs8f4Z13SjTQkGLkwqAWzDpEdwVyq7HmVxD8z2+s5PDkphGjfCWMvN5hMn/8I/NWzjQtK71giU6
q/IX7cG0HUuozyK1ZiLMalZsm0+erg9aDxZ45Ry0jmyu3KPLxD6sJNdkXbYvDVWIxoItbgbR4m5a
qaoV0vZXtugaShzfWREZG6gJEbvmZC2RnSbM9fAsnhQtLx+9CliToQC7aRI2aaS6hxmHy3AZ3nne
DwuqyHAYrSKbzyHrrfnK4pVw4JAkbs+nlIHyWeJIxj6vJqgLue/qR+9td3JVtlGryo3LcCUQh6N5
GB8B/vyNaOJNjyfmorvMNRkJhBNewT0DZTTx2OZ0BWOf1fugMPV+dfItrUIA+RH/l2fc8FXPj/FP
TxTSZ2lTFnytafNX2hoYJhBCAh/cA5b2n/yi3grSpY4aq9ySOEQ25Lq4Ki+g1sc+/tZyfOJK7xAU
5U8cpVRJwa/nyrdbMldByjq9nRDbiOoDiOMMQMMmC/pEnsDUyVUQ61JRhXqF8q3RbgnHkCC56Not
XSFrGSpSqot8DeL7ZTHw4Xw5gq8FKGtLsJBpteNj0uuVC3RMKJz4lKID48Ps7qHD7GTRDdJ7sfAL
XFg+jeXp12fBFFw6Us9Ct65FgzyECbtP53EdmHyLKj6/Ss5K2DiUQEVYriFL2kPg/g690RS3PU0V
ZpE7PU8JRHjXf3zj3exndZ2PaoO8Fxghy4svtVvUhEzlOHh4aOIz7J2vQsvIfHH3HCL1wxIq41PQ
/Jh4PmgixaMhD2rOa+5ENifVUewHJmLs6fzu78oei4FUPENCa5YLyOohZk26X6/eUd+dCFQmCn5U
4U9fVtquXYtEkbDbNlMdAeCyq72zr7qoyjhjuRHJmNPRYwMXUhbX3nO7obss7Z7RTM8XE7RO82lv
W8mEuQu4hiSKe1VYpOWNvHCHoQkXVZHBf4gQziryy+g4BXSAvk13QyKHLFvo1BH1r2CFDYFecIqr
V/F2GzPs76bZeWE0TFHgmq43YduWNI+bOhYAU9l8c17mU4QjMbqFycaQRC2zvJ7iUEc2X20+9siE
f18Kz17Lpy6ZAEX72zPQbh/OiB9oMerF3bJ803nYceD4f3VZIuc110cMJuTbfniWfT/X0EjNdMkm
l0BKvg30u46EAX9T/oWTIaCHQpWLhZH+yjiONcjZFngXLdiJd/z9YXcktYQt9B2Jv4Ko1mpE/SFG
vqkLbwjIKbWt3xh3jiC93LuxeiuzzY27ir5u8YwYQC4v/hDu5vQ7DxuodtymyblK8LKxW7tdFDWt
CPa9wicReTumgU3Es+ezeW84+R+i4zEl3TM5WcFaIBumg2czenW3541CKuC231k5QLJD79tum3bH
diPcmZuPokMdAM0fIAhEmv4/StOO14UWLLmQ8b8n2j5dQ/OfbRJNIzRB+vGRxCGqAdO4bwNyYrdX
srnPDVPjYq4T0QAJkfAIGTGd/qVHpbRbsY0PZ6bZc+gy1OdaQG3zuZ3FhxWy+250dId+M/pe83C4
N7n1ArmWpW1gzumWmJ6ETBt4RBDrJ7gITgP5zzcP0aLPHizVi5O76QD9NeW00dUvcP8/zNf6zUOf
v9+Ss2ATBe9Bd2/gmlbYlumJVXajWb601cLm5PuXpNKwIRYD6mR29TzeQcnL9FC/sJGsriDKA8Ja
MVaCmX3zfWKajzFPLYAEkA7/cvS5c9pF0Y1z83dgOJOBrVztVC9CdF5vnvqrIIZqCsxbddVZcUKe
XMQ+hfJsZO6rwhqgwHxGQBQ5xFPBdAh4zDP2B2C61sb0fbX7J1KqAvI6MtcR0yOhUsLjq/tRH1KR
p4N3p1n77k6LOB7pVlw00vj2OIV56fQ6zpDEF5Uw4Bj6znUPCEnModCEHYhpniZL6i1Yxv4+Hz0s
hqB0xaYYpG1PmDDbqBOF5IbtO/fVaxCw33O4OSmL34SrtmRbdEVfTC00i9p/czw3o46YaSAYXmzb
Qg7kW4QIy2cbp64SUdn1OwSg2j5NAtefpAZcvkLag79aOoyyjoqtPaa8ciMwa3r16/iXgPalx0Mt
iaz7bZqqrevuu4N5GYqItDhKJ4wXcLvgjfx17z0zJ9vsWNlgqzhJd58BHibnX3YxdGqhbkIGs1b0
U+0Ne+B4gZT1ti5V/r0FeI4PLz8OOCH6HoLgGiJKIkh0npr07n3wriAaa7brK/ZFwDz3kVVxw3x8
KlszlOBQ8d9qpvWDGy98t/Ig1Hs3wE1Vn9jH38cdOXvtyhpAw7yBQeQZsdYud+XM7jCdO5MgSNDM
59NttIAC9E9XMEMvdMe9TXzjwjw7uMfp7YHiUkSuDA9aFM7PnNoTLyc/Eu2e/DI96KT3dgSPC54B
U2qsWwmWgvaEyKBEyT6s/s54T3nxIDIcxa219Vkn8EdoI0K7AqZTmdyYCpDs/N4BjfxmcUWyf/PO
R0181CTLBlOYg2rttT/txekL9c8vZY45csdLqAzl1bh6HCeu8WGa2gILTLtxiVujT4Gw3FZhqpBQ
8gBNnDsGWAmBi6Wq1StazWJ4T1Zsdi7f6UQC64s2ihUkgJ8gXXwT1RC47PTOPaRKlRINc+osy6Tg
HpROgnRsLHW0ADzqN3XmnceuOiRcLEk0xYuzARQUOdXZifzX6dg4RtxyjtCuT7P7S6A81fgtZxXs
EIjX7UbrTq6wrniX38yLLSypoQEthZWw2lKzIDRNLWTL2NgohkidpWXRm593BJ1G0xS8fRpzfpmx
74ZWH8kKCBR+0bLrjfQwCj1BhSO40BcsbvNlbeJ97hlhnqD6jIYm37PuDWl4A1ylJt+XYRFwrc7U
nKO/XQjgkoqnf5ZG6U045XrZE8GL/T7te494WrZiYTN9+Seh8NjD0qcZvq6RUNkxT8fUGohyEWGi
Sce3g7WyknEKCdVXumneegwCkDmCv86X5AXoJTaIo/8DfCyiKEl+O2NyvObfXqK6JhhADfZUurY2
1AkTqroy2qWEB4tkQW2rqiz2s7R3M3pWEz/N+ueSIrquUd4zJ4M8EQTR9Uxom1jdwr8q3vBl8oVM
PurqYufRv9gYmgm0Red6G1Tzu21b8HoEPd5eWrYB6ctKyZEjls1LnyP0b9pa6BY0+ompQPeSLboI
FxvHW/V2Lo9Wqm3crlMJV2F0tGtbgAhowu8m+KMUmMSjNwwyDY/Beotq+QjBWzoK5cyjnX/rVL23
hH6hLJXLmOcFiXeo1E9dKNdy2ivq3Fp2fCEQEX8w7BtiAL2y4aPJFwaIzZxPtPvoIQ3ged4CC0tz
kN2z1b41Py3DJ0PzscvfcZUpkqZ0rTLAAr2aBV4KT5p82T4/HJznc+elLpZz0iz2hHRLHU9R++Fs
jf8nE+n07Ah7TGdrmf7P6BViJh2J92YbobFBaZkZQbnaPdHOseEIKIc/BiIotbsJ1jJ5xXOI5WU6
nZQGGjSTCwULExCNo8mu5xH00CHXzuzfimCrGa7fcb3WBeNq2d7s8jsY4q6nRvqLmRH2625KSn2w
omYVx6xWjGOY858Z/Si9EEJ+dIaJyxykSIlEQFCFWe4nIZ/Y75mSIgu2tCYWQYb83uIX7YxGQSbB
QPZk8Opl5JK6ayTiX+G39OOykNN/jraoV/0Gp0fDA+BxJntV5IVFOmya5GAfzMFQzbeWtTkGLXy/
IToTLGdwt4y2W9lopGxqDyCn0IZX/fP5yaYgDv5czhz2q2WVS8qx/49d/hY09z88X84QFsf7fSsz
LLiD7Dr0HxBMVLF0REgcUeffniFdji20vpT/2zzfoIgHi/8KdwFJsFMqRc8Ton5TRrp7Baf5BbSg
n+0Tkam0cE9igF9Uslpq/2XnoW14rcDQhrxdwY0vBDfQhmdUPAy9DY7CZiQbgKKMsiBbo+29qqnh
WSD6t9kKHg+yzE3xab8niYtXTFk0Ioub1M8km3SsBU/kty0B0zObCCSTEZ/JMZem9fYswVIqu2p6
md5mma829zF+CTNgPj/Y8s63Lyq7Yt7wh+kED7HsMZqP44I0PhVa7BL9nq3feicAduzFOIl1px7p
6A3bSIwelpCBCFprE9vbepsf6Uq1Mc56idMIziV2+K15Qvc7OIy7fGFCRhrQXwHGAByiHZErfEbl
BXJqoNPwYPRblq1tA+HT20Vt8YdLT0nZPhhVbZFMjKPtBrPi9D0ahSIcoQbAp2v2veIZu70uD6Xl
EDek6pfmYeHna99m7sUyN8gf/HbMNrVGRlF8l8oiV1bJHzXzgIDIIR/VcEjJrhbVMlAzLugNsv/N
QiaoYQ38AKBGUvebfBxIAta8cGtG47fBSULrqb86hqpiD2Vsac6XR+qDIFkhgu9iq8amT57MTioD
99t+Dd5kRpM6bHgZqilJTFuE+oFnJ/9sv3i6G869/mT/SJYti9XSAWupd8P3hoe1OaNzxfh+WnHl
HrDTr/JXyvEaqev7H4KiygKW9+yguhDKk38g7EvDsXIoR/VMDNtULMzBmxitXf4GQveBg5xG6DKB
1E6G0X4vwAjpV2GP3dXSo8soREGyhbZ86FtdPQz6UfOgBrA5lRLUbrNUBKlEzPHe9wqLKaRzzqN5
VH3wTxOErmvnrtYXVZTIyv3Z46pIg93kgl+HYOFH0xJcrvjxI1TVCMsVzcZajfGgbdi+4un/+Hvi
OIbETrgGw8CYpFGVTch0NJmcHz7o2J1bNtM6HJ3y2mYnKLH68Hxy5PAmzU7OeUUtlyA51Po84Jdb
YqS8nxobax+ZJETwo2BxCe/z62NKCwMmHPSGW5ZJ1M5hAjLhVP1Df41rMuJEjksMipC9ISQ8oP2N
mCOxXxFCFqsYAlvHkKtpmlOVBwt9CoPJubNoOfF9CY7ksedobMqPM+p2wkR8NWVXc6XoV0QErrv3
xnR+Ghk9rKKL3HK6udf5n8z/uo11x2zCJLNSg6Cgyk+2XwwEfEeShrA5rs4xf9O34B0NwCdHEnMi
Y0rseWIDjO6Cuph9ILEY+VepIq7v8rFM2e7L/OLL2FkQSvOQXx939FjZj5aZcNPVAcrcT5Bl3u9+
DsrT04rP3TYbB06UN8n8rZAT+spAdIwSx+sPuEN02FXRRbQ51bZeAiDaRVE2DHmg03l53GUpS94N
4reh5ZMdsU6qU0kU9jzEuFjcNPM5NzBL62MJ5R+4qAn/6wrCIt2YHf1w8mkoXb3dgtHk6UOPpZkF
aRMjn9Y0fbIcH4cEPVNOKGuuYLaVaceJAejsnW7yYVx1k2RP6tMhXvGdUN9qyR6BLpc/zPeIvZPH
3k+yzTC2jHQ09AHpqqsmf787rIZtslo75bP/FzwbzGcb/Es4zgNMgoDTYRGRPaD94UFlcn6bya9K
wL2AC+tkfco6/P3JdCj9KgnYajorTa7XbhtCRgTDEzd3vsWE1D0/iwbcB2szYfPzFCz0ywtIjH2d
j6VppsyQVfttjvDjN1UPmR87ORK5lHIiyh7i9a8bK3u/oGQiZ+vrOl6HMK03cM0tboXishjg0mE0
pQs4cJcolkUlfbtLBUclJg7V4aBlRmf7EY3gOF19ydAZUDZx19vm6sPAZ+3oLnZKI9qmk8ibUWi4
H9/yl7tvFBw4MYLJCEMTW/SBRf+TsPL/MIsjC8dSn5cQC0mFlG56DhEeSLs0vi4zciRugZxO0PWb
mKnpG+QWGxz9nR7pIBMMQt2W+YcRDKWDyAH4Mh4GPKTbB8hezBFPfr2gLSnNGevuNrkfzWnBlNkr
wG8aM9eR2R1P8FIOvTeUvtY/h3MaZMTwWjIooBd+2y2af0n9JmRv4lmy5UVofab2gfuIIlgAi6L4
lsAMDqBideItwapaDfkhDAahZu7XmCuvZNQ2Sxf3uwcV3LtTEU/TThLe90iPCXyrVzlhzZn6BGDX
UAb3FELMggqxWU1AA6GvUV7yfSc0AAjWWn1n8iBBbE1CqihN/bs5vH3sLRpqfKWXU3Z8aCbylqLp
Oq/ND2Of6E5KsDztJIJy0DDvSaB4ziuzOxgDE0fpLSrJN4ob/UBFiScoFEczcP3/D/FS7UYkC5/B
fhAFHGVXSzjJVIk0d1qfDien0J0FG3DvDAivaOasKBw4nPH3iy59fpMXR0+S2o7gYPRNR+L+AHkE
b7OnKLP/kFw+pThhhApWDMIEt04fqBMpzeJ+oIpFzRPr4RzC/QSYSBffJ5Y6bQ5vkhDeYZLD14gG
I+NcSrzaeZ/DKok72rTsAQlhSCwxkMVFWnZXDc3muEMWxt6a98dZpgznR3f4QDxN9zaUNXvyAGnS
reYrpE+2Gidg8f/AkpQSZ5a4nsreXBail7TYtzlkXEvids2nXQ3iVlz5CXESyxE7MIj4r0QxuFKK
Gcz1fWuKJFVIchME/C320w9YhKiwXOp5fuq7/T+b21UpoHKGgUBMf25L41uOURxXCNbfcH2StP+p
KarbbVJtvFkuyrirqA4XPS0ETCm55dMwZU0ThlMMDKLYFEyuhTdKJMMVnFlKe+5TqLddT+KVkuxO
kHoHdCwnd9+6/T4UB+I/IsKWYBzPqM7CPvlwW7m0RVovfyGVuabMemYd3jhPN2qV85nNU8ATQO+y
ceDGngnyl2ZhXfR3O+ZuG8y8RXbeLjQ4UmYH80DQbm6nTGjKtB/bqdLrfu8o3nVRlZEc+PVqeiXZ
jb+gUs5ZIuNcLdBvEU3U1S0pSD9e2ib8sM4CCxtvzgQlaC4tPCnpFWx1yYwVntHZrIAbQ1UUDfkT
CsZ9Q2XrBrL36Y8WRd5M8PUECfB7G+uq/YjCfkf9q1AmszG6fFFSKF1ePC5mY+LDtUjLKH5ZuoSK
aMcEN/Ju3dkJHXGBKRpNdDqOHens1CEC8Bi86HKZExaRgV3wHkvyFCy7/yFePBhU5AIBPPYRTGvx
vQH5TNFV2LGB2WxA3vh5v+Na85dPpJ3GY1O5HgLSXVrXNiB4bnnsPcJ45U+/hvPs3L5bYpu0Y2s4
Kcu1I8zCQIbeWUkAcE073xdU0oBIPtaAoe7n2FaThKctjT+RsVvKDE+YhS7DvyZz06mEJ9+n7Iie
XAWCo1JHZFycxXJQpnXOdeWHGxRBaGaMlPJ+0aOj+bfMAtEnkaa8DR8Ousa/BNBzRqJdiC0I9zih
O11uC4Eow0m69MMjxIWHx6zP42exGkGC+uxARHfS/NvTp6PH6ZjgrBgwDhmSdgLcU3K5iOiEzC/T
uQwA50gc/NvMo7XtsepUd0UIFvpVZrP5/kR9oWdLH5hpB0dphqerd5onw0Mb2CYh69OtEOQukMF1
J52WJMAv+Ohi0ALv1bfOFygOI8hV6WRsHB798po2rHc6zMM7bUaD5SjjHnwP7LZiSOfVZaYtmzX3
QO+Ol9/Ir8JlIpkvbf+q/serNB6/dSuXaqBTQVxUnJ5p3VVFEbM9SJ39j9Eag0SEdTGvh+35dE3A
FNmxdcXoilyyISmo+Vc6+urymO0hELKXm6p+4nlyNdsHOvU6bTPvksBenNfBU/g4UimAqVxj20mm
z13dzWF94uGktn3kJXDQJOxXQm7kodz35DTu1f55gACqu8GjTn+OyoT2qVYf7WJMzjhkCLh3NBv8
DrWjZZhx+6wX38YlEKxou5WD72PZ4lj5MvCcDME0xmeMhk+e7E0UcPAVqXbNagDiopfVh9a437m4
ZdL7ZTtX57B/a3yo1u1t8doRVQm3Lj0+OdHO8eXvg9VPXSJJWu3wDYD6HFs6oVFUlnWs3mza0I/Q
X+78CPsoJWG65UonD09EpFxf1CVxLaqOZEv4tQC6V3YtF00vm0XCig54hQe83jrdB46mXfX/yOdE
dOrPp5Py+GP2BXhRqdr/t0h4Y+avn+XJFw5lPwuhjU29Yn51zju8yrjKkLXwuzovQm03/FcfnGwE
LR3f0qC9X7TJei6VIt4BEXU+HJ0Sq7kU6c2LZ00KVUpedjId9i6MqWP+Li9e7QpaSNSczMmSTQjP
93dix87YyUcCvmXxGNIkoMC6m1ij91N+mH7qJDggiL0jE79i2iXak4zQYF5pns7j7Y6nLJeXFkwS
tqegeFViIVt5cv31RYc6ZqgBbZ9wHx6dNVM7rz3VYBPlFo5LRW27KHiIxTtO+bysAm+9tWAk+BlA
9YslQu7/KMFXwGqxjOPOsEAqsSg7U12aFkQQ0RepEjmNEmoXcTY9onk1G0tCZ+H8DNJcESX6SJU3
L9X9LJ97QLGOb1YmLVHWase2HMJYXUa/c9sYdoFvvACEipfJwkn/JW+D3wzOpkZzTAJTXgkW9BZZ
hl34kRtno6/BEcpSiQXD4EmhHm9Z9wl9F7zsEJWdXI07HLXEc83gGees4D+E/Myfd9Y3Kfuf59X6
dkfuyuDw+70+ejm9/6B6N8+w9rCp+t0mCHSIyyid2RIv6SD+VedYzXgFKeI+mZSCM7R7yz/b8V1z
zikmgjij8yVEYiUjQso4/RxZaHqiLwahClBKGgABXvgvjN7dodPTg3ZJ820bnL7dSuLTOYSNTFvM
mbZbCClnvzON8Fk5VGXGNKCVVU3AWMPpB87lTpOl3B73IhNz3Sd1Mw0iJqZr43h9DeckcWN8qN2x
7ElJn/+QPzHtV1JbTK72vYx9G/0G8Z6JB7zPnFwhLwDez+bYJwKg0y/IyRVq5IjIOrU8665vGNwO
lNMroDJ/h4XJtwEMZ7bGowsCc5De5NIFoqu8qt5FBJkS2p/bRGdvmnyfr0X24O3wPyIgWWvngvgv
Pd7Xpv8DxsqViTswJqdAGGzShCsz3T76fscuau6mIV2dZt2AeuOzlNVhvX1+z7xARI1DfREwvbce
oxtB4D7UdsGbZJ6d2DSDvDnEfJu6HHY137VopNYbQGwqZ1FwgqByj3xphRbMTONGtiMusLxasr+i
U1A6PxNhgR/LGa/7oid5AA2wxv6Cn2o3DT56p0rQ6XDHbrVWW/B1hWN7aLEFRsDxgM7nxjg+v3wC
dDJLvuL/h/DAjdSQjgnKFmSrbFE7Acap+u0k+xK8p0qv8yNzdnBUzJsKCWNv2FjGEpFGHvse9J/5
2zf9ZwgqXePlFbQrF1m+Wv54uwJ0/NWHIMDw7r5gRloqFriJ55uFRcmCf8fUzKSeI73lOo04GM+s
N6YaxlYYX5yENil6j2LCtVimpsBh215PMbCkRn09slSaAqBhjCPTlYT/3OiLFCTdmJu3fOcznhDl
Tyb7mG9UkErHkh6PSEltfvRlau+NbVijAoRpvYMuFZCGPPAYAlRjr3koeYe7034bdBAZRS762sZM
s1EBKwIfojFA0f5zNZgoile+c8vj6QMaQQ66ojMLdlQk4jd5jVg77GxRV1dlOdQxAycMEfZBOwZa
ROiunIc4C648GMEq5ujLUDYm2Xlds5kpas0QNHApniX25+3U4SGaBqo/30+4fsYsBapWGkSncSag
IIRSdBlLr6grNU66H/kvikw9LsS8D3GANRtHuy9f+Zidv+gYiU3hbrDGeTzvHBnaOYhuP7iicpur
5hFnLp475fMrjt0fwrmjkLHnAQLVTQwgePEl5SV4VZHrybGLkxFWnh33HeJ/y+tkeTkIGHGd8wAp
0qoMIMrt0jS1/KXSkXJiyzzHpU0Uvpm/7xRUWa3d09+3v//3R/h1oBtMKRi7NNyKuhVooT8UUANw
Or7tWN4OCHNIo+KFlvuaI59RrCpRoEb29SGLS8hkM3eDqMQfme7r5HBncRd0CUT6m6BNvli+R2Ig
uOMOjWXm3EYx9gnQUc3wEvP7mIMScC0ip4m8Eq4sVZvNuMRu/SWIW2Gw+E3IOMnKaTVsGzufezTm
PyiQrWgJWsqq00SKKYufU1ix6yLAmb6ohfgGA3zQJQrA/d0Nkna8Nmd2GBSDi5hdikgu/0zrNDVQ
Lj7U7SRVP3uF9kYmP1qsb2Sx7GVqwnqLlT2yQsqKVX4tGcE/bUlqv0rzG4YMBvTQwdw4H3RJJ9Xl
LuiMVFsENfzOsCPa7b8CIkJiCOYsTuaQJqWhcgmuFbrZBH8E3TFCBlTaTFwoYwStN0fB7WpDV60g
JQhIrd2O2JkFIUFaIWjonLKExfrAlYpnU2d6l3VHod3AoztBxiC2h40BN9t8mshJB0VoZiXiIbsr
a64UoNoe4Nv7z9YHUXNOO2Vh/XrcDMidAnWNu88VOKoXX7IM/H1HtLGG3ldX5vP08CTNn/tW9ojT
1YnN4oHUDmzAMdr/l3gtsYZ5xzMm3ClaZqDREfSjYj/Qn9uKAgi945cv+bCDwcdyRJSNUc0l/eIC
g1jhqW5mOGFyEdsGipUGW0/DB4KvXDDLzXefiFvXfHrJUMZgRtHhXDhndv0EiWbkji+wl5VxsFQy
D3v/uP8qTh7eI8unu8qoughw4L9mktNPSNgG/5/Z2USIE21E65dr7jpIAUfEI4T1AzzYcJi5eada
ka94AU+B8NlIggAtCy1dCiuYFTWSxoTgFq6GP1qAhNGuk/qrHcp7EgGX4UX4qlSfqQVn4zAzdXQY
02pI1a/wWjaS/seMyk5mwgs45wNuKNc/7hWICQsn1D4Wlh6lwi4wIEtVW586ErDM7TuFwbeki1mb
SoTruhFRULBcR9JpQ0uX66EmTMzx+H22mVU5pLitIjipmgIAy8wGsWLR/UCQaGYQJl6oekeXcX8n
6U/rhp00fEAGHze8NwPeBzYFEVzt1s1iymYkBNrXW9eyZBWYpb1q4zjEGN7yAVfQ5xb/FCIsA/N/
K/R0houZD6HDu+ixKOhxPFWLnAi+xyxRoLBdvzv9QPUyAGOjzOXugPnwQJC866cjkr1bk9gMKATU
zoldfnS2uPGWkbldShZs3X+a6UO5fboQx+59LxcYaGSGTJJ+P9MCz3flJ4up4+lrfvxpdSmbUudK
R+b2OwvRZz127oOwuPWhyGDwcBnuEDdHBXDEjzXc9EgR81oCmlwVRGALOYgHTZadbewdIu3KUODN
xXIYn4+1cLOeqVOV787alMoHUo1SEe1wB39tNVJLzyKUSQxVppAeBbXDE8fKCeJ/ssWej8DLxicC
pPwTs0N5H3G4+FrJ3qIacUJRZ1hSyhFIiyY8IbfWVBvuC/FH0KfAPiPeyqRmm+nlSyTgz19eU4s+
kpTDQHyalzeHTKEQ6O7VvI0VNV38BAlAfxNZK7VkSFLBr5PK4dAVPs3BE+Ht28gQLKtCE4U1i7PB
v7vu6/eDAelUWgYuxo2shB+QbSJZOJXdVsokIsl48IxfPjatBQFsPWQC7pLQf8Zt06IiOC3YMjaB
yyggBj3yPltkktBkGMobeyhm+9jTpgnyyJcB8H3XuXi4g1o2TLdlAMnNjah0gFrF3apDaeRV7nv9
ai/O95R2dhSF+vpXcluf6O7qoIv/W6SN5HXBfDkzeXXjCDnSzAjE7SgMT1hlVzZ5amwUxq90PPQo
Z1zRvmN9N7pQDyeaci+ZLgzSdMbbSYckMGipbEt6DE58imbLN1g3nKOwfx4RIQMZFIKbmwrK/LIM
DGUor5M5b41R36O/9jV2t3RNf9dZH27Pqdcxwjx+fwUNHoTjz5U4H6wCPMx9ptkLvdqmJoI4MBCM
37i6tNOg2hCiQp46cTZx/EzQknUBShmHtOATf4huz77x1hS2A8wAU166SXQ8C6mjuryZ/RiFHxTq
TEdfdHgd6MeMDIaX0WAYAU7/dZCvyw5O2RUaYOQAnBlf8+K2bCtA9eR6itkV30FKlsFDbxxrH9Wd
uHSFvmH9MHfD6dMxs5nrIhrps+1KNxBkGQ4iVmhlpOacs4Gj60CVW4lDVhwOWNYsXcaqPz4WObg+
siWoMxvfpK4S5KDArjQ+1IUrfT8ueJ/xWV472rlSKdDZ7EWB1NyTLglNs+7h3H/FtzTE7zqmz++U
fQX4oNfg8SgweKe/iqQCQ/Cn30QgKeDR/GE94V2xv+sD5OoqEtQDRrkUyZ0EegFmMwwX3V1DTcq1
gJImyZu3F+WquMF2lvo5JwXydQOocFBqXlacuCn1S3LMvFoJlUG8GCVe6lpsznMK21YAvHAcJcr0
RwE2ycDTP4Pcw/viKD3SFBnMgCKw9H7OyMxZZAdYtOmb8bQi0gn2mgTBQHHp+CQe+EqD2z8cWUBk
UYvaq6tALSmQblsBprJdR0A6bKKkB1GdPbhj9hsjIufAQb/cmYK2hUEzXjvWFj3ugjtT+TbURfUK
27JbK1ZRMbyY9ywJdX0qWxVfpzscAujBaz8g3i0IO8y4nvRdEN85P7ujEUWGZSXyJWrZjWfU7cpM
2DShahIctq/j6t1rL+811F/HP1WoS/ylTvayqeXaEelV8GOPNhSfm4u/WmFjoZ2Z2u1lQ7bR5EdD
pNBiOcGqyg81IKhmjIGacserxv9reMgEcZsrPNyfI7MOzAo7dDhiLAoIS7QBFmOUsZ5m1wVNo4jV
1k46SwifMlpH4G4osWzglkWEMjBIV42ckad40a9TN5To+X8YUMi5+xeZ78CwWjElq9VMBp3EVMc7
U+U79wPaPhbFwV2R4qi6ScF72SAhnXSi8hpJlTDgIGHHksj6RIOR2pgdBfRn2TPC/6zKzcSoHZTP
BRpdk6nZ1PW7EKMk5JgBABzb5oX49cmsiX6K/gDlmBA9OiIfQ6FQk1Hn6lp/UxQV7PAYKoxWesd/
ZKySIi0XuIhQYqsYrq9KD98DS+OAmU5Ni8slXo04BWy40bUc1uzeHL0XKP6ReH4hlHVyFCwd3zb2
R7dtcovp+LnTCWzEtRGtuln/Me2alMPrYVzlieab7pnnHuLXNjH2NzWm0LkA+Xkrtc49YasSR11H
y599+509qGEOch7Wc61ON47d4Y7PURzFoE41rAQQDr28RsQWSpm4UiJwHqiYMgLorX8kkLLT62GQ
t86TF4XzoO3h5gsuGql6hH3S12wO5MWY8SDGHmxtL7G1ezTK7I4ruJxkGpCkWzToWN5C6B2JNBsV
I1O2Y6B7qqMprUc7GyCc5h22csu1WM5KgbPkLhxO74jUpJpNRyWZPyd3Ips1aaeEoDbu9cLMxZ/6
z+OCF4Ar7eBY8O8voH5YVyaMMixl1x6O+4Jx/KzdGyq3GXEm2vgYBJ86469TTKkXpU3TNaI5ogGZ
zta6uLTUWlTYt60d9zqWFcRb9dU1T5C0NvYbGMoNowrir8Q6QATxv94tGOe0amRTKH6DOauvzTXH
XxtzbwBcGVsL+8hSl/Lc9ciuap6FCKzhJAA28XdLJOtbp9JVbJY6wdgTwWZg3glt74KqovmebL9x
9Vb+xae2qMKdycW4cwNR/0UbzGucVu7nnmCZsb5081DVkVxV669G/OsDFRF5FIWZlM5eq5nC4KBQ
4knyrJnI9Gb0bcjOSbRXjZXryYmq6x8HCqXhoVehefJHrHwyb+K9VxyP3gxGQFN74esZHzUnlSSR
1MA2gIIfuhg2ekbugdsr/dQ0BfS35YiTVshgTLtCoOBHc+87FPnabQU7/srwfSQN5Qqb49pV2ZJd
lAVjbAUfQJEcyveKwoeJTtyLhzHINLpMP5kquayvwpyvSQt92FE0bHMLs/tNOAZ1XDLkop9PlcL1
sa494JfZlfWx1kR0iZfmvkySU0/ysr2S2y3ILxzLE88z6lwntp8HsgNBrO3NnPMU1AfCqyZ/LDLS
uxOsrDWivozUYMCiDPPujYBiowzeU4VrWhh7mJbkjwlKrnMnlLlWfNIwWTsmgWpW9dFYuusNaatX
C+5P3bETE+HtQJNWPE2l2HthbXgnzeErpWupPNbQ4eMSy+Y3qAzYArvzU39430Q+dSGCKp04ZA8E
oucWE4yY8GMo8z9ey3m4cip/zblEgNxRB8J/JwINtGE3W2NQSVoHwVZ+ATVtCKJ/AJAPzn6my5Uv
FA4iwT+GvoML5uWm09kXUZ72HQJVhmU/BVBVC2U4IA6qDDte6oULwoIicpNAQeDq1OUpepmZaWjY
EBDEdbuHEqVhH7dyIomXXfIpxO35C+mYnZjUkffVsVy+jN2mNRApX0zDGdR5MeoIemk4QOtIk95U
35Kp6QCkZcoVydCM+52nmbiMNm4b4guicPGe4kUtawh6I3/p5Q1NiE5QO5klwGbH0F3wirdtYN3Y
SeW4L45HLqLCG7s93qfe01iel21FQnQpDysT6EL6/ChRVkF/Yqwj66ACAzh8BrCAe0I/GakOZCau
/FRnIsymBFC1ZdavN1UGqhruWsceSvubWBMamrSY5MB4IWgbA2V4ZKT0fZTjXuM6OUX/tfGdkrPJ
j/mWxc8Ar3PUK1RC8eDsmzb8u28/Ro543HdFQtaG3zD8uJbAx8Tl1Ruzdp0aDIn41LtB0+eco/Vr
m8dN/SbngJHua/rmWEnmlDVHGuQezrjxASEyh2eNRGE9ayE6lix1KIqonrNR3Ny3MrPBsc0KGG2J
Uyal1yGjS6eXZLHDvstUieKsRQEPAFojryQ25Utd3+iCgGEJXhxC45g/GRtWY+EwD9smQe/BnuuL
yOpyLBFtHkqbe4cnzLdj80BnURQsuntQprH/blBHZkgHnZj3MULMWL34H5atg6pZrZI0CQ/xJ6BX
Y063LIaS1CZ1dDToJ0Z2jnTzJPKcHVCb2J0XJqGhAq+vVc6NgQGfVmfWRAtNrdHlT13jqhCWrrk7
JyFZk/bnx5baO+rfiblIKO613kEpnBlSLlKjsN0XphdibCQc6eqCPDDYFD6cmPTfh7fK5pmz/Woy
fB0BGi2oQ6VYeHjQgakwYaGO8ZrV+aLlqznJ7Ca5VIlQ5/wPy+8x0t8Il5DZw3hhnLrsBnZ1Y+WL
CYt9KTDu+heDq2Sm2YAHzVqwZa7C0676zFJgyzF55ApTyhdG3PPwLF21aygbQthqdXPuwkUr48qX
voykYqmxQbAyrw7K4MzX5skc+LA1PM4z+AE4hAD2aqEdNvI6UCHksM/ZzaiHPRZZdh2vFmEjLeKJ
nSSKaNRrGO1LGgPRyVEgJDmnZStiNRFPtgTzRNoxqEXdYLpBXWO2PMC8bgE5JdTndYBWGYOqrS3H
hUvfE0XxJolH8s7Rt/b1pRTb/ukJkgzu0vqPsvmM95AXc+UxIMgsRnmKa6Fy+JWAcpsGQOT3t8Au
lYPA5+JowE6Wfs2laPhy4v/oElBC/AlwR2fBUjtbKyuOJ54qX2YzOsT5XTBesiJN3Yl0mWkLqGFa
L+baSnowGmtHB2xxkf46zo4OD2cGPRP8EynAarfCM56CIG0HQ5+9wrq92r9xfqYif5pTzOvOxGrA
prs/S24F/Xf4odV2BRqhMC9Nw8abA5ZDcUICjQNFWG0EFw/UVuWEZvQsy/0doqTVulFWAy/AbMwm
PyWL/crK61iM3vDtRJ5R3n2vFefajS1Rx3kIQrTTPh7njwHhh9TwoWqTDnTzdkdQJg+5evbNUqfO
M0PvTOz4w93a6ypRptYKTzQQhWS6a3VKuDrJ5fMfJah9P7YcA3Ap1fwteCPExTvTOekLmOyA2Uan
VNNS4f/Fwv79Hvq7BHhuGU1MUNgJUu/YSwgU+WZpWUHHpRhftBOkxIS0foqQh8q77xDzc85Zp8Fr
4q6Fx1e8cOdDUpI2f5lZIYoV2+iAKIwyHF+m2j0u8zK1K7CmSkSVUAhfG16MfIauryhsCI4EKzzb
QDrXYbZbqYAIZvdNgrRGJCqlT3ra7lotugduIfKlKCxWHuW/K85/D+nD34LKAAzr0qP017Euhcge
+OVfVsYzgMQHjAivSPK8M52fCCdbHbl9BKtXyXJZ0JI1dRUx6mYe50Gf7Or/Da/Lsd5FWnVOzzE4
ECPyhoX2dELjpXYgCUwC+RW5Ue1qv7OYOl5DpEjy7E8KzYFQMALYtqC3+MkkgwWoJZIhTFTK32rQ
QozWyke+rLmU88kgDp2zBqal/FZtXCnQZ9uQdgYReGg8pOuLwqQaiXSQ0oz5x5vjjZidS+nOJIv6
oAIhRXdB/qhGr3t2f02uPJPzCHgKmrj7ehsbI/UBo3I+ry/YAmPdcTkWJss/iY8WFS3G4Vv679j3
84UoOlUUfKUyLK4KCGeM69JmVSLVCJX9KxgsPKn182B4sVMTVTixPLg4E9ALU8dGL/SsNLzw9L+l
lleYTv2uXk6vQCxMRzzVW50PC+sU1RRlPbwKPu99rjjb89JGsWjVq0ZL17j7l9PpIh4pBbol0LwV
44PjpfrwsI7AoeqVq+G5YrufclCBy2Dab7xbLHh1hGp9YS7f1bXE6nSlf4+qlfzF0I9Bt8umKbPr
HP47xGxtJEGettGybCPPetL9e4pwzsYqem/NYcAmwyamVjXhffx5V2jFYfw6mhQg8fyMoB29z95t
r4HbmaDWwCVo/OqrMDyKUdD6mT59kwW0FJAjRZ2qj7D2pc6ErNETbfo58mp3B7vrTdSMYsH6H5Rj
ZLF25CsXVFwnymgzGVjkZRHaGz6Grx+0+kh16HBIxEeekbyzwZfXYlfDzHDe8i4FqHuWBKUoAr0N
u7ntkqxj5SDYErNfyPV7/C7GFBF9K3IcRyDLpIQ7mP3BGyRSAah+0QcXCUQNrsmrF+KOQ77EJiXx
ZHF87Zz9B6nTE2TQjZJb+asImRhPVaEBtK7l1WcwmIsp9VewyYNdTQX0O6xRt/ujQaYm6zftlrRC
IFVSGwuHK9etY3wfGIxD0JzP0WGoXs2UOonw5W87zTAHUdkOnhhaLz9jBwEvPeufHR4JZqdo26qw
BtswC9tRS1ypKK+f+kwsABIM0KplzmGegg8HFC/pmO96FlH0CjMZ17NWmqVxcJA9SY4dHHoOWvhS
xMcduCyAqI1Tbs5Z8YI/q5G/tMw0BX1wu2FTgHdywJ0Zj4Feub8gdM2h/DN1yL+fLyighD02cPtp
br2r/md5CnURgWA3JW5gKVLEJdcPXBXNsOLWAUG5hJJoz8G3BdKsMQrlG4edf4OCiNyXZIUYAXP4
gJyRFH7tr6CW8nMczbgnzot1VqPT8tuUA+FWpJIkhXoLWYADt3zrsdcEKchS7jax1ccmt4keUXso
wSbNuuPdessGtKHRgxIOOa2iUjaCFH1wTOwx4xoZMvKzgc6P9zgNCYtP6yEE1H89KOsT21XRGl8t
Ky4nZgTSwi9SZJBINC4vvz38lcUI8VJwB/8tmD0Vg/mNSmpYdlME3Gi1VXwYuiyGHiGlyG5sJXoo
slMqfareb2W0BDIRd8VO5ElWxS4eu4QTehpFX3sXTIny7FGvQ+flplHdGgPDcZcXAkpcPRZ34hJg
3+VP2AoecW+bN02z5/IJe3uJGs1mnpyBcKIKjEzbH8SdU/Nnjz8V7wPgz1CKBIbBx4z+mDDPGJz9
rfZiXMAuYy/MLGGhOp+/qQXQThg06WXGeZbZVdATQsQsiNEJC/+sONw8aVAytFqWSyiI+I5eVhx2
K4PrJjXYLwYnBakAFl9f1PruJNRpSzlxmrD2+u3QFA7jou1cBBs2ADxLBCOiW8LP5pl8usFA1f/A
FPMxgfFjEtKKB/AbvaAV4gCMqK0b2aAOEg8IFoN9Lp9tgqts0R30suSZfwUpg3Pnb4ZEbcWW1AAD
LSwRt+QodqIRsvvHk5G1bmyc5FIUSHJ1CWG1UnzS2o9l97LHuLMdeW/UPDhXzLNGuswQIj1lr+mA
yOOfKsuiwzdaKP3iFrhEBrZbfrsR4QL6ckxHod2P6a1lpOD50TliItsSvJZnuw/4lMxX2HEf3H/+
j6QvP2AwtOpkzc4gL2bPm13bVB8AVZXy6tTMv9ouybYENBu8eABTqFJMGwL5/FlGxWq6Kby8P6bK
ETHssHVFhDdSMm/3jT+nF/JoeAusRRFC/11Avs+S8M/IJIGGoxaA/V0sX7ZtCd5/dzhLSa6BA0Xp
CDJRXIc0a7XwZpkREgUVqbeITh/Zuu9lBmsDnCRi9a5ioUmGsvv81QDMczNS5OgkuG8cGaCnz/xp
/e690BQolUcLD25CsekecQXYaAbgO+mhYcVv6b/y9vrZjpFz3HANWbXUyt1KLxXz+OmjkG9S6xZH
Qu4ioos2NOO+VlA4V2faMNdjKs7Tbwmxy0VlRxcmIDvEnoe85Fy/VS44aBq2j9B7DhSHsUqS192X
e6Oq9ERohFn1kAunsNOkGts02go8VrlaieCnbIIgyMB0gUtHq2H/bLV15182Kync7ll+V0sfIVn9
Tr1HizflasASElDCw6m7uxHjflwZ8nSdwP98S9BsvyGg3IubzDQ4Hod8GOnYxzYLdaEa23q8SBln
F6oShiPGnAUg6M3cEcs5udMQp6mj+mSqJ/CXYa/gFypd2iTcFrTzAqQhKQnF4VIJhI+UrsfwSNe4
tZWu9qM03myW4OOyo05Gy+yiPzpvJFIcuSyL417kT8/Wrvh30lXGrUo4M6oaaPX+wA7cXoMg+Eqr
3iU/ulJ91CTwkXvYi9butG0COWdUxWJLap27UYGUgGNZKNwL0vPT21rWmwyWYm4Z29BOgqU75gUB
uvigKBRvmm/ZgXThrmAkVwZQBYmJHaEybULSD1KgtKE40ci7jVhBQCIlgTujwc9T5i4Vzfy4JsGj
W9ixF8gZKE8pNtLhnR9h8fHmnkZx54pST8Tplqd6mjjTU3Jas8RNsnyDrbvpOQvY4bt4cNoRlqvp
/acp0r2afOr2Is06+ngsljhjhtlFglDOTr+MXprP5WH9UCjDXrZZUthmrSsUOTH6qpEULuajrDlG
e4UHfy92hkx+EgKRxGsrSv1I7qKr8agH+Yw96kolU3AbZ56tDV8aYQBMWvO0rDeFEk+9fzmjrIMj
RRk1A5stvyPDgHHsqztBZBJ8yIABMRr2971sqEz0M632mVjpNVFH8a1aPFTMOirmSav1IhUaIy76
ht+Z/RJSvsOpkD+iRAeHQdTwr054ctDX/Pb8w1MDVYdoIlmUu9IMykGjoxzQwErnjn10Bo5sVFp+
Y57SHi1jDFSPAzv7yCO0dPa5s1Qq/m3fTtJX6ZAArlk7cXGbg6r7wquYvoBeOLdoxhfnu7gMQelt
yFlmWsCX7THVVmnkcB7MLTP65EbvAtPTS6YIIXNN+K0sy6NSNs617MPLYcg8F9W7wNksJ1RksHPX
R9rNaXUh+HnWYARBT/9BSN0LLrT7YBFKQWUYohTCqxfJqOMH5VW0cSeX0aVLcolej8zghqEUdFed
nAlwPPYPpkuujL+i58TdF76E2/t+Mjh5zcA2vr9zMnDe19OatDg4vNWNVZgZwqdOAMlnYYR5nMSK
rQbsqFrs7M8Impp2sj6YX1Itzj1rQ9USGD+wMG0SwPnwumqKjSI7RFuvx1BvJhh6LPntalgvw74V
bKweZw3Giv3oie1MaXudcKH3IjxfFydAo/4I+HKkjgXn0wbgZgOxYPb/NO5DZ05v6m1P08HF0FHJ
jmbukWxI5wf8fOv2XtP+PEm1HTEkBB9xeDSQosr/Nh/NDm/Wth6OaCNys77dn9mohVf3Aatem8PM
o+P9Cb16Tj1YwqSTHy1LwtGlDB+gR/PVlPGjkRiMNQjnat+/Tthj3YXZSEJb6s4XByGc+aLurjdk
Q4fkz4MiwO8i38BAifm3CRUNpQHZuwCzQWifHb6EWV2OSLxaCRuev8FjT/AQJF+Ze3CL9uSNWL6s
NqVYvrwpVtDyFFmNdjbLuCgn2u9e45Hwb0qg75ytEq6ND8E+UDNL9xuiuoTBbfkWvSzdLlDtCSsq
LQa5rNowe3PtMRLdDMzRYnkZomWfFpoFX7r7oYm/OK70HmYDgL9eAG/vXaimz4n8dU5I0I2tgdkb
8DnzezWjlLG8hlBwtU//x4JjbEGi+u3v8ol1+o/qGnoVh/RJhQFmcMJdo/CZCSp97IYJ2yLiZTPH
7swhcoe7LOH6erkie6x4/2qOb9d7SquXDOc1GwyCrJtSc77C3FWR7ACK4rBZ4YHgfbNziwKrVYf7
KPdGic9y2wOK5CbI7T/oEnnNQdBPcBKb2Xfhqyhs2JNnnnvLCV1RxBOBLW/L7QPVdEjNRRECu0bM
O9+MQ8AFOFXBk3+EAVdsBbgbk+xtE8AZY/zcKzDg6IeRYV0yHQbmmTi8+3P1O4wNRbhcvP52S+8E
ImmJO8mRQYn96alb1Jp5vbeQ7hpy3GV2vnyqYigmX7TvAONaz/gHitCRVH6rEyYeR2vWcIQu5v8z
xoWTZhNdXx+9jDfFGUJRSiDjztvFZiP8hwL4YUUYyhsh8Cm1NWqhR+Y4iVsQfOKdhvPus5P62DtO
13lGI+oi6O81OHKE/T1ggFssNMST1Tn2NZGE6aSsaHtvgjY/qUxZRk3aNlRHLUlliqZtSPdhikrj
Bdq8rIR+Xx7zNsTPhJ12SbI13KucJ4F2z2hCUWHHsZFJ8AZIbZqCugBCfa4cVfwlNE+KZUsZwDAm
9WUtDD80Cv/9Bkrx+K1Ajh5cPH8i0EGRW3blzGLzcjZK69IAjp3ngnHI9sy8RlZi/GowmN2cPsc2
qhPw4/vcZCIb+cprmgyLVs8iLWVi9KiHNH9/PmaXrWCTFhVyRmz+RJcYJMU26+Nimu2urqKkBfWG
437WVYQHWqtR2+GFWkFmAFoT5YJxMGCsDlxa0rfEKJ5Eq0Vej+8OLTn4jjrVj8enAtdyHV8i8zZf
1/mJeSUcm6pEQzXmu0MldHODvEdEEIKmeJJCcitn03ZhqWnq7hc1IuajWQkggJWapj0kyiv5C5sw
JddN6Y0F8ArtATW/MCpOSTl7gdOUqvlUBpxYQHX+KH7uqbDaXhKUHPo0SgcPvaFGPBwCH+L1tqBq
1KJ0amA96gP9jotOwq1knmA/86w/lS9XKrND51HlQ+9hE+Ere9GTcTpnWjjLOe7vREN1kzXEYL7e
yz2W30FtN6wwoktfrBzJRur9Cyb/JZCJSDRMky5ZjTeDp+uwEoZHvbfDZEsF2Ka5ycYLIxzegwdU
y91k/fSxLGxR7q8t9WhWAvdmxeA6t5iWzIY2gOM7FFCUPcwsCscHBWy2rlXp5kQmmdihyTF/YAgT
+qDKMrplbULZBwWptNIZ5Ac/qWtXtPGni7X6X7geMp9YmxpubkXdrLKwLUw0crRGnmDN/783Q+8m
r9N7tMDpwbH/+pZv5I1e+PAq558lytN/ob6hBCwT8vd1OEle528smN3jqHAvKn4pDadPKvkLJEGB
2jgPjGyVQAkkA6E46xYZLhBpmbURBPNPEyTXydYO02twgSdJhNRwhYjtrnXjpJ0Ca9ERS8V24EOi
h8BMtIJ4QcJP2dB48P6WvVAj9SP+eEk5/+xinXt5TZPieOWppLJSYrqvyN5D/wFQovDhUk0x0MEP
kRYFYtIgVeKDeh1mQN/JBU2l5R/cdg8yoSRELBeoPdf9aBVWT5xWekmD4v5ED0gw+k1cGsjiScRk
0A47rAgBagoapCAdhQA4bfmYsDAizmeXH7/egHqvrZge5FPDlSYtlzNfZ8n5tphg8Exb/1lJWY3V
jXykvYE7i+yW/zUocYBJTTOJfXIo6BeRoOiXdc1ySUmMp8KpDKYjIRt6blWqgSYQtzQmybBRy6ud
vyBNzhMQjQiGjNBJgnskFfbHlsaMMf2kBIQ3FVRlYVuKXl0MaDvmN2mNpVa4s4oPQzGVsMye5eSC
k/zDfkzy7P8wZ1g40lptLcCaW+OncdiHCSiKUpeh33uwDDdiLWQj+UXjF9VSJGiTRPFFhAmAN4cF
EUHO6h0vc4bELYCGSv0ZKLoC+CpXV9c3qUX5nwUfgaEqnUJf1u3PsGpP+rSNggbf+L41jhKqE/Nu
Qizr7BejJDqf2gJPBoR/oHQlxlNh4i3qA0/zxRaeA0581kvhBRqwyNQ7mjQctKKbHQXo5aa1dLF4
Q7YDWapb3MbKuA/jibMEQnfsjasDXhDI+yqjp+MhqxSPpniP3Uah1ujeAKYM6uYb9SkwaJnyr+1T
7yb8WrlIaC6OT4biTVB3qUTyvmtyvPSIlpNfnvAly4+90Hhc21JAWUHkQ3nvpExr4T7t7SSw1L6f
xHF+Qxrz5z0HklRQFPwJmseUgJFwEH8BIlfhtyH56SVtItl6YFVmiHWwl/Ah6zNE/MissdPDpwsA
16da+rcnVbV+uHjSpo5Ht5p8RNzmqCu2yp+TpH0yqJyt69dJGU85F9cj2a3ACqOW8q4bSpbOvziA
sc2tqY0bD6fApy0g01QivnwTwdontD8wWF23Jc+2pYxbV42/H8pSZP1eN+bbPLQKPU0K2dtEVOS8
WAwH/NoBwWsvt6QxoztS40cBhBcr6yxPfbgnod66kLu7w8wxDRAuZRSsL8OpL+EZ1hP4wOT+hZNF
lHaw8tk3QqBkY5vYXlk2DsXfFedJFshzldXsYtDAwe3PVRkTartv0re7ABsRcRXzHI62P903bVvY
YA84mJku+n8OitfavjAVbXEiv4wJ1jC2p1JZ9PwKUP01xicfmaqf2TCuuQF/DjLkRiwhgtcSqHif
qGsmk9pvQAsqRdOvHObQG/vzbKEYcqCAE2rmXpHj6iIz+Mw1I66AmbpiITuJQl6KLn+86KQxE7uk
vseyIM72CybC5yR0shPYD1VLKi3GMttY3FJY0ewic6/g19B5+jRGvItYlJ0gSzJRZJB0JiTBrUZZ
Iio2ghXDtAqXNooKCAk78xhtrSYmMcXRZMlAnA/3osjY6NZJYZJpqjswGGfpcVV9mIF9esHZjp5J
SW8ufHQJCMjqV0K6MTpxswimmUFB3Jrcphvk+FuFWb7cG7cJkR2ZSLkzjH1SqP11cQ+jJqKejAqR
mLj5hh+5pgqtNwvW+JINLJiFMnOHh/Qj4+cL+qwG1HLstNy1uBSyPbwPYwmmYEdE+F6IOc37c3qr
dsVGkZy2Y9zTX73rKiDLSOPZC24X4sFCeJFO965HV0ECtP85D2dtk82hvWougKrCZ4UWmvlLvDFa
wArnEsf6Jemka78yKzh+zUEdyTCIppgaAAouaK5iteOdDSv/hJ4FOIebb1eJNAGrhFSOQDOZptOC
8mdKK8Loqklagjet9ko3NP4SdhxNfXGCSE52n9CkTpbhQ7zOcUSYuFJDixdqWcslXIFSFucZIl6l
pG+8woxkBTlXVFsQUJ42/iugs+6Gt+vrIV8/b8SROmMIrHyd3Qv2Mx0S+iBLVLvWdK6nohERMHB7
Dwozj2Nmzi4e6spgH99S95aqj922NawL4tajKs4JBHTp6lwFrWgDTaz1rQc1JpfW/YeZqQBI0lrb
xmWZz18nexgScCgqTDW/tnBAXaXtmTpmBsUP8QkAF7e7JdyedH+iEhmDZsPpPl+bjuAOPTEkW9uy
RUcAN7FA1+JFjM9T3gUWKDHe7EPbz0FkxfvRrEKcWYrRsNN9T2TmAKjYlpNPkHVvBUDEz3X0zo1g
bssPL6g4Q/NKQ1XIJXMN4H3212rOUjYUugB3Q8fQcrkOk6boxhRcR7GEvlieR74ojCG2LZ5n5QEL
Md9bvuSITH71LW8yziewFML3tZwdYA4Zj+swDptPhQssYicXuCf/xXM/IjnCZpxrnJQMhgZFzYTg
sq0/7ddPuaR83urcb+7wCMas3v4IT1HFDaT7Oxfjmxa06vrL6+C9F1SyWixhbLhca+QtlGkMWZnT
cs6ye0hdstRQ8p++tkWwgdtPGKPnE7DgqUJs0jD101ObYuRdUFBohpg6pAbRMi++DR76bhbI/v54
k/JQKypXfYNzRIvlM2nXkONPc/76pCpam9mv8KC5y6x+NWcl24Ci6T/zL5tUQDnrFaqu87FhaSBk
zok9h2P2UGFFE6ZfNH2L0a7gjXSsZhWMYI0n90pXLOXHY0kvYGO8F2qWnDEsGgkZgKCMS+gtqWh2
z298CrfMSVM51MXYyGZrv6dqhMPsBgWOp5ltg3Dm7+Fvx/F+Sc0NTnNwmoVzBKs7Uk2SkOlN4okm
rEhNyktQlbVnCobh+BhQ+PSzXKOwvhuWBxLIpczcLYLm/COvOFA3cBqyodMmwJHh9JIwwNyy4KRb
HreG3bML07IJZBkCorDiEkUYbTQvHa5y0Z2P7kCtBoJWcD3qcHitwEaa8zQ5QoShEKqmkiIEAD4L
KzUqZVv62i2V42tHsRf+EnHi2ja99wSu0eZ8fEVVdHWwTBKCcqmVeWGCq7YDUZX2AANhr0gN2yL/
fo67qDdTyBzlCUJitFm2JKjvFFc4/iTdiRBDbUcYgPzCPLS97/UdSFgT/TRgKVg6lJQLX9E+B9fN
V1xKGPVWqBBtRAeIjg+U3alvSfDFds0noeO4g17Hq/mspF8pS2XpeQ331vD/HEvxq3B3FGjfPhNK
w3bujnDKXVs/+d1RgWzR4VjxdMG26COo3PttBBOyRC+Gsl58zw04PyOZVz2ZkcovaHWntSyiN7Ft
QPSagsCzxu2aa2a45FApXcvXRHtWpe3DpcFvf22iiL+/1v6XexW9XRqEUmmmS3JNgMaV8myl6g83
xS4OtAl5QNYgBDaTxIIu/24NRVxVZ1Y0BIxubagoQCRXtVVdadY8ciB42pTSQT9oFGOSZfMkbCXC
53lRxpk+mZvoYfZ4VaDQ+lt+UDaer+wzGqA3LKZQ2pOfDxJfG0KQxZ5qBVgoV4rNBW4ikg+d3Fir
vFXvBXOx/G/yX9J2W00GoLaa8YdV8Qa88Vr6fWCr3m9+WUur0h1oA6o4Tnr3PMpFwbpnYghqssr1
JQEnZOS/3DiFnIRuhAuPNg2Ge8xbpZjkf0GJ0osP2cst0s40DwKrIefjHXOKjfIzR/erXfmynWRb
4K0q7ElVYQyle1yNQJdeuKU+FAMtpPQCDL11HUbqk0U2vI1XXmhXr5XO+9GOgBS6ut8lQZUvHEyM
JRduRrvb2ugJrPXg8yAd33YykLQhGBGF55nKuP+fmHLux3Er9DJvVuDxZ/BjPcFLdPZll7wjfv51
zpyD9V83XnYEA+Lvzkz6ZLKe8wtlIiky5bHzlxRpRQLD9TO6Ju6uSvQ62Chr+7wS7gumz17rKMDX
Vn1GdQZocIk0qNwTW2/qGFqY5pFKJg1AaUAUleHz6PAFMp057ihpuxOFb6xjjSN4gs5ZIFfLKOOe
Kg0rDlLLcxTpzs3V6V4rTR8Vol5UdVH/omi2ipk5pMvNFsnIcoVp8uXmNfwFQiY/pfiYmKKXfEXC
YwfxeAa3JlLPLHNBVobnhkfiaWaM6LKaj+c9/BtfLiMcUIVQX0wRGGvaigwb2dw2UucJJkVSOEIf
4f/DG3Cuv+k+zC5PP5EuMTDW3zF9cm/wcG5ovoM0n+Uj8Hha+MKGYflEM0jnsztoA6awCze7vAO7
YF6PwBmAUHPrMznsmu/3M5puJldKeRAmyIxFP5mEwwVF6vIC+o0tiQeK6QRCFjNBn1vxuHLnT1cK
4hDIhkyMNt9BZyKGgqMRYlwfP6FQA+Z+/8kJaljvcUibOu5Xs9Pkzjrk8uWxBpNAyht7kHUukafw
QhDR0G9Qi1DKNfGP92Ei27NGUxxw4Itk4WJ+4YbhZ6zH9D+QPvrxdcDTaKs2eqUFCCo+rcbNZISS
qVKrUpAMPmhNaHu00jXTittfcZSaOJvkQ0q4VckR6UjyBU7yBL9PsIGQf2X5heZZ4uTF61zTkf1g
EQlVCD6mwYvgcn85JfDvvDpPA4nW6YaEBYdJOc+RpybZEzr1gKy+JQFxS15qiDiRpbReJVQh6NXA
/+aOUeAZlzoprnoOIrs6YZnRZ2EtGxg9kE0LeOMiSSBQdYdH3C35xQzP4Bfeq36fU2EPtld/uozp
pDv38GesFyficRXGNd6Svt6dDSxK0sFb48DCY8DoEGNnT+n4ybD4iNSkBAERvrGB6qTQ2azC8n4n
sQEVWap9APpnBWHHRh6it9KZQAsCc3tL9tIQaikOjv4jY7iLZJ9sU/Gsy7ELHlr2qnxWDbLSjaHw
x5NovEGBk/uSpMJNUAMqWhvyxEZL+Wq0Jynn1bMjj/wYVApdbHqDio7ZwhvZ2zauuiy8jklWyuHp
n1EgtgomBIa1XCN38kKW4a9msFk1kMpJIhvacxZfM0PNPLEi+3amcLFOlZ/eKkRVd2Dp54DAuO/t
+tR6nRUwZ5h+RoSfkBe7jAjAI7aeD7kkKGyy4zBixyg+/nDDxz3GpAZzRu00Hi5NXp81ea0fFYPF
Rc/ScA+L7flpT0l4iWFi7v5vzoITThXDCVMoAJp9Gww5FC3B5+1tDZsQ4zduzD4x8Wgzcgm0fHsb
sOW8ofWyZ9z5RwN1cuULUYHtqo2U/8Zc82tCW9EgTRSmaPH4Q123xxwur8kTmWCGa7GjvTyt7gEx
k0AnpUF7Rv3eGbe744Mnslu1l1F4DqZXKFhPnonfLcF0YxC1ud9MzWA5dRLf+G8/4smRrXDroyMB
FKgkL/Zb4RH4MAUps6GT9HgErzVI7zP2/mU9VZegxYyNl3+OjnQyyO5oLfuFShRxvWrc09bo/xv9
RQrY4jOrjEu+QkrRhZZcW1RmZpIV41Cd9JT4aGoUqN2WyF9ZllJmZfYNQz/aSW+omhTA8RC/tP85
4y77nuP6Kiwu02YEWrJ2p5Yyc+ZnaTXNErVb9cV6pBiX6luVBl7JGR+e01WkhI0ym+qOpLQwo/4O
YViX5i9DNYNsTroNiEfWrNz8Dvwuy3bGZaC4EjucDdV2egNT0Th09T6NJHNn6V5aHmHCFz9cvZK/
gMpoSDZPq8UdNPqFBRuZ/Cnzie+ZHIiM09pv9KRVeOzL/PQaQwJUTYsTclOwv7TI6dhZKKNJ9NCL
8mEfs+KNhe0tGUDLYzDRpuaUw8HRs0if7QI2GFMTBSOciHdUC8CZ0UrUImAJ/4iO3nGupMLjSbFV
nf0aehG5zfDMeV5MVnAyt5e7mWO1pEaLvstwM0cRPzkggh+VpAKKt5tYZCCIwQHpMj5y6EjoQqFA
wTUnLff+RbDO2mwTwGcS9U1te3HkYupPCTFhV9xGXe12GYDPJSAYQK8Vm8l4EZuwZDOIYTFyrJqt
8pclpN6aXwLVV/yGxe6hwxyeLslxUuT8KFGmur2a8foqc317BQAvJeg5zY6knDJ34EajwV5usYoA
Dig/Cixcv8th7pR5OHw5bMORDA2k+MYkUFZbpibHz5Ch1vdXAn4/gKV4G1QrMoTM7myMt+gK1aL5
YaQLZdr9Y5Kq9l3Pv7kx6oxbEAHveRd6VMPYxQS8R0EN34o+ye4CepZVIkG1VkPUrb21ZT7h8zQe
EjZs6+R+81R9xUz94E70Uo8aRq0RoEue6Z+AIBT5seQXTEiWiBaS0fu2gcUHbz/dQYP82JxIjLdB
W3WE66H9Vl6Lu35f6wXCCYgW9USzttOzPSoWzOww9GfYAxQTMNrxnNS6WAfAAb1hYpfxxgz19TfK
EfKv4YwHHC/UuGZpkukFXJhVyx2ae8iwMSB4UoDPMrVKcUz5HZyziqQf6IMBOBxyNKsiqPAcg4yB
yVDWF1lkIeSTAXi3B3vSeKCTSLxeB2jtIGCae/33pz7Jt0mND8SRhSBtZWDx2xj9tXyovsdTK76l
ilV9Pu+WmI6UuNTTGmaTabNC/16E5yBNwEmCR8hBDiHJLD2evpGMqL64XyEcoATwtps+FmOo9Qs8
m6x9VUOb2VgZ8ZQsJgadf6/aSIGx3nrxXF88lpyT/SHY1fS5eH7JXjktkTd1w+ZrOpjNtaksTC86
twCUihFo/ZpNTyKiSvP9hbOAyJyzQ/593jCaEIyMozx6JEo6X2NIzV/I+kGnjoG8o+kBWyPV5hET
pELnOJDsU3Nq242X06+LHRu5QYiDcP+qcxlQI11qp6s5qGSMXMtB20XVUIOEKCqOeLJCsE7b6Jhe
vYs34CtI91z9juWF1PRgwjBQxtNbMKmeHoeygIh+bEHWR095N97QL8L8/3qevfcj6ZfSUI6LxxOP
oj2X/R/ATZyLksw3xEsXoh/5h0VnmFWAJEe5dl7mcW0KWHsjlhRQEmOxN00JnF49wOZHkSywDJ4n
klBIUtChkh6UCfg4wk3Bx2IZmKbAgttl0E7kqH8QwVvKSMpFNIkzsf3LwRvWNPEcuxxhNMr9Q9nL
ER+A2TDGjbQJINSLpvw1wCweuVsRfB+ep8OiaFV4SxbSnxi4ADnPLGOHcgVQnNzuhUAR3S2PwXRW
6/0t4643Zl66lWtaxA5Ez1UcttGebJYPic3zHd8ynN6esnrEBLgyltxMj5WHq6AlOhZXmPm/pZ7t
tcD0IZPoXqolpTgLAZUl1PrZtl485kc5HfqC7AQXzrQPEqbreHrGZnDA5xgQS6BiWHHG9G+rX4/k
cyVhKEAfAnUXPo0DcYHV1I/0nHV5RLFYegFMO3PBFp6tYi/tuUM5IwhzSjRxapzre/61PSUxvJ7v
x9SiLOv6sgNWl47UTFZE99gMXq9DegUdQ4r5glUJTCE0h7pFBO2BSD+y8kIVpn8lMFbLDePo7l8N
KM85dGZ+qalk+2qzUy69CoDgV2mVzuOK0u9evIpMnV1Ds9hXTFe970QjeFp9n5joDBdeaMq/Fy9g
pueKyVeokfC4KXuuJZUWyeOptvoOC/9+exftnsKOYVU1O9A0rFffj2R0olH6mN6Ys46CSN2q9OtW
pLJYgGY6zzzooCxKDq7FtTBL7gOobkoEHSh880HhAQhbqpSLvjnfj4DN6eIaXeyRy/u/FMyyhIvF
2ZPtsp02AFZ0kdy9fuxg7Rn9yyI4Q1gh0tqbVWJFPxr1MSsuhJIn5g/9sfyWMwZW7w9QfzoP5vr2
xBKQA01gGH6EbsZxFp/xcRSJpk7LXDOeKbDvBvxL+fzQMjpVsbRZuYxi2ya4SuKvvf/n4lPZahJT
gzTwr1hI1+8O4/YtnYG/nDH7QnsMmd8Abl85eP4fqtQlHpWXZ7J7hwuD8NTSdTxHNBC1p9V/438S
73OZ9YUHUES1WcJSKP9j7JJdyLK/N38atIF4BSB+ZJo8ZeqeNeZMuH/2wOSK23PEsIoEi83hcoQY
+miQdcJsv+aHM5gAGcheI2kxcaGA0u4qANblIP+nnexBHgcqExtIptpbYcO5eT036+TrZCjctYqR
8EcuIy25UM9cWB9MKOnlMHVSbeXAvFXbNgW+LGcr9KCaEwt/2WK1yYM3/l80Iq9MYqnY/pVAjWfZ
P8JAGCqRh6VbofHykL9LFqC1154p2eyKmeaL/ZGKmbQhue/IYC1krpFL9IMcVmPyOPzUNBpyhjDl
U0DN2+NuDHgmZJuDrwzNpVGezNvtuwngF2zKVyeQEd3doe3wHMExE9KWVGAzNJGr2WfuzPQnr7+L
yn/LUi3Em5IM97XXDsJVwsi9NP9ONNh7SC6gHLI7OokzGuBi1hfIsbrpnUfNnP+NQraLT9SZisPU
6QAj+gIDp8K3LZUsOn/RZx6QRGkksli8o7oFjTriK2yK7U9Nbr9lRMasXuVVSupdaC2qmQqatbnO
xDiDkMxAExXaggRJ4qgVGoEHktZ73jS/rhLwx9Hs69T/IcfFBa03CR658J5BODYiEVN+5v3M64fw
1q2Eao+1kY/1D6WN2b8Iwz5KGK/5KRFvimICPrZFsYppce3tjln9jvtrlS+ywh0SIfrtvneypyw9
PxXVjT9HpngPEPzxbYqz4xbl7w4dCnPZd53LQWPAA0rwCuqlZ9NPA/h517LPBrlbXT/f/ztWf9N6
z/eyYvzcE4x2TgcNwLPe0+HuDI8vDNwF3DgivZ112jJoMO3/JxrbyuU65KFK/nRcFoyDnf0jMIuB
9tUPDQ7of9k1CmLfWZ/oiHM0uLJeQjcGlAM6jxwBWjGU5V4XW/DxdKCrlXPhhBVpg3MZ3Ca8kzu9
QQCGbA4oaaneYTZOM8UeA0FyE8Fwfw1KkadCeUqhDxrWlYALqNr9pr08fowT/edOcVW6B9Vhk5/E
N32dM6E8Mz1xKi3dsKfxGXlPNQKCZwTnSoEvPbBRiB6bAtYPUjxXjA9lEvpLb/nFF3mBcdpT9s6q
ZcE6v7PUOFaeIIEh1lnO/R7I0fzznyYbYmbzR0XoGTVxN5annlEzUlpd0DZmkeDteluIfZkbVul3
pm26VbiLYjBqUF5uyLBkdAWPy5cbVKXRQylMRflnWN45ueafAcYC0Y2w+Ipmt0G22e+JBWoM3KBQ
gNmUI7cM1dyS5IQAlihWEovFRklE7fHl1k/M4TV5cwOrb6QdSq1XBjNouGimf31G3hv0WpLESKIR
twHXgg8+uGAgFb99oJyKfDaJSqs6FctIzYNPZ24rAlnDpA8DGgpJyq75Oa7NX368nOTj1xIfvfIj
yCi2JFF0yrH2IYnRdx7DQ/hZaB/au+kCBEIG+ZIR8v4cUHl/W5ze1Sk6An3qeM5ExzVrozuxtx0X
xWAHNT8F9YI5jZn7uiW+YUx3jdMWtlvHDavvReknLp0bExo24ovtX5GulvIkR5tm+HFcvPq1AW4K
yXLqthj9o7L65KzHSXeyGYD+E1okd+oX9WtYy6w7IvduB+kUV9xX4HqM22AFVFuQOw66J8sXsoeY
TwwNd35nlPP9e3b/GWmHrexoELvsb7wqtnmIZEzYFVGV/RaJzw/LSpnb0eykYgLddQ13NqgRjR+o
K4IuDV13wJ4qNI8sj65tiZrsEz3WCJWOrIoiAX97XtaWglBQOfZ/l2ezz+Qtm/2tC2FUTCzOU2QS
CdjhhdhGpKsyGiXOAm3Dt9LS0HHfeH9bqGTnUSNtf8BB1vBO8NDB4yb7W2nuvKC6wA9pNbBIc5JU
GJX29AhMQJ4zPzEl4SlQ5h4BaKd5cJO+lUKfeBoWzamLJ32kVsncbHqQw6o15fISpCXTzBkL6LfF
q2ydfshPg3Ukbykd+EMZd6Nnpz7uETGrdOgP7MpXSmhXvPh7CQGKipnogFYMtUIpFBur8zVx9uOC
8yNnqrXqdPVawXTETDHTO2wy+TwQf1pAP8/+rifC1h06mMs40o2KhxDqA4uDK+29Rp/Z1Dq4eCzU
sFIzrkF1LOYBEujCQybLBEdK+5Yr314xvFmZc25qg2q9Vn9GUVnLePSHD6lwGqKCiqg2G13ewq2a
XiOGpqtdtyQAL4cA5MAqxoUv85nAruyVunHCUcfxMUjgBxoxCANl/2dYV9+xOeNOPiNfUpKQoq6R
G6uljyfkXsbKY3cAg3Pr2qfM1MtgYtC1ES6iziv8jjja60uFbrhojhSPstJQFM/H/EPQuEfWGSNO
FF4/5eg7hQLzs10Y0pHlBHibBpnE5ow5Zk6L6GrBWHnpGwnVFPc9eYMLtyiz9qMy91Bp7jAJ2uR+
GvDF+hHUjOUgFU8V8PjjS8YOf1Z9NSKUj50p/v4z7TvXXc6OdSdEychTu0qlYmBhma70UbwlA24O
AoGwoFX15ByWCT8PO3FKsmWNhIVii1ZGafxxIsxrI1B193OI1XipV/UL3M1m1tcFsA5BHz30lsRI
lsbN9w6WXoRLQjxG0w3/EE7mGRNflxTViKRyyinMeNVDfT6gvMc2uxLm4ER9bDtEc6NGFaNPwkou
wRXZfjYA182zkx49JUDdIRv7ZN64+ZVj5zOzZX/sJQFiTvJ/ww7TkfoJ99ERYKpNnm56WScI4nBh
6vh0XF+PLr6831wgCKJw85v14KYghOa6sXYWlF+7TUFpShayALWAPggwdUiItj9ZFvcqCzztPCk/
gKxltapyjHQ/QMyWS8PRe3Dak4CKSPlG/jS0za2H0GJ+ig6gzw3+zuIqdbHgvyp/irUvtRehsA2M
kTyPNDLES9QymB0kETuZzs2dxwLA3hUeHTl6s3Xr0bAAxNgn8Q8m4Md2IdRHBrkOus590K9DJ5ol
4gKPXBiahXRoxAHRknEoWCn1+jHhEw4vIqjuaCgyZHSNx7SPoZtWPdOtyE/VG/uiELnG12f3jOOI
UypdSLy0FT0kd+KtQZTBs98bHP8UIZKIbxh56Y2PZc6u+Br/8thlmDXRWZKn0VLI5x/B7cshWz25
tz0OS/0qyzsQw40NlBDLFMtng+btZjR582HtYI8J4P1v1K5giSszbfutnDbtACPweDDQl9Lo5ZJi
bvNKo0wZgdDkgBk2TRr3vb95P3SjXY8b7ygVYZS6wi39O3v+R72HrMEVI8LPMAOx2qWXfRxNJfN/
IUQ++H5mZBN3IfimDgxS9bGfSE8pgA0fc14iSsUPFC34ROWpiqSqtAfefM2T8PWT+nsSrtiQC9uX
5ymn5vLqY1r8fF9iX9wQbbsxNNiGpSJz+9+LGShsRazqgzOBEVWt0pYiCUMZCdDPVC0c31Mn6j4E
W22xGHM6uz3I9bWx4Sum2Aw/zOm75W5OgHGWhUCVgJ229bpoCs9CHcOTwkuYTif9aKHK8qbfVnH5
aLi8UcowX/+Y1H9hniYpRnWt72Dw9X/T609FaAfL71HF3ieNh/x0tw83cDbu/bZpZPMQa4pIp8YU
DXmK+lieX9JRCnr5wwmZTDg751TgeZSje5jSXOEDkdxhjdwi3rTZAWALKSlp7P2hV8jGzyu+cOT4
x5wRdOa7OsO3T5Zv7FeywIhZhySqT/roTK2q/XcFJlURBpNPWIfXeNqpmoz2zHM2i1tBJAZFDXn7
qokKVsmf82e4samCw2HQaGgtNc1VK7HvurL53g2QHIwy5c2dRNpoTylxRlBhB5AMjkls5Plziq3X
zz45tkEMN8AWHU1xafsff1ftvpTY4BPWiZzuc+p2BHkHj+HNASdZt5gkRkDPYlT0+PlMS2BeQgOG
mfRX6Utb9Ji7mdbBs2pk9DJCxfg70oQYLzNMFSRiswXZuUtN0JrMIkbjfBA033u3Dg4H0q+W8q3W
Wg4wOWi9OUEIcoR0yz6tCx4KwA4EIeNxbXRvVIQqHwkz1MJewVhY31WS8CjIQmIx/KxUDxeSr7ch
LVtXzVmjpw6TAzO4P7XCVTspYkB3RnbDrGCuSCBsxAISavf+vLaVw551fNoYNcpOLru7hTCRs5la
+GWh1+PmYEFZ7XDvAzx4GKSa4s3uwbFFMcJ+Tpe4nJhLewaw/tXn4kFWcFU/7R9C+z+/6+94eW6M
0S9pJN056Pm/hqqDHBzTk6AIaG4fVyAUUrtMK4E8jFmYM1O8T6wvT2jR3k9dSDeGbEhSU+5gafcV
lqoGin9O646LAHELmPFUE6qlLuFp2gcnubItqhxTPWyR4a9sdg406lSLESIJjJej9M+PuGZ8HC24
K0g4zP8bK6B4GxfyW0vsy7yjlvBioolYmQSfr2iylsArGTE0juwDkMUp5SOTwNEcQIMATKbMhPS9
qGmjmEJTWmqlQQLVWMm6IMPkzt1eoffvkr8QP63KtR2+mCinxuiyM6AqvzNCnEBQHsCwi0Ik3RA5
K3xdABBbnpiz2WNZxYqZ9q8/Xqp9W4nutUPXHbWEK9mNdlw7VGj8k7EVngmK34kaxPd7arqSwkYA
L01t+7u9bC0JQWitmPMlghHNapCzLPNCX9wuaj0+HopopVjU330wmx0D5nA14skqevnlkFSlauSf
Dv/+/n2AnUYyE9XPVhVpeTGHO66xS2vyNjrkFWDvrSkTyPzV+V/n7GUTHQFuQdqbBor2vWPj9ob7
OAuJRdIjeO+2jgQqkA1Jd1kYcfmqzRZGqUMsYgNm/KsQOnDvyfqQf+LjIz/jR4DvUEiR0BR7dIiy
Gv1y3jKOFyG0oSDyFBuU1sGUXshQHJ1mxbb4Wm1cTo5Ir0MVgUvlAmuVF8Hxk1KgeNRBl6ApM7Y8
lMUfrztGHVMCuBdHM9b9ikr1Trzmi1u+tXLJrwQPrQ6irE3ve7B+BtUKAEPM68LR0CoUgmFsGrHb
1FDu7j3WSXuanQT1A+MmdVZS++o9l4PfR4GpJXXXVER7OavSdyRo29CRRSmK6QZa+shQTO0EvziC
qcXiULAUfUwmB0C23fVPcBuEJ3lq8qm9v6EKey479VFMjRV9HVUzC8tWTWasnZGiQBcrklChXh0Y
d/RJvKJ48rgSsXVElNBUR5d5K6KcKheWk/wZInLgAC4k6iUOX3YkgDCQLEhBXbVx9tC3QFH0F/3f
STkNcTgqh7rRIHdR/qTaqMIvnoxbbYbUC8Y3zNv6lKsryNgN2v4t7EtU2ebsRKvG6Q8UEbVgKq61
QEbew3FIdvinYpVentTYrRme/a0PBYwEyc8vocaxAYE03DFux1FG/l2ihgXOiZ6viXAIF55dE88w
TWaTyZuec2nLUJ9nzJjodRsldxPmNE20RNtgEKyvGYT13gx+8R8jggOOV7kHBVuXnmgJbj67pSHK
GVw44n2fHAaiUoxGTI2QebgDpBXKcys8DXYMqJBVhehdTOIzgfNnG8gkVBJfJ8nWrEwxcZ6wHrbP
3cYEVZrJh5S/KcTGyR+Ma2R+bJZqCHWvidkwCRhv/eSPGxyy1CCrXVjd75nZqSzh8nGLYkYSjeBh
0djZ07TutGgPpAzB+7Uq2cjrbVeihQlR3Mxt2hYbUBG2p/IYckPnTclCnh2CpQUU3wPyb+rX117b
wFViSPG3ckwl44B4ZgxBPsi41XzoO+3mXNVyk8o1Q3YZcTfIxapTscRri9vzfymrNr6A4jOnAU00
nTmljufk+bqPRe2FKnzjls9tbgS5SpLmAl12c3blb13wy95i/diFncB7Z88AryAIdVjvKmsc2rSe
IAO5QB3WjN5NGr9mho64HhkIqSSY1kTFAggXOfRo0/pkvd0pOhZlnhp47x3nNKj+z0Mpp4vw7rsL
993/65lioZ7vnVuE9dBQaPmEyPvjMz1YtNfmcbZvfrjRaTBjluungKNEmfFBLKulxEhul8PcA7P9
BO0MD2M6S6SQXSuiugOZCJjW0C60ib2nQR8I5dhiXQoeCTk6gMuMshum0T2nr9TdaRb8kxCdtKbZ
WKIW4U/zKwW+LmUBRFAVXrHjAWw+tHobf73xTlx5AWJILutkwF5QfnEfEd9Arjz/TIlagqFk4ynO
20yN7bl7WsXzqx2XIZpXYSJR9Djgh4x/IYO4HVX6zDi4fbG/jOJdlbRLtJ8MiV7fIKLizie2pQm5
5xwEfRn2/t3vxpCURJu69dqtUH5J5dcVEfRJ5Tn+C77+SwiCUR+xVWIe8d3zQJT+tdJ0CizUiUwM
rAvgfMSogPeUO4oToK0vR1iLIxos7dqAA7nQi388hpPk9kCQDTUXYpY+GZxREDnEKZjlzrq559B/
CbZTcJRnpUfZRiwF/KmW1GYxaqNdbYebaqdqK92SDK7SImvUWydlltCDVlXBpM3LIaksBegsM4mc
IaVNTkkAOO8AtV7kUfW8S4MFCbiHj635aPbxkUB2qGuG4LVgLM61kScd51+LTw3LRiLescxxMW9p
T8Ghfl1lMuRzbv1DOlyIkRHwyPKtdREaU/OFyRrS3KHN+G4nHywxQ64GV+/4MkJPtFzADJOf6Va6
SFKbz1ABXfc5oUUgrM+mNnkFFqk1Ji0J64yIeZ4xvsIaRSpCwxIZCFmo1rMH8DkoNvdgaTov5Wee
CinL++KQNEfvzS7OENXA22B1lBYhFGoMa0B3EjduPZiHJvvAw4FAwhg2FUYORWyILzHuxYn723OC
slkGvwtz38HE7IYGdQwD35BbUlGgzR3vPaZCwPp2YkaOJ/Ajp52pjqxCYSB/m5mKDU95FON/31jg
M0SDZAnLCJv2Mdy3CM9TCFZbcwXbSAlWXY4135Vw+2SE+s6sjG97L0Si/DpltOSD6WsI+BkUmvpw
Ccus8SxJNr7PnSBQZWCuK06H5HxGRe+DjCjkOjfYPmdYmTYWf7L/hSvs/qiOKnqDjAkYIf9Gy8Ch
/ppF+MW+m3Ud6uxoPSOG2a9PpMW5onBDhRBNzwAbvW3EmqmjpIsOga0FBp3AVlJQqDbrM10ZsJZg
a8ZZw4VkD510UPSl5boKpOiy8TvmyAYXl19Z9sjDO+nSQQwVVjbLPVBanR9AoBTp1tzEyUnpoUnv
ZyYB/06CeC0uOK/M/gcQ6wSCiFNviJ3NZWIKjlvY97ggdl1UHsfRj5yL9NQkwmTmEtwp+UdEm81a
1M9FdvxblhOpItbL0fgSL4/fpISEkeobD1dEEBE2XhgiQmiXJ3I335Bk2glFMAauFIC/kSa2NyZB
UPSgm8gzgdC7f4ZtzCraQ1pr6eDbUMfpvWAKhMfiG93ZKeiT8F/gYpJEFvRRWpY4MdXggsjoLaYo
BzLDJaSjc3Ih8Ty559menE1+KlghQNAT2dmPBbu1f/MuhwaDvM8spXLplge8/ZMyDfce6u1+s05+
Jj6790Bt3e755v733Q1yqP3VUeDi1hgpvMDWSyU0XMhZimnGGCjo1aPBLpyNPZuUjhffuUf+XX2k
oU+AqYa+lo4T0XHPfcqQUYpguR1zaZzYf/n8RGR64xEOOI0tsTI1bUBXrELm6UXfVBXSNfwdRGeH
oepmXZrsQfi16nSQzbQ34AfmOVQuSEfbcAdKRyI+CuH3ACu4u2rI2XTUiTpqgrsa9yYhx22y4aH+
Uv2B0bbQj96NB+wQ2qyM/05ZbAygJjHojoxYDXn+PtSh/GrI00hSQlTMMfRL+NNsUb6aNw2gr/Ei
/2nK9Ko7B+avckCQZ/vs0FG75aHZkpwLqmGy3LsGzf33Li8pCwCrzCKmHADvZ5QyoqjO7rTOZquA
U7+TRGZD78XIzbO+srKPEL+zV6NsWKNVX+UOVT3Dm+doQdS6JF+P6zDvcprqe2bBmzhhbA/jB4ih
J/24IqDYrXNStZ5VMFpSITBeTc8fTyQh22XSgm7g/dgdz/Opl37Yfnh5/UV6A+eiFAet02DiVQwc
3hspJuSxau1jK2YfH3PN31bPHU19DYl82x4kWTmZEnQk/3GVTe7mObvrRunPMZlNEebbjD9KmLr3
kYFmDdDJDWMcTXwNnFWv9b9L/aIfGCRiREH9UIlEkVZGi4m6TGQTZ5vefdt3omgAsQhJZhEEwUzl
b8SY4TdsV2P9ydAtO4uhBdXL4z9PLv+qqzV/v2BEu5bx6Vu2UYt8XAC9wSsmaaI52AwHtJSKB62T
nvupnFkVi7sFwsBeVVcswecdho7CaLiS3bRg0Y15gMiv7BnazzD4lbIYSK8atuWjo/jYM0hbTIT+
VOVm1x0QI6PM7te+EVGVpGdQH1tcm5OwUyZirJE+6aO+lqQfdQCcF7vEkZ6GQDgz/Xak1LchDCPt
94oIYPVtsCtjHAVlShGcseWpMYMINu2GKD7ndxo8iztavEaraHHqMVL5mu2rM6SO9LzeUvDgKCD+
osoMpShxK4oF/W8dyd4rMAkANWUb+BuACU4GYmuZLxpraYAlmaZh6jakuPDqrCE8PBtQzrm7jPqM
z5zfwewZ+P+xNjM4BE8C0l6TC/oBGbFnu9958jSlanyL8QU+gseYq5+yCo0wyT4vxvx2YHPnFY/J
pk1rkwE6i68GJyLJ84AG0O1Ct7ASfa6pr0KVMo9dtWbkLdBg3ZFxUFBODE279ziq+g+xTNoBNsuU
Q5zXhc49mCZXEjBmXZVoQm1nZLg7+KtzVI2/0wGAYmTagjGNcbDTYExlDzZBTJLDTOD+uZsyPlsy
AyGzdti2+p1TIKMOU1BNvZdVL6Hx+OZNrNqfxkfYkT5ZXf4WBKtlC3nYEdc8OcGjie281aW9+RtN
zSSRyXOzLoM/tDkocYG9ZN9EEqlczBmRXiV7GRLulOeH0YSShehgQRzfU1Xj/CzuQbrG8e8q6z9Y
y+BHMu1wTTg5zMnl9fwIpNrWrZ3VJvtlIPaEDrpP8GdMtwOEC1uiuT/x9nrkvwQqjUfDL26lw2bl
zsjYiAG0e3MCDP2AJt1fRU43Ei4IsGOPCe6Ait/HAb9C74CXhTQg08jZMCAXs3AO6Bd2SkvOjlVR
6m4zarf6ePhGUiau8WvJjQoKt/CbwrBqIHYWbEKr+F5QkdjqKfR0aS7MNO0HTRsJzdwRnxDWJT5k
zKLIYpZUG1ojGactCb18RuS/fkENd5E+WDHNGNGVWmQ7pbQD8yn+7YDl4NF+W9seEHDJ48CJXJGY
0OPkdXGp4Fm+8s6O5vgF9SQQ991A1pxkNnxiBMEZH+VbVXRae1lUC31cuWudtygNSsk8QK5CF+Ub
6SixIo843ctqz5t4P77U5eKUjEFrAOTcJbKPnuouYHdJPgJ/6Z5qaDPvE08CclTvlihB9GO1iNcw
Xf/OyiBCSa+L2VhjBmZzyX97uKB7H3KBNkp6rKJ+jLlROulZe6EpiQNvpvfEJyOA6KAKYBdZ/r42
kztQiCk5sW+M6yEIPLokPMqnPpBkwRFvZtFBzlh12pSxHs7KfZU9PMTxzUM2tS/f9e+aCyuRIutM
VizOCJj91IdNUgF9GyDqnkJDlm2vyO1k0S6TMpMQbyiwzNSyMvGVAZGUiE0Y+NLKZvoHZk5xI3nq
oEk3qFqRbBGTLwH8GtE3lr4WNxud6fgPOtn8a9Y0PhzFgLpioNL5UfHZzQ1mxai4HOvwVPPCzIbS
7wVZHPB92jRK9ciiNU/Kwte7vIzMep5S3LBEAbHFJHM0f+4Q+iE1EbrrFNsLdld9yy1EanQvPv93
R0zpIyDWb8PbRlyy2+MgtzIYshLdCabMlCGO9pUQKs7b/WTOBItMkRt1Wt3TYm53IEYlbXCdCCCV
TTn0pU5UKjXYlxsKgoQf7m/GtU5NgplbS3siT2HN7WAziTvohVrKesGTGtGZ6hzhOrlmljudVzgd
l0jm6hicwRHN91Z1Eg+lxeFUtaXilerCMRoDqeD+myWviPewgvl2mwWi+r0UP9mSbEvmjdSyElQr
GHP2VKaE+o82qQsi5QMaXW5918zUmiURsRC0cZ0irFcK7hZ9yZXdKlsKlItjQkTkM0MKgC6Yvltx
yZB3dV47Nr/Hj1K5TW2/WP+IW6R/M/TTGnnTxs+/9HBdlwc6wSE8zoUMRqJt6hpBLmsOhsSX5jHG
cbXYmdYEAfhoJMKofNEBJ2lh68Y8hV/IzYWeCf6eM4+Hpz5DfIqU1Ugj6mL7GRtLyHB61g/0cW8V
WEYrog/8u4BWjT0Yu3g74t0faaw4ivIe5uG/XPbdCz1Bi7+uxuSrjHsYKK4a236kFrUREowdrqC0
7rSGqSdX3qKQYStnuuuD88mD29pD5uUVw4gFF+uBWvfHa8R8qwI2M195qHEFrssQzOWkQ1Vzf90J
ZNWO1HxXOHeRKLi+HwLZ4iQWC0mouiuLpNlDPipR70cRWr61bS1PJfVQw444xsGi+staMb57rZX2
lKD7iaUXTQLfQ18ntOdCPfVXoDrV/ac/SoJOcL1/HRRK+2GgV5qAhk1adJ1RrCwCiQkUUEqahcDD
c1a75a31VR7ukuEVI3boux8LfBp8e7Tufdi43SjVeAYqt9bPCl+RtaLs8rEMupS6ZmBsDOKB/1Ha
PGFMZNpswVbgoQgeJ61uE9FOjEldKIqk4wj9kO84ljGaXn/FFu4wV96pGRcfntm615DvVZFcpmtC
BIO8fGBidC/Mi/lwuIk8hEcMZkYQTjcol/5fpvxIiO+4YE2hzpLA7pnReW0r5uBtZ6oh9STOIyRn
27qrIk+m2NLUouwPlKvAqBGeDGyo9Qvp4urR0RM65wh8abupX/hoJf3kW68/0AsgW5ElJpgxTrVT
8mdo1+sW7Ki6ONuZyI/ccRfDXqUrbP+T0XQe1xOs1ozfxwwoNc3M/MzIg7OzQZgAAwcS5obWMzxG
2NJ/vT3ZNdmH9mZ3eQDYwmkjxb+BTRScjh2VNOR0Dyf9fkZiMQJZ7s13DVsJyPmxJs/tssI1YRz0
DRtIzDmVaUx8hnmLCDZXjzgUq4XJZ/R7MFwEZwCY3XtbK+BdgQKfFMRgejHGK/7p39QW9YZk1hdm
QY5nio5mK6EzAgOVBOeVNSQKNus21onRfzVsSkTJZWLISPb4d2JHXTFTCUFLeFaa0kCSBQp0Lxuu
Qj3XKf8Grf6koiqDyxlRZxfN7jM2Kk1g73xU2hWwKj1uZ502iHORz5QgTFj4vWLYjM7ytpUFXPYf
2MT6h50mt+BGQltadcl77PnNJ5TvjgKJpdGmZClhKs8nYCbPdB94rCFL90s/0KgsfMs8p71v2lPV
E2aYC1CB/ra+3mEedavJ4iQ11hULaLp1oZXs93PUqJ06Dx2qYu3LAPbZ5SxCiCYLlvmE7rQcwjob
6Y/wYBi6M8FHp2/HO9uDjkBgmEQymreMJuqAjwWrVk59mNcmeqR+OSv437axpiyl3IdlC1cHjGzi
vyoAnl3tJV1nQZj3OKEdq+g3WdQ18xn9pYMEt89u0ugnf3p5huxhaU9/LMd4mZSiXrz8tk+RL4Tu
/4siSN8KP708BUTqouivoEMyRRHSXkxgLHwPIRLUrMbNqNyNOWIB2581TC3F8JRXYC8pVRcnR8jJ
RjiKtKwSefPmDu3LveoI++71rpWDxpXgkIgzJ4pwKk8zEoeDD8EN/GJm6Cj57wVR8a6z7fINSh53
Km/xdFDEHSslP5Ky3U7hQSbxhOdPcwzLAeR0DDGv84axZayuUm0t1gWeFaQJKIZH2rK/wXy51MF2
uIbt/aFohw5fjjLvfm6Av4blwJkvA8sEgDNBzvgp6k2XFYS9CTRldd/w2rnD3egMZ2eNWwczL9cD
R+5UBt0qc2HGZjTjNJ9w5qdLovegYAVlR+5MK7I0UbDVvmjeqSf1JAUQ5+79UjRcCBTYEiuuuqfE
sMUUcPGQijqxzH/Az216M5QLT+paJ7U7TUDvXF0WmwgTyJPXjsfeTHBiP9nfcvrzvzAZUYhLsB61
8ny1BXL0plFaLslsF0P6NeIZZuTSV5E0zc+IX43Ax18UUjk4i1O5KKW1EqMwXh9UsFHDuT+/6q4K
U950yYfJ31EJ74CcPNtet1Rz5PVQcvjgIsU/85S36XrT8XDzWLUkIxbSg3T0wCukoex3GEwPzWCZ
dwULQVbUKfxwx2Khx1wx8LBmDpyRzjtUmWkUKNY5ALhoNFeIY5q9tkbVYJC/g3otT6BQpyqqjWZq
TBZ/GXrCATXunGR9zvxO05AK4kDBARh6+U2A3p3a8V82Q0xFIa6/fmrhDHiw3LE1A/MiJ6um4o6J
GRX8/MFAOAROFPuV2bQ+QNSb5aY8cI5PGG91cU32JxqIVOMg6mAhUxxT8T4iFowDVuTw6WtKhxk1
BI0u5J6NVLHvp2S5bg9A/MXww263wjGxA2bSAXUOF8M9fy2Te0JxA7N0WibRq9NbzVT/014p9jco
AXBZXz1oQOmd1SGBPiaDhFBnanAQpNX4aN6Ev1pXcT1hk8ljIfojOUAcJRXfrKOXQHRQxBzl6/fl
7VshKBiA4sECIrPbaL1Nr8+xLZrv5xD5xe6hox6VeaZT5aA+VswXtPCnSIL/+w21fNhxCLIGYKUC
11ME3pNUJCyE45zh+vjgmt88vukh+7Rw0zPamgeUbBCyLwpcvXDy8WJHPuh3zQAgYgPXhgZRhSPf
riBI+zMsmmFmQyDqt08l+YXPj70VRllQor6qzxoE1ZX6wqP4gH2lTrcBbz57soCyGYYkKQaHGCdP
tX2q8z03VH/lzAjEbC6s/Yu0Vygm72gdOQzv2X4B0YY/Op7EQL5Vhc4lDUH9PwVzFf+LigcWG6cs
FG50vNtOSPMmfMx2b5wOTR+NpFIKPJ+VfkcYyATAElfba8cyX0IRgu8G6cn7wtwGv20mujDyk8DG
I5XspjB7kD8W8rOeFgiDoF3WGTwQukNnQWQYeGCJWuzq1N4UudWSiGWZqeo9iaBvGjieXhvAOfo0
kdoioSxIzuB3Y8WKXpdJMm1avZ9/WL5TYOJa3P+M6Ko6eQwiccwyGCj41b0QsId373EkmbhErxS6
meMOzqNAHadd/xinqNloH51y6H9D8DSU9Zo6Gvq/eNdiztdk0/W2/lLeVgzErIFdo+MXlMvO2KG+
XkLYpMlEqMOE0hLg24FiKJjwvqAG9P2FdLi3RHhsMg9wey/oTKAn39ZFeEHCRrsiwCfOYVHe8/ST
tLsFzHXylmSdgsLCVbtml2I2j9hD5IcsvPc7ef+2lrwRptPNHS77CQkXqJH8Bk0xw66O0XTaMRXE
0v7mJPpr+3ioXVeh6cJ/POJQQFsgDBpJYErkCu9lbhTrJ51jLy0wZGH+PpFPJ15mJ2CyNDjIouCl
B6jXEE3ZSPhqq/Y69Gr4fVUtGkcSKCUsXvkgvmjtJ1glx9EHQ0d/t+sI6zYs5bZ+p8Vl3G0a6v14
Dl/FGNeLwMWK15sDaheyfj2TlYboRNzfzsfZUqo+ij1JvlwSPcln2jlg1VYZ5TbYxjVAZJjUQ9p5
ImBF+yHWz5ut3eMFILvdIkSDQjSwzf9joz0igxnATEvgZ7Mv0REcs8XYnlOMAckYXL1vHruYraQ8
cfDR8tXu063S1nHBFNL1H5cJ87mHZQGtJlMV7jfkAFhLh0ZOV61AioExUqimtzu7Y8YAzzlFdpEV
iXxinwhuXQunj38XqhWQDRXcUTwvqm7OHukcNCcdGnLH6oLABF2svK7iqTi1A2x8VZ9h/C6Wk4j4
u5Yy6iHvclPRsNi7GUVNUahre73SpAzaEoFeHOQrjeQLBbTwSBY1/8koyOymG8goS4q8s/KdeRhR
t9J3e5d2pLaBnItC27aDByuZ4HiIRbajYILrwEd+gJ9WNHZDaf7+TZup4pj/gnjRmP5vbmFpcVRi
KQa6Z30Hf0tKTztL+K/KDl1r2AweH8KL0pRA6B6sEu297rokfcO/FcH9wo1K2TO4lwSPgEpHMoxb
x0ZO7LvC+E83QMfkMIDbUMytIfs2/hPNeXlN8nYVGfqN4Pi+RVhjwiwkAzK1mXxQN8R4yprVCkfy
ERoIrxv47XE3OcX8AVldcXMfB14MeG1kxa1WPC6UWszyaD4e1aDAUNOS6kk4LEg1iHt7hfg7gaw8
pT8rwk7PsyQWu9d3pLMsHaBgq9wO/1ZkU5EZcUKbq708QqIl48q9qzbGY0KfdIeWSyzLJ9llm/nA
WCjzrADQODwbgs/K4wWf9DfX3YgEyIlM6xK7pr1FNsavwrlRKwxdErcF1qlkqZleAdef9hq13gYa
qTZrTRbc7wsJFt/zXrga/cIjL4Xp9hSzfpq5wC7LTQxtQHBC/jRF4eeZI6L+ParQ/t2XmCIdyEOR
NswUppn5aEl59LcfCwthORUVLy1EzoYUsl7/AYx+X9WhE8MrQCxcJH1J/WQdftXvIPA/s6A1VGEh
cchpt0b0mx1dP7xG2HrJqTseX0IHzDhW7/PfLE2+jS5U7tnOMZ4mQSBEqtQTBaAaZP5f43evSI4H
AF9niBhiYyPuDds43eQLLIKtyuapp8cCgl359idKy35OLw0ch/+/tJAopgvrOuYZVg4/D3EZSLPL
7Vc3WAPj/KEfTwM2N0T4m4F/WLzEn4Naoz+eu1x5CZLAwDXMxX0a5Ov0WJYAWr0oVjo20MpEbtV9
v6n33G/FSMv0+zGO6sTW8ryjx8rAQ9O6UKvEV1fAyTl1nXI6rAsvCNWyFMGBF1IzbCrN56sqmrFG
drtJdMefXFmTzmTlu6lI8/LqFe1P7Nvf1lIKzysfM9P121Pnp2M+G1YLYxVapXgx51V2nhBpeIDg
FRQgoisHD5EsB/idssZtLINwnlyxbFeYHlnO93ZYcm5TnNgrV+vsiMqlHCd91qp0yRlJteginDf3
QYtPv8AQ9bIuJf+7s2EUFlbCS3K3PEceFnAqEIxwWIQmfkmGorBv+/wWCYmby6Ev6k8qrImAzcbn
NbLEcVlZMOXqONqnNGgihgcVIwYVG+PXmNIyUrRFNAYIW+vK5F6U6Hf1dzFe3omxJRz58D9orWU6
jv9HM3n84iBPkb/2Nn2IOZCFT+FYA+Ux5iNYNbHJHHT0AXPwVPjjSiqTpAh1lJJ4Q1v/R2YkLqOb
bxlw7kGkWsiViX0c3ueeTUao1/b1wnfYuigccHetWdk2uypLqATs3c2cFaSJGSPxxr9lNYARyS/y
Se/Z+Td+6JNZtDmGZIfU3HrCwoo+xvlLuVQ71tVN8Rdih7SRuTYZ3qRLf47HoN3EH39XbuA+3v/Z
aQW63tI5e54W2aqeEkO6N8yRFhFORrHLydSNDzEdM4RVv0VcVlV/0rXz5Hnsxydyouiz33r7BUfr
l9sO7Olw7KDqGrAb7itRuETy2+d2Tn8nImPDLHDkiqeX4fJRYJXdJStzP+Tx+M/I4K/ftEoG2dGM
K3vgWH2E0QuRxbt1hARDt3ptaaCaOl/zzKnG2UiwR8cMBEiQK3eqpSCsCpjqG0PoYixkYT5laWFB
UoJsvYpDIDjxVJmcNcmrtCMHXcBKMSMXrFigAVRvVbbyVC97cKAHrQqPQGr/YSNKHA7ICDiDRemM
5EDyw66lIXwVRT09WNmUA++atcUOsZRfv//5y1FAl1oag1sPI8aVbn6YZ61nT9Uikn2yotjSQV19
/tt0Vuu78lqN5wq2lIaa+JdyzHQqGdPrxw5HCVmW1y7q1G9BdDCUQM5hgBD/O5rT+7ZiVygtkWBx
9S7DmhGiFOuBF3NJg4ohZOpdmBICJsqRHSG3OSKJDz8QdiMQKen8ITRjzKvTXSDDH5b82Eof8giZ
x7N4ZGyPAcy75jEugehvalBJ2RgWJ2D/+xrycT9ARvsSoLkeY4HK8sWVy5ZMzivjKo/P+xmnWgIr
NG+Y34R1dfO2Uxb9eLPgL9h8WVctDRydfn/Cmft+YOs86njNGJUrHVvesK+/R/x3B7yYPqokuSVV
CGRxOwDD3ZLYkmAiheN5qWMnwVtIcKF6AGxYH0MZwWldahfVddePu1PH/B8qf43S9/wmE87+mLpi
n0CO84fkEo67oF0Mpu7BbP26mHpDmiT36uirDmn+PU3MNWd19bU8GGbNtOW+00HatqIU+xlxSeh1
WNT1ylBey6Pq5z+P30P7lip75QAYaFRoKr/9Mb5FvQGZiD51m8vTuTWQnAFkVDK91XhdlaYLhXw+
jzhCch+TCjFngRMoYyo0snR/zyk4V7zf79D8JQpY//ffosHghev647TbKRhR56187JnJ/Zgo+lgT
iG2R73IlzYZjrZ934RRSOWXl7hdLozBC5usjT4t+EuOTfylE0EBZ1DVWCQ7bqJ+EzDVLNLtnIqJl
BA0xELI0OJiJ1nv7e8CayFZUjZgV1FljdZw5O3fz8N5iUSLuGXJTxinikSKGV0lutiDPv6YlWFX9
DpA2v3c0czXeqVd322yKwdyeG/BUC+UWjAMFdqfVe+9MXsVW/DsRTFQ+ruokceRG0z7pDFYupEtN
CsaUsQ+bnBZod+zaUj81ID8pYLZGr5grtWuC+Rs9zX9qquIhKo+O8ExTZgCAFIWkoJNydpN2RVz7
DUzjwywQnXffaWv1LkTkaNikRVaTeqGhVhODO8AGy6oi0kgNDLeyzR28wkOoJgwiUbxyN7SmrYyM
HP9A1thKVgVOJRJI5n646ccNLF6cqNC8oPfh+diB+rmoqW6qJRCgdHqCYqWBdry1kYB3v24TT2Va
NPPI4KLrtyN/dwPt8cle/AWjpM9nBrNED1v422lOt9jIaKg0rpH8GMjVvj+nOD8MuO5sFVKewLPe
9ecl+uDFHD5ongVn4jb0RXKPEaKlbDDAuf6MEzV6W8jwJiisNdZaatZuOkDdnSTiKLWGoj11W6+S
LvguZlaepsunNtuW48D7fcU/XnTGNg/C0q6z/UuXi13fVa3t8qGgc5tkSdmgRcwXAPiaIpKhmOei
lz7VE0q6e6AeEq8GAjm4ukCw1hb1iXFUlxnZ4MteuzUk1Uy+3iAnZd8WpcLK9TgH9jzqdp8Irv2H
W4miRvfAza6+UdIvq2aCyRgkyrTFzLaqDz/ChOM45qJk3Zk7kupW9pe/5xZGQuUTLPhDKb+JOjAV
jYTFWGJgY58GBFZjfmYr+dqvnZ4tWDGQRdmTWjh9JBp0I0/3NKtGoFgpJoW1beNCHhW18AEzZvtn
roYfVVwpKwtL75Hk8EqvihQLXmomrcdXdHlBSWQTEtJw0/op4tkz2yKH+VB8wQbLYC7BrKTeIxNx
WWYHn1DKHb+KPrFxGpkEMNQbZ96E7aHOxKVBQ7kFQhoh72c3IMfyWsCL4BHhW4Q5iUcuHF3FX+ze
31WEnCtK4i5WPL+MOR+jSXsa2ZCFIUmv2yyhA5+yOcUVtGoOShqoQxZCiaQztwzoi7W/fOfvnv/T
xcL30wHumnkGHNwBxTT/bU/y6WVBPfonfpTszbQeDkYaW33WJKUtPDRWsO4KfP5iAoRuG8G4pzqm
6oXI58qysMiHBDKqVOQlTKmYigakapsSvThBwL8/cZqAO9W9F4zwM2In4QZrc5En6HDVRW93t0xB
kraWTGDeVj1FVRm4nZ9zwymJDiLdk3v1WTWYpuvyB+adaxryBiEDdSD8pdNtwQuoSB6YjxMvRUWq
4lgEKQ/DZkpHCZ8/LMK5vd9WF+PjYb0x5tbmGHfjDZ7H9x7YT6B1KPKl6EmHVD2o0siS7olq8u1C
WeR3NRmF3bfn1+TN/AN4kzlLDgHTNvroI6lPHD7kEYfPiUBQDm25+xVxYOFtXw1nEaSS6YxlyaqR
fKo5W2dVPAIXWzqmOmEfTJVR3g7arjbwGshb6NBhcmWFLsJuDjHtgV0KDSDS+0BBwG1vjgp2ikGT
JZziqxNE96reiz9qjqGPEk4wT8NQrTp2zBGMoYgRXMraqVlejzW3UPi1QzjDm6c1sXo6f3KMjEkK
L7mo9WFjNeS2xJrL4UVge+X5nGo+vjUAIu5AU452gC1ubPiIyNqDLLpuB6FXcF7xvMa7b8ZkFsbx
4ZTL7IqneLYEbAJPQU/1jL6dVSXckk+yl7tHEM/6nBJMTxyW21VkahNUaS8MuESJHsAk8RQEm07l
zn6YBKP26hh7cnvGWDR4gjPvrKH11sFstkP82TvxLt5UNs+CEhKB2MHUZh7NzQC81fuv481b3Gja
SPROjMy23/SnP7S+0QIRYLlHaBUgrU2IQXkQVs5qRrNgsYn8PIQNz1ETYy/wqvjwGd+IMZFnIHdu
G547bj4DsRUEhHFgVgVw+K61IF/+VrFxOnMDEaGiq4xTD+xzVloBtD3a918QU45qIL+pbMM2Yh/b
ArsfuNApWSitgIlSV5DsEL2oUFPj50vXojZ2amsGOdq8jxfySbbdBPNKl+KwdkhtbGZ+9nzwQZzR
x/BDlFUeIYwfLNuSsxBxXIDyLLSctzvdKU2gvH/L5ojqA3tq0u9FLUJen1JcbNAvZxPY1RPWalHf
j37l6z4nP6jry15E6JhfWui9Ivjj5nU3NNV4CxfwHFYOOHiDEg4N9JhmR34CHkpHxc2mlHXn1duJ
+4yPo3ot2r9C3HBqO5OBwYnnAHMIzrhND34NGLs7uARti5jtJ0EspyguYrvyrwWryG+9q5mp8SRm
OWubEu8DFu3XruWuvNHxQzrCeDoxpmj8F4M9v/k4JY/VWQFhei+n61DbFYiKIY7wgP7dLQ9eWyKA
WfY1OvV7DKgIAEQBSMrIx+AYdmfodQBz1gKPtJOAMCct3Xz8pGXJ8mvXn+hljEePzkaQ2MupNl//
6I9l6hGsT+janIpC+wdF+YyagPKcIGHnopQY+I/xuKHO0eeoUoPSl2cFvVdLM7UruXGyGgQwbIWv
3ccPepuI7yg2uoO6eUE2LJu8BVNiPt7Dy42Y7B6ewCDqy4OAz6FkSAdBWBt/JJo1nTC83B9RFe28
1G1MAWHo6m3um8TJL02vtizuJO2P4/mtmFyYDrkbGDWQTPRl9AITeesdA7JEEgMYryF0rubpLDCs
63Xf1gg+noRllxglr97znCophe97AebO5TdB5DQ4TrirB7rhS0vyoenneT+Hl8+4fq27/0dMQCvq
bc1wL2OAFHymucHzjj/g48IMaS6i0OTCGLI3kX0VRHVSC3TeAWJJO4TxJwc3kvtgplnY/tl1nhte
woyaNHPxBGzhQNbop39FxhhNXDaivxfnSMd2MugbrpAysB02bJN0x1aCFtG3dOo8akh7CnqTZhSz
XZ1HX3GT1JKqZWwnEiAXsqR7iorGQRApJV2LUYhWRE946oW0gVTJ+ur5sjmRCmaCQGaHcYXvLj/C
MbCaarBBHxWeEgECSCGBubtrjEt6eM/2QS2mF0Ql3LlwXYKYbBwAp4ucxvNTPqlD3T9tbsyD8QCk
U5fA9HetW291WSfczoUDxIgG2xVY5hVTq11iLqRsuxmUwlDIn1GBAJG+dFzhOFX5gDTVGMK+ah45
iyX0MlEEJQ8Zr/b+DDKSe/3nYhBgcDgiU4nG5rzsRcuiE+Kqh42Hw80jRKjXF/S+K+Y/V03nSgmy
6+WuW1xGw7w4d//iQfUnIc+n2sBolNr+I5Kpm6m7nX4lWqBZQysxDnwAM9AjpJl+fDuMRzzNK/t7
aajotZStTigzPHLRczrKfiui5V4Kd6c58FsvWXLRYAc5DePmJQgpRlZPkEyXgdlbcLs+2BAc8SjS
3RfsSOk1XDECcqPW1mEMou59pMv2OyE08OqYEE7ZpGZ/RiJ/XpqQ3f57Ze0ElMgyY/cHezWke5sB
/zypVFlaEi8P0ifflGyqDFuYNVWHE5iiqM+J3NL0kZtrg2W49A6FA5z9R7pn+G3nyCzcPltvbsod
kSvmfNmlo+yDqokVN5HsEyt8pdnGpcwRzH6p/fx6OmeiaekaFO++P2OgCLFKk1z3PmnV20bk/Hj6
NkEzFLAUlzIPLeoq2ayNwnNboEEzsuL1zHipwnRreqtMcbliU1A2VvisBVMWbRl9lWk+i7IRrVE3
lUqsq/NIW/b9/pSbKHtoyWoUQqqWZ+Ds1BnCLbJD4Thoi1ENOrGeJzJk8OmzRZwI08hAdxksia2S
aDxmJ/2QNfm2iAtKaB+y9o6JgrIW/IJv8JxFmVLtRRQI1UMgwZufvnKFL9ysXuR4FIujr3O0JvqU
1kYAkZgt31R4CUUJgz/LawuoY7SDzBa9olKZpiwvamAjtzR7xwQCgevFhvPO0BtlXtEgvdvv4bp7
6ezidU07Dmp83R+/RVTvjOPqO36sFngSRyfMZrq0DFjLGR/B/iPKTPOTJcsYmjujTRYg056uWMMD
YzgPmIci5/y4gtjaEfNzjp8hB8IbmTxWeAERSSWNW2aEcn5TwUeao4jHDSqt7Z1EExDrhGJxLImm
im5DDpbrDfUpmcht/mi7ZFu986CXfBfNsfhIbCjRyGTpm2cc8yqHwEoR4fbl9Ip5oRKIh6Y8yhwu
k4EwGSieNtVQEpJs6ImgD2ChxFz8+MfFPy284n//8Mt8yxHsjiT+wN9eXqGNC53R93bsRrI747+L
M9KmRyQPz65Uu0pWyXsMSwA4LwQExoHLaCEphG5WDOy1frMyIfk1bv2jj9GZ7EOa/CR9UTtz/C7Z
PGtcnib5+BPrMN1fxA/bArtZ+a5SBHRqfzVpuKe6S1uMJ+nFeLU3HeXNFm4kLr9Hq49HsaVcG+ew
+ie4bv6I3Et4ShGlvSBNkgNVRMrlWCXh4ySrF77UPQscOP8lGuk0wFrzfCg6LXS9EyiJ0302C1eI
VzGvmDgooxJNe0sSdOBNz2D9x29V9XfQdeqM3YPm5nc+qzS5ooLyKCv2kQ4lUTNcUfyTnLBv7CQc
FrpnGWoyWnVlM+0pa0TXvNJ+hkoiRTCRTIgN3jYBMl/Yq7LAeC5MzNhtnAJy+aBMAQ8R0fGT6oM1
X2Kb/hWM4XAclv/7U2K1Cd2jbvV6Bc4MpfuzFc0CqpEq9lsjqzsW1DvFs8ck2z/w1wSq4orH6aq3
BELOtz1e0+PhZT3WG+08CUQ4EFgJgWVg9pNTW8aaE/eIFS9L5u4rmGQfJ6brKKZ/GgDaBQ0Zyki5
i1WnCZGMVrn8VFubh8oxg2/UmlVb37tVNlYBjIa2LxRzqZz5NWwUHXgtYXauEB5ee3iy3vSkfpzK
wmyzm74Kfzk9IzppCkNz6rgfST0X+gtdX9UcfGOtMwTHomNaDWpt2HNxa1zpknOrw5Ccvd0hTepb
jN6aDAfmeNCibPvYJczRiCo+STIAlsEN5wWxMWuFCxGTW6hE1nNj76WBZY/zUC5FPCox2x8s1FMo
q+tVeRc/3Vgkplyjp+VfxjLmvrgkUTyRkpTs+9uLWWirCmH1dz/O1xEiPrwowaHoAWQoL0sNPTiN
MnD1rVGE/xY5UE8YE4ZarvB5aThVWoAa2m+ZcXexY35svB3MFDOTn/mZik3R+KNqujrgvn1GpFVB
aX4jwqhPuRi2Mvx16qxDB8zSpTyX85SGbxUtHH993/cQGC8O3ba6I4OBCJpTZ+Y8kvlSzCzL65B9
NVfOKRYDFz4L7ngQXrWL2FmqwGSThG4ZfhH/aPQD/8DZu31bxviTi7Nz+CF70hGLgHRhD7Yv6Gn8
d+L/QG6hRR2n7Y1OIcMc/OzJaeiKgkUc4QGiNYZP0y1Lhsw/ncqF6kKbkuGcF7wS9mj4HDfz2wHU
/9VgKxr1BW8uiP/ccoxJnU1re8r0ZYz72ir4HDZ26hdAof7VfkhmmSiE2axvWfsyOyTIk564fBIO
xsUgOsyQbO0dC51BvsolQMyBeADaEOLS+HE9sq0piFbmuKXYaV83tw8bKxr4Reo2iLhWT5fgKIgf
lwZC1hM6zY2QhNXzDFIDWBHAeZPLuKNDyFcrqb6pNA5/HtuJR1far0ZMd3Ac17hmmVBx0/kU9lyu
1pdKwViUX79mMuska+m6m+sIk8qbUaEk0Yfl5RVnkbVcLYpx3FucyoUu4XRF3PvmYsTPsK8q90Zd
5gFzfL1HuAp+86lqSUU1s3/saX2Fzb7t/PxbDjbCSbiEdHyaCnb/ud0pYDtJYI7QQSOEhDSEgQqg
guitAINslLRqO9fdVGIuZmLV8pjxUqeZXA1DFLJmXjXoaZSNH7bVbVyd/4+Rp11enXrPwgl21B/R
76nVZBxjX7lfownyOIBPMsp6e143/4hNIvApd6nvsgmrMKytyUpdduxwPLXhS2ZCNq+TKMViTz//
yB73p47ODWFLX4zyzwcbcDecbPo9DEUe/TnK7okO1OfzITA8ZSql7pn/hpAq4jAu5FZYc2MZs5gu
Tudj9r74XN22ZXGmFn+srjZrT5gvt79aaS++8k7ql0ktZ1RvIHRr0s/P1fCseOIVqJaLVa1f+FTL
CDn/k4kEtcV8RlVYAc2m6mcUTXZm4BS93qNq0t8jow21DSDJluYukMXtEIW3pRiyKUbrsjt8wXS7
bxJAmq9hMm2E3NfxMkpl6+wx7XYZyTU6rYVFHR/ySZqGN7fz0FBNvZrIFSKOQHUMTsI34etGC9e3
RJSD+Itu2rrGa8kC+JEiKHe+lT3J2Ff1FJXbpBOPYEASdGnRGI1Fy4Fd2FbGhhVSOAGtC90wZRir
QlBbJXDihaMQRfb7kHSalGmmR1g2tCyvcG1n7D0DDCq9tvxVthqV8oX3BpT831w0tcT51/tRtBWi
2QUFw6LMgF+hzZMxhCzYZ9GXT+67ARoD98scqR1oenBVjaCGs+eRimc4I1LQ6JsUIhBstJ+azrHa
uHVjdLkXVq5Gg2DZcLfuF3Lpv6VVTDhhvqs5MLb3WM0M2nciWX4S93aAu0U0H6BdFqLnjqZrVDyc
WNNF6cabhkq8VeGJjaiVFjv90VLCuCuuTyOq/eteW1A8UXCFe9RI7wUFCjv6UfMZVGvqczztpLt8
q5//6idf4X1eUCRZTOmCqKXsK+QB8Z8Suly6x/AZTnOnQO6rCpsUTKcx1uzrDjNSpQ0+vCGe70x2
oKRnb5OPARv+ifXbETewe7LH3YURy+FDnciVKPBbuA7V9uxTX0ozyZxK92ky5VMAigL7zvgaZ+Lf
9LHmlx4LGB8k1l6/a2fcuxJNUDlXcsC33oWUckpzF7EkfJBWrI+a0ftsRDxAj1ld9U1no2rQwq/h
71jQ5BzeGKXbFxJ+kQwVhGrIf3uucbVAnE0v0tJUH7613a964biycf/WepeGHY1K9H0xWxO+yYIz
IhS4na1VZhz9SM06teITMJFr8dKxhiQwMW1y1+cGtNDsDIygZUnioJ+MxDJFnPX3AtxINPgfxxlH
MoO7S3cDXIrhL7ua0DzFNILyMOjZzYp0tgdNiGm9Xi5dkXpnNZQ1GrcOJGxmL0Q29u7WlsbzMmWl
P4+ITZ9Hf3jBcJ4gbUoTSYdXV0bBcgT7VnGNHd+RdP7bijxD2daFebJJGV0yfwVKYF7q0RGMx4im
1J2+eYZIDe0YsHkzoLxgtA7iFCLcxuylGMawF6LMFsqTXxIOnRuuczcQzPjZFXbAYrjn2F5uYc4X
NHaSJ2Pu1rJWKuFMaui6NSBkZyHo+DMltBpdZ+YxXienvGZWr/ammBlJLeu0Zg7FNH3J602PrPRg
lZqlsCebCvTQW//1/tq6Qe8HTS/oHHp+Xk20uoayF3F4kq5v+eDujOCzeNjB3zSznk1Y058zvLPa
mYb8NvCt/tf9mDiUce/ZZTyZWTxVPFTIVPnZvwvDWNGg2J4JXuuJsb3fKyfPJTUNs+18wH6yKOUj
XnkiXNATBqTM9fzya08U/bVZsgro8L6PmNjPdWUGgtgUYC15ECnK+3tlfBmm081o8MsKAI2LsmAe
NBY/4Niq3IlDpME0E85FSH+p0Z57XwDLMnC2N8ke9cs3vf6ZmrlkWleqjQRQaapJndm66iYtECHp
OQxcZIjJt6kxFJ0C6csgCsBiMlz8szEIwBB8/b2mDaBoRiYCrl0iwn93WhbKkJstFkI2GaYbCpyi
9f9DXfKFw6As0kZ+myHQ3fi51Vof+HOVVA5NW00qSFJcOLdQHoZk/6XeI08NK8LF544SSxT+EkWg
Q6JAk4I9vW893ntRN21nWnjMKkfcZq1dev+1tuo6AQnlgZKRd6N/gsMaSuEJ9FZeeieroZ9bSEJK
8coh3sfjYYvYcTFPfm5L2/ZI9+P0VcfxE1ZgRSppyOV2D+E2Lx2/wFR7FCdU9yRh1HKPHwOkYWHt
C4uI1Q0UWM9lMNwg+uAvaArfd3+zECOV+nEBKmCKNfNpL3doVYNiYsT8k80cEEXM7pTda6gE79KG
aIEUpSiXv1vvOpcadpJPiVgjqgasq0/O9vMGQ34x4Lv9RFP7GwSfqsnvgOMNcxDyOplKomsh5UyP
LJLlt9PJyOLQufS1LB0y8ufsR1/4rmksgXgD9I5HEk28kcMWSkQ+ncCd1Exkob4+T26Uh08JNBoK
2XpOJ34t4aFBTrH4+PJP9m3IM3clroFCIGty95yt9cz1KtOqT/z3aIy+T5VyegroXZ0YBD9obRuc
73XK/iEu47P9qZ5nzf/crzgN89ukoIupyuk+AIQCo+3QmFeizdTVjNWC94LFbG0b3nKSTVt19HtA
gua7WTmmfG0meunm76it9jWe27Tqn1hGUOfTzmMULTBYsWEILqoKM+ZZcGk5MCED9IEPV2JsqDdx
wFsfoNJn8kA+FlXbiXokQcDYYo0oOaJtrNdSiZ5URVqMyrpF/0dnmEclFGN3kc/zN4mO2pcYZgwN
9/E/9Lwgs3FE7iW48ku4FVoWsfiqXCIH6mPh4UCgSWO31GSwr1I94hYDKDMtychElO5G79X/4q5J
JinFVGVKN4ilmtBNVyg6C4ye3cdtAHsYIca5uwpxkC4+GG9Of3sgOeKPsXcjWq/MuhlmQNdlztKI
/jp1IH+aGBtcbDfeRNXMqsZAlMRFtfM+qM/mLHkWQBgEL0JPlQF4McjldpFvPfbCFRA0P2QQOpf7
8IAMHInTS5g+Ip3vkccBNHHRRblU6QDEcP0AspCIwJJ+KW64cUrlnNd/SDn8y2dIldiVK+iGh+zp
negFsI72u1GPVtSKIFDBeZDgiojjk3fPvKeIwT3AfWXcpFlyvQ0VdKLq/58znJDS/nvru1kj1e+s
e4ZmKFl07MU6RRuQ4InD8BYDtSdvIy8Y83k6KRjezAoswQB3xK264pf8F0DmH3UYG0pUx0gU8i2Z
n3quIG6gCVUmLGYb8e6rHeN7gPxwYInYvlrMAEJW97wBEB7FWzYCFrVliOPcbULfrZCAyF2hAKUV
znAU+c/w2JRTtnfsYo2Tr3x4Vjxl81S+X9CWmez4B2HMxKWihTcgSVPw2TnlJlaBYiPDsfd8YGtw
QgASgX3EPYzlnSYKAhIWJ7h182lGFEMVBk4FAcN1gBQPFiw6seGKkSIxE/EsXCz4gmmMHKydkzUI
fgPEoBAXq1T1Ye6jXDtcHFq8wY7HaSDxf/dmQFcYmGmZL1kuT1JGOH+BphbA73WI5gvsyNHPasGE
05MZm+gD12e+OzXYCTAMvaD66sN5cxNcETpa1se38Ntji5nmVcS7sEAPhOo6fnDijD+RskYHfp+e
Pm3MhdXhlbnyd2MCJl7VZkR1qUdIvREArTWqzpok7rlIavf6Q7Gv/HKtZW2+QlUw9Yi6cCmAPAE1
p/micu15gUpbYMAG6CzKSvnzWLO5UpElkfVBmupiNhM3x9kAvlgXHUg3mqyK9OaIV+3bLGe5tFdp
Qg0wOPCiAtXC56qzjmp4gXq7wkPFhOcA8gvXTVjuUaDgstHclhxC5ExDB/PgTjC9L4B5XgQedlgz
gGdtCODB9D7IGjcmt6SAjWVLfXw7Hzq17LqvpF3IeI/VdXaJeUiNtj2jeFsnULO6R3buIRsek4bp
LIQXIvhAMmQgzDj7i1K9iIMztznxpW8CaPpsi2YoHynv78wbLHla9wXdGwSb4K7XsHM8Nsn1xnbs
WI2RO7EHb5ZHi/6MKFWabZVJhpqZ8kDdP2vT041UzcWXgY94cLbiqeY+yTp39Brrn821G8d2Ug05
AMSDEQPloDllD56uDJMO9yrLAe7kqh4h+fiFoxBhlU34Iq5kYkYzv8BdkD7HbaYdu9ZianQF1tnM
o8FzGCpIyHAZuOxjrw17u8lGahxpuME6T/a3L9DkWYPAnzCmLpJ2su0Qt+zSDkAA4bfvZZ/uvRoX
/UKW4Y4AQaGQCQFIY4QkCEWjoKcixta166iArzvrw1HwzqG77BJCevqglqu3y03Hyt/gWbmBuLvB
yaC6JRSsh24IgOdqyClamzjOaD3mTrjZB2t21bAE3WhjfcjVi74JerpuW9FzIphIt/9GZ7l1AoKN
rvbSQ0IVLltSmyF+0Pp3H7LdZn85xVpqvejfIw/Eu5eD+ACjOp6g76NNhn+PlZq6N05nYH6je5qm
3sMHhm5kyJ/o5tclOeeAPtbmZYChCJ/eNcz4d3rhDtplJYL+QlaiWxaczScAyVfOQGBJmK+85Gjl
WsUVFOxY4DdB4wtoG/45LtS+iXjEJ1zPjC7Ye5X3TfyaHM1ClWSwjQPiZWS0cHp82rkVPfcXluYA
bfRFCtpQ/fr7Q+fUtsCh9IyAA/V32E+kf3uUUS2GOllna/yViUXp6ss6tXd3kLwJQutISpDGQyyp
noP9A9MZ1A7+zt2XAUeVg0pUzX3Eska9ue146YIwIQFLkpQNC0YRgrYUv+h5lOO+vs0TCNSnfMIh
Q9KObd0tJ4W4Ny/Tyh0wscUHXhqMqcF7iFuy79RfNIYVpAVoskx1UoeCSUm+tlMFka2MRvwtUJYn
EqlopzGTBz6hwd6tS/S7dPj/68LUOS7AnNNWQs889Mbc5FvoLKEZdynrcbBr+tAOWrECkdENK169
+ccw8T4vvdPv3s838Z1CdMhgSIeUBwVj2vMKYbl9XndW2D0ciCzGsMLpo2klnOZhpzNDu9Ejbioh
2y93IkzbJK8nQn+cdAvrowKwXLEPgvsDYlStfgi4i4rxj9f9d14/hL0yfGGRdlu+hksXb/YgWFC3
bJpUTpOsm6R3hFP91644XzQHxZelHtJiRiRk2lMgWYWkiVur1CsMDyMecDEEyEp8HQTsoarqfNT9
P/umhIOmIu0tp1xs87BRyar+84+MIeIhRSs96jGowby6nk0UY2ygYV7KgQg5N9YwRdW3i/ibKYZT
cPc2hAHaVDkucBRjWFBXFbY58utB9FH9rkvRGDuMs73TX6ECHmr9A/5Al0+pNH4VDqJKbFB8lzul
g8L7HTvr/pB70C068pU1nRf3PXC+SZfIS+NyG4hckNiE21IS1WX4YXHWPMXaRxKxALR4SN/g2vXx
JzKtsnQbNWw1SxxMyzQy1SvN+NhDxrZbKbQJsrpmf6GXNfHbTGOlbVP9TZoyi/yxM0LBsZ9jzTHV
TXKDtWSpUd1AtGe+EP1j56Y7QYEcuA6jIQh/YlQZPV2iZO+S5YwWqedmZ0SEWxbTMBQf483f4mJf
pxH2rLD3Dn1AJkNXR+Q9dgDJ5dUPa1XX7vHp4l3LFD+2bHyAJeBH3wtx1sO4p1jkRGreS0AQoFe/
T4A4J4DnV4npmAL8Mw/kMvT3670ctZkeWjpTyU1KntRUKvMtnkSH+LUKlxl+5yymqGButzA+r1DT
xkO5g6sJDloNMZCDOFA2lntpwMHzT8YpUNCD5Il4vFSri2izQtU9P1Lxk+3ykNuGxNl8ij1auywK
odoH47H9+5QS9a8d9X0OJ1eVxJIiYYnNAaV8ZC4c/GLrChzaKGNFNTAHkWhEKFRnTf0RZbKNv2JJ
4nFjzXYkRscj4VrGWKds/ATYiARTLiusyRG8sy52Sd/f9VCH7jQ6uH6AGOs5UhK+ssNSk52QI6X8
AfRAR/teGQbz+nAG/qfliaZg957vBMjMktifkxLnPaV2gCwKgRdImFxvI6sGy4gRIKOQz9ohM62j
Svk2MyozFhW5uk3eEjEaB5qTQ6MXqpm0yJfKHOIIUjzTSTnbY5fRAqSmC2xOJ8uWlaPgl74rtFGd
+dFUyWcf+ZmKzA0ObKYDZMBKgvY8zDXcbH0qoioKM6CP6TS8S6SPQRzdcE6ClYRlD4I6gJ/z37ad
KNpZ16nYjzfjQP3omLTBSV/OcogOCtxnJHjj6ZRM4suO3Ga2esiGE75WcQPPXXwts0y9D3atQLfw
ifbdUoRiwX5QJREJ/jAkfTQJLHkryPTA9QncOgLuBf+uLhpdlKWwvze7K+FDKUNxEanso9B5vlFs
JjOWser8MHCRh7rINH8wuaXTRO/Q3b80W8as004zsQvxFaSwGkqZBuOk133CGqxhkDlmFmON88Wf
xLvmrgu1RdKd6sGiX+RqzuVQXsHayg7u7bLy6/8uvrkcTeDGjcc+uqLOFMOmJC8Py6wnAq2TAMWc
aU7+nP4CyTlpWWoh3saJucSfx5l3o97sizEmEjdoXdk2P7mzsc92flkTBFLkwxZYZGbEqxZu6OGO
JisP9INC10Q1YRg8u4R2PUSK+/pSqwnNbFf632PuNy+Srv9J8bNzXayzRRaHI6TnJqmAbilBr0ht
jurVrxCyhTcQpZICBj8FqnjzSOL49U5aq+JePexGDnQOdfSqvYoddQbTSUxG0wlmDQ5VRZBXqT8M
lzxc2Pg+qlwXcv2z1Xf1VvUvS6GbViE+wM2KS1PxNdK+0dEbEZCKJg70ocCpdxRjW8dN5AXj1/cl
5nnOlWJZUfEPqnGeaBC3A+fJJkOoVVbFxgskZnu85fd0KSbkK5rm5etV4LNpTKcy8E0HZbSNGxhr
OSMvToafH48+138KEKcfHRTk8NBXLqrnQ+flwpR3PkGYwFrK3r3faikqOGOK8ye8r0l8QLkEEw1n
qTqchEmoTCH1cqHV5Bn8iOJTBdT8GQ3TXIzq6Lp9MAssGZ7m86v05tb6h4oebmXUIWHR/b20mrhD
sjoIjzhrmai1Obdx8EUju9Uhmn33bxB69mari8qTsqwXP/EyrWa5jJCiG01CAVN7oC8fVUSeXjLB
HroQRBQ0RhQt0V6nW2qrDYS7Ssk2Xjr3IF+vAbuv44BZF5QNa8wQzhG6WxaZAWZPeF3EBXvzXokj
mAvYm5WCPQ3zYMtIi7j6XGSuLjv/jKkPYz4z9tqoMSHXZ2SV3g8QsfpsDsInv1D6me5tFZCjYUE5
PR9JkfPvOydD/wK7HZBJLN8sXqIvGQqAYB4kO7WTnyFYfUA0LEhagLeq2deDjX5YvhWdDTaXF2x+
NHdfZOzGgsMoDPzTEFlzdg6nx9CQAzmh5wJPPBJ1iElOMV1VAOpYZMV/tehpBVeke/zDvD5VUPjX
QGYUnPT1SS6idekdU2yOriMHjkqlmYK2zM0ynjCumulB45BiVOrUjQF195ppur+CRjxrb9S0HuSP
OGZ0FetttXPJiJkItxyA6xmHg3VH6TPg+z4eq2e+Z+EeU1R0HBRj/34H23R84USK9+7mNsVzWXMk
3TcrPxyrLi2Hhm2aeG8V/DFP01VstcmpzwvjfDqzKe/2FP7SRsaKJ7qWn3vifu8LRutcLK/TOGJC
5O2VWQ0efl41IiTwFlEzdMncmOdfnzC627sscnF7XHJX8bCUmXwulYuv+OrBPBYIM5YMwO4haxne
sSsQERlig1xT9IXKk2HszMMGLaqQQSm7jmMiff3PcK5x1g94UiSWSJ+vahxGrXMACAMaPHFNxMMi
I1vfwL61G+WKnLeE4RSoo28ZX/8f64ohW/ALbVmLAKqnGutMfNNGfnkYSdP6uGUFJTc0OhEQh2+s
Sk/3HJtQsubeYyHaTRfifyu7q5/gpvlLlOoIy4eddBJG6X9od1o+2wrt2SAACdPsSF/UuXFtp5do
6ONGFxenbUX8KbEf9e6ID9e5nlMTb04Pd0/RuI5sHT8jarQtRep5ySxz4274L11PnonnunZ3jsNr
+DMaoFhehnUZ/D8UYMg/geMFhLKvJb8pUxFyXZKl93EEjzz8hBKClI61qRPvlGnK+dCsOBBM8bRQ
w68rzgSj/GpzhS0PY8txwbhlUK7IVoQegD3/sP3SEua85ZDT/J/JVURoAVSjocLp251o+0wX5DBe
zBwsIdQz5dgHFnGQsHIAmWUmLatFIX7cGVoh3i/FTRlj3xmqzL22qEL3o021FtwPwWq9QHCt5tKJ
b4pVTigkISeceZhmiGBQcEakPzIfDkWd7ZtP0Qn0NqQmqvhL227QkTLJcXhlxkXwDIkf9wcjyAAW
/OosC3LTV2X8ziO0khashM6T+iD4a9nc1x7gGly7tAUvT80987GJRYIStbi3F+D06Ub+YT8r6rBo
YIvG48qyxSHwvtC92WUbWRkDXAjI/XQfDq1epzxfAItFxxG7ZanXJrteI16Yw9QtcqG6ZTMb0nTY
rXLmoVwG+VNBOLHvt3HEHBcSUzWLv+jQmzG32gJVDNq5pv6zi2ddh84BTQ3t+fEgyxLUk2bnk1PN
8q491sJCmmt4OFBacIOAYyY/gzsQwA5nfUYxRVR68rJx9Vo8kIIelyIutF/bmjMkTwlLEhOAuDJk
+DlIBt0C75wYzU3ipQkPx1T3aSwhX094cSOul88/TJ/FihSaSzxKINqDspDjCWQvLG+kvw2LJmrv
VJaAolFLVnOt+EIYpCh2zhfK0KWEe9gIEVfF6QwKYnjkYXM0m7NI7pPiJMC0hYpMV/RgutzNxy2J
JoQGuGv1HpQMid/L7gSv0rhpp6fyqA50S9sEe/ytoPooSjG6bCJs8gNgvlTejMdp7nffsRHCpyHa
LOL05vQKhLmqz7a7twDmNrg6/9Bdy1FKpx7XDK9JIvBvCofNfm69TPAymcP67UCfilrCB/xEpUc5
312fYi7viJcXCM4yx2/ZCbluBBEFyctE2jxHod3QHhGZ1lOygfwFU00WyPlEZ4tLMryvoK73aczh
rm8y9WZFlOZMuHp/K7lNXpbnKnI7mEh4zL8+NniWxtkrabzQf+LPVdjrEKlqoLAM1wLpzJQt9Eq7
K+TlUG/8EBONsMUxqVzs0IjL2Ylp+co3A0NXCIp/a3pXki20vJCJPwSSEbtEdNrYeseJZKPjyd7G
S31F6bTEXeSkQfOdZpIMmUqOOG4ESdaNUaCuQ/BA/r+WYmN9foh8B3G3K8plXrckY8TkX6zO/Dh8
m79xQ98lefx5iRQ/YRncSCTlBtHii7wRU3t3lIS18I3iJ5f8LLBAPXY5slPfizhZw2t7m6VjkOcG
xe6gRsM/nTPqLBPl4hsm7CzuIQDmy07WuuLHregj9G6+++SZXQDIOYc3A1gqNUec2KdqWrHalzXt
9ty3BkmPb5c1rQZVhPff2sULegnpt+oAkon6GjT1i4MBNtGKRoP/hgkG6bJdETOHs0+rmmoBxRol
i9DPLyWXQUlxIO0ifEnf7sC0AStlLMaFb07xOwJfEnINs1JS+xWX+uebyCaBsS6kzBdkjypTkUSi
VcR+ZhA3X+wlSq3bzPFzBat3XiApHSTTsjQxK5XVn9UcUWx6OsMlFd5S0MYx94Adge0Q7gMqeq5g
azahkjvYUaPNSKY5r+egXUYNFkmiVTchNvsgOOhtfB0yTQyJ36/aFfzH/xnztRBzQ7I75Vi88IZq
ARWlh3nTjj3rtUEbORUP24UhXq5OOro7bZs4d8mXwb0HdxpIQruG29mnx6ylVShphvkkGlmuxOzg
5DTBuPj8VY0SPDjaF0Qg58qEhYkdBdrVxijBIT2tv991bMKjOlYvpEZ4DYtK21nB1rVCMOZk1ba+
MkJ26L/rJQWiMzDUr2k+ugngVJdTQkRPTzXTXfnwryo1O+3DqnvTBZVHpLNyUtN/XOQAHiav18YM
9rRMquPk+yaZUMMYiaR/oR2xmLNhrSIAVFe8L3AY4efXOqGzPo/IPmHwDJJoiLghcqdj6Il5hT0y
SgerR37OB8swzHSiBZ6+6SKFZqXPIs/MlbBMAfzi70EQFXpw2hTsm04qFtCdzPNLNeizRh/vRCJV
8uO+W6Ah0F93XG3hIHUMiqaRYzKbzrtglzeNLWHHjvjtHV/Zy45nbcUxI63mhEiW//02lcJRDY/8
cAV5UkpmiO5ld3RqlsgESgBt1z1fXF8IuRgpTbyh/3+hNuMPx6X5F+hBCyobqC1lK0+4M07dxvZX
JITegUdXZqbXNi6KjVp3KKEjgR6Yh4LJ0p09kufRtUj3xZsjc4sO2pto572Vn7LJjt95/RPsvG6o
0AEvuGu8/w2Az8Y3S4vzZIlVDQ1a+2QR6u2MwTQEtoF9YL+tflCjt6GrBl0SRl2nNuWVXND+q6u9
z5qPb2P3n1Zaq7/1ZExSLn5dW4tH44u+PslP8nRNcSh5mKX8a67S+FDo8TUV7wDCvHnIbcl+6EwX
QRenqPXgQtzzphp82WYVbl3pItZrnZOEfcq9jZZHhWE9QApemQjykKUi5wmHaDvC7hTsHsZMgkX9
wdf3by8w0IEDu/vuJbDAIEqWp4nm9OffifDflnr9/+VK+NTR4RYBlPgaaQmPgClxrfuwrtf8Oj5M
SM0Ccmi9KAx0ZWMxz7bdDJGRqskwgk/Qjza4bq8hNR9FkjzgadbYvaBQzg74rIjq/sflcFCvvhcf
KXrVQ0qsaB7LriB4xV+xmi56NjWZifk1q4iPknEY9IKh2ZLUPPaUUUE9MxUXg805FL45tn8eWUNw
NzoB2u0odQiYxsE5U0b0XhfG++53kTO4uVLPtGJNlj/28c6u4MFnqUgtDKmw4iutgjdHtPZpqhqb
VCGf/c7n/d1x3McXEa4aT5pSDMTyujieW+PQtdCV92aj+OOsIUM2Hzs1F6/07b5w6IhsZsqlQSLI
AsdKPVGCsGrxWOrR8zui8qgQ33jovm5QaRxfl69AWm8ckG9BGUq4sXtNvMEt7qHOOOn89aTfrJfa
jvMzLWjNdZ9wsIvlrTKOq+Q5p7r1PrqUYFoZyHVdyJn7HM6wz+lqHhFSqmUVY7RiakvGEFoCNWSM
e0F024H/CUmzsPj8uo9fCslRRL+85pmGrW+10mZEvfXMeJl+I+R68pkHdW8jv+hPNyDI10UDx9rg
wcCAC9SUfhkzI8+xOFLnV7HLgh/aUEvEdQt55dCUV01JJJm4Bv01E2bjZmwtJsWtwXCjVN+duIk2
7upCWkE4d2oNu+6ZlA8ZqsF+ELaVPam15UDq3V8ZLuOky9MrVmaCvqmegQ35TPfgXLnZsUbWuNZ/
Jige3foE2bOucFHB6sBL6BZ6zXbIvhFg2E9tkzHYp+62eKHMHO6THZxXKICGPLoVw+n2I/nycmVK
0J0tedsem5034g/3BrjW7WWrAYaBsKsji6etSlKNPkBQ2jPOAjNh5KkX1xZs5Mcv9RrCgj6TA1C7
5VlrIJgaGJQdzXicP5yraXgpDnj/tLnOZhd6iNMQjJoUwsEbzx6Kkw92bjpp6wpULJna4viCvGJX
SMa5emkZ+ug5zVlLHEahZJRFLGe9RiGqW1RY0oK+/zTdd7CwBpOS/zmER8qykekZA107Jesez2Ki
w5ePqdiwUn8DFz7rXQMAkJKGCfxU5WITIOuZpY3XUz9A8DVBjNJ4hMYqd5PK0AKDrKhAJU3+H6HB
qqPu1cz5mdrYPWBWvRFubD7qJUxrMUm9Tx3Fbs6tQfboUhZvGwN3r9IF9G67FcjwFeYdFelQUEZG
P+lPuaMhNEUbHufroUJeYPK1KuL0ePLkNZefp+SVp9vQ8nUPuW5Q+jSG3RlrgvsdToSCtNH70wgU
JPWbtcB4MamYbc6hhpdbxX9B4kGprhv3630dcjACbnC72FRioGWZw7qs0YP4fGRgfHf1nR5iBF/E
pX70jGwGz3espIXIY4eeb5OT6nvtOSI8/JrP9CDHP7py9mtlADWj1ugZK46f7/uMtIL9YkVzVBwk
9rDSFOyPHMetvGSQIJ0jpeOEcpcVwkJaCNRZht6XqEMHIFAebqIJJYY1RKTvDG7Jh3cCFn6UOyI1
bsWDf8WN9MWRMjocuEhq2TOzIu7IF/ZPfJr+qosshIi1yzKeN54JY2/jHU/091lt0vUgArR0K4ka
yMgtYeH+NG+6jtAEVy08eZB3YACufzYe8qrNfBBa7OrfBkuckGpEuuAft9FO1WD7H+AaekCuj838
bnNRiHyGsMEl6OeF0mgCqkIQHO3P4tqoKy7jMLEkHFB3c603cFJ3PXValWeJZeucyZMxYWPcUcg0
VckSY9qTnJHMuRJ1OBOkmIoTPc8PlaXdZASsVovfJJ/j1cVrOJedqbVl0nZFPzv4gsMGOGhkFmNR
wx1t+8SGwdKD3Kg+KU97tHjSpKOxlGthuAHhkF5qc06GaNhQAbdMSEp1vB7wdJTlgSXs/Wh5tOJe
G8Oh9iHenH52Kjuv3DX+YDRhtaePnXStpQrkYCbv7Q10Jol/mdEqOoAS93SgjVQbJrR3MsyH7bHd
yvXqApzU8q0V9La3T/2REiVEU6bmpGNv8wLypfImi1P7LEYIrZF/hW1BAs+gv19s9bNR7iB7mjgA
N2pZM3PmYA4jX8vWr4wjw7ydCAq/zO24ZycNAPzG394LcfnprRDhH+e8J03DcpkPXkbS9uuGbcr8
AlS6UrHn31tr6RlHo1FkAdi43M59VAKvCC+NnvXbjmIxS5GkZYzVN4tNXnf9spYueFj7ZLHAqV+C
OyMdaQyVWhDZi+Vj5uBNjjbts2MasBtuM9NNoVZRoGJvP7VP4WziapeAB8YZWGKoZL95VEChH3+e
QOYErmsV3uSVMfsKDkM8vCyWWrsG+Hqdudknrl2SuAgHIcoKyF7q/YFk0OBLbP4/O1cmd0R4DEj6
tJbpXNf5ZgGZniWd/ulkDOInoUUxyQz+94ic/3byzOegiH43UBmg7zrkcUrX9bGFEt/gtyM1mdYu
FHnEiDCheOUZqg1NGaqzS4iB6biC07NlWgBYd1waNiU+LKUrp1Fij4Quz42A7jFXKtG6czZP6B1z
F10S9U4v2Kxmy334o2loYyPK22UJAFcjJQaZBDNU2SlrY2h+IEN+t2f1p9fd2xTxYxVi8gLT8u5F
DJv79lIwuYm0cDsyakbkAXtBRxcwdOdb9JeUDW23kVeAE2Mk6VwWxJW9nlL7XN8A/3ZkHwohrfwN
nx0k/xkmqk5hNb86OKbvYJZDI0Kuq7pHP+w7A/olAcTUDJROEF8dnQkgYHHJ64Fk5E+j0YTboZAl
0lzjif2OPhncnsDajuJcMs+DYw8wwot1zdYYRsy4DcBBoqLWaEPdVqJmYCNQsbwPGPwQ3ZuDLFOx
zHMpCjro9VVkfpMX38+L4wmUsJaLCygxQgr19+lm11qDQ8yvJBbqTbvqZYt/VNe3UDT4FNRlKgYz
cNgToCMvCmALTz6qzu3RgRifvvMvXKESao+rMhXUKeIdhS6FfGvUzTmB6N7czvueMRFGvikCJPcl
NIlNEzPzTGHh5UYVs9ddTidvxIk2qw9jtlSsDeIIvJ20IlRenlCI02sprsWdW3XZf2SUITWvxw9H
B3/cNJFNDgvL6u/Uw3/Bmm0s7+vym8wu0tTld39QL0n3DLGkX1fmnYxxVdjN+vuoaZAzA3GwMGVI
x3TnLf5q63cfxPu8FtN5D/KCsmpA6N5NZXlOyIvNghaJbTyYDUjdtst/2TaHFSKlVVAdNEZA5C/V
f8H2kY8BT/2ldmNMw77sYpEdKIo9qLKWhLA9TxHuBs40dh1ww9IELHsHM+JVpx73ZMOeDooPz5I3
2Em536pmjl9zafx0fvJ40GvChGpzj8zt4ymiNp90WmdTIciAsRcBqunrhSfCRQFPORmGpX4vbqds
1wrtsANeMgFjHh2K3yOu6wGjqPw9+A4zOlOdqY8M94VdeNljNtxNecO6Y5NeLcnD5W5wtK6S+ocj
l13upYcgrD+0X9OfkWGBuOlq5ScvCOhdrRPSi2wxQ1hhLBuuLh4epQTGxfG2VmgtWBxJ+sYNAtxl
LG8OJlJCMgSHTiun/Dxg8H4Z4/8JmTa+BFqsWuGXf5xAEBSLqTN5gWZKNkzLtmAy6yX91jGk2Dx/
1P5sWV4kq/DLommP0XAyouWI2/E3JxsJKlWJmhK4gym2E1A40FGZmvHsdN45+zOlajLP4rJoZpjU
zer4fLV/t6MHqzFzIUkzNN81BmOrdtmotIJeer43tV+7sVFrJ7Bua4ufmEnSw1DUSHDLy4bdtzJw
CAzEWtKxoRsoOOEFd4C7PLX8Pfzuj+7uw3ZArYBAEexDjhtllNgXvq3JnymnUFyBOYFbJilTUqV6
QtuoEwZjmU48IHrI+LYGkIeDKYYC4WwMBkI4R2NOpJMDfwcVO8sN7dhstnBdTSz/VMLO9ZGqtsPA
4LvifC16qUYxXwVXugYIFDR/FXz+KFMl45SZac3yDYWC6nGTlv8DhBacdO4bsJdeYjjxLaZkLq6i
dbJZu6QTdjeOxGLN4ZJE8DJtoNN7prBARvYiFBhwHsLCOrJwkQ1jtJ0tn7AYPDeyfbp6w5+mAlrz
BQ+6mXcELBLdglh0f+Tv/201ZoRuNBz5dECrxb+iV2efGNZQhsLMrPtSbgaD3+KQNf5p7wQ5AM22
L5jXxoIb5uhrG7fqLaKT+8kUEjVKph1BOAYfizNPWH+86u1SrPLftTDPwUvcTdByCbIaDHCXLHu2
HUcCEH4Xj9XFtb35wr4NHtUaDjtsRwiR4kqgTF+Dnxit2PTjwOeXVhk8UYLETgybb/JTaIo2TBX+
bYjeGnAwryZagMcX74B1IV1anJPFdqzfpkOt7uULKmkMEhU0Otx1X5aS7p+l36Cq/PhViwXRrT0y
1EpYvhTiViAxYiSagUDQfyGALXajTb4Hna3emjvaP7obunhEOWXLIn1sWIN49n1Yj7Ib1dUjBNKB
l3yds0haePakB2epVt3BnJ8soHNCzx563xxUD7yG6f4xoq+kNPs8FH3Y64OtHioOPv7AlaSfqCeb
tZamvdP/W1ZjUUu7e7csKvbEuIuyftxuVT1b7i/M/gP21Vvw+MsKy8o5Kum26uHjyxLZH9Hudomt
vnSygMT9zreayd3+/zdNBUBRRrJZPNJ1tLedoSzm8jXZyCAzCq6VrvYmmRxWdaUUQNzWhv2yajpL
XU0RpgwxF+6e9Ylixy4Mq3RF7Bt2g2fMTTYVFiuxgAzHLMHKYgIi4YD5rYcDQJy91zSE1e4H7Dqs
hQZbkvqonJulTXxGfUchOcPHh33fSkkdjiFhjpwd4gp34ae1GkeIZ+XVH1EJMtqewUYMLN50dfjI
+cCBGBxlhaG2j/yCjRL7Dgnd1iTYDhy5CVhpNsF0kPzpVT84u4/zaz2N5K7htk/XHd2k/yFq8dX1
rj3+Sc+sg8lkt75vFgLRWgSY+2++QXLfQR7EAn2He6/dvuhYWlcGwlyy9FHbVeZha4s2X8BjWnVG
bImXNlOVSQnYB8kWnuv8ocqdnqD+H7tp8hNWE1cMQZDhNNU5fcOfR1X+ew+3PtW465B7OBXAI9/3
9IsXZMdXVKVcwbNcI4Wl1R+cdfncPp+AtNHyWULPJt+EHNIFmdRl9X55cWh21K4Dssc6WrOs+7Pb
NRP2AmFfpMTkZ/a/rBaiHLkGKyIBImPZTTPoxeP0758pT0fBjYixRDylxUhxL3Qiw8sp8638A1dX
N8dlZm5D2G+ulPR/wGZ87COMgx08Icp5D/6dbdGJFmgMKaq31/tyG5xgLJAND1ASFPcNfGCaxmqU
Pj6MQvu5Nuh4I0gFEhs3H2MvBXBPuDj9EvRCR86Wn/6VXi+37h12Z/jqkauH3Y8jfN4UOE2u/bzo
wJ+OQDe/jAtLmawbOBZtbbtqfbtG2sCI66kv8A0jSzzpPLEZAgXo3FPRDruLk3qYJb4fn/CeVVe9
VE6NLnVk72qTC/pnTus3xtCjl8NwO+AkXVj6YNlwzv1weVvTjz8LYmMVUad3GJMLgdEX6loZdAUS
AKxddbP6CkwBYg5Rxsd0AP01GKhwudL2RQZaWIVvFqL1Qpi0jsJy9Y3GyEQneVj1yoAFPjmm5Wxw
p8gx60f1lB52VtXivvm1b6X5a3fz7LrTi/yw6KItiJqUry7g5hz0V12t8UGQwka93MC0Q82XPiGa
rSwhpili/hNR1Vp1suB0bi5B8u0EwESijCzKCC8ekUO+nXnr4x3Zjqjq3LhIHZ4SzF48be5IaF2g
xs8JwdLFXZL/g++A2VNe6VMQKJGvwiA3EFebxME8tFS9POxhNV5C4+HNnjuLvL4bGhHOTuMk1dxZ
I0MzV6d7kOm9JzgExZqn9IrCKlxD8Mxfo1DvbBPZG0INNKKRx5+FxrP7NAIpkw6pNwWbEyuX0rU2
gE2KEhWacGkNJnb40FKHqzh/RVVjd7j8WcneluZzxKCSGB3/lZwzENGiS81r35vyk6kCWVrN1PvG
xNzdm5h+scKiqjDOwcAcjAn1y3rfRaqx6JGDuzH//JKECkUXEGSyT3rhEocOi5wLahSf0ubSSmMK
u1+lYlrzE/BfpKo6R62GYKbWsgOq9HUwQ/d8dmRpKzjCbXI7hg8z66Z5lUSd6AGcwdPIQIL3ti4H
nnzqfv5F3kzd+9sZIsjB6hsYBfbiCgnUy270ZW/2v0/F8i6ORDpe8UCvy8hmo8E0Rj7B6HCjJjor
nEWNI2YyS8xELsikr5s8mio0FmNjWzoIVrq7rhvEUkbPfQOQUehSgY8kuTl+hXpVcp3iTI9j1ZUD
3QDjw29iFs6mp9s6epdtsa3cCR6iqjwXNo75N8xheBLxDdDwBVV32jH/YJwNgK129/L1oLyC9h/b
L3+FRav9+CPA9rkluBShsl3x9ctcRsnz7a5aM2oAnqDj65GfGOtQDIFh28iojgphzvtoduaqxkYM
324zJbjHiZouRZ06QdD0+CMfLJ2YnTkoK+JuHLWI3pJMCRG7ROapAupe6C+GGEHmoeJaoKlRcF+c
1svJ2G3TEkEd9TUNgrDeLJJ+YCKECCnUnt34kRjzwXGBq1erIekQm+qdQe5+9/tVwJbpvPUw3Cuv
cB4dypr6b9XYjFef4Pu1/7S3EAXKNETR82TIrdE5jYxl8RqpqusDvDNH7DkLgjOnCLWJCZ+7b478
uj28Spr0Z1rvyXhYcREHlJbr2ATY8uIUwfDiZdnLYvpyqUMcdI5WRkkPWHpazEZCj3Y3/jbKyE8D
FQb4gSqsQEq9dJu0eDiHhRB7Ly83m6lmKpg4w31zcLtw5N/419zlPH3EUeoYTa1nHALiLI+/mv2q
SON1HobWREf7/fOybGnM6IxUymQvYyw+X2WdP6741cqLJquMRo3JXAbQV1T8CwfF19/EbeE4tNIW
TLdP7ZSaptqCuzsmt4PP7z+AkgzqxlcIjMHB2mbj9YmSoMpN4CSI5yXruzJOZN/lDBtfW54unPIk
3PgdUUm3Vu0INy7tgFVAn3wyfVFSkxqJuMsodfDS67tbF19YK+K7rjCt8cRm9qAAgnqIwFoH6d0+
1gWse5fUv6xNBsXI1Ia7bpucElMb4C+GrP6OHyhRFurFagUNcg2UOmAchnksvp4eMagnsEV6EbJ/
3aUBPYvI32YOc3+njQstnyXiAmLXPVkhE1+zMtjnxgTcjeqtkoaFO5CEgcAQHeOHPZDQVbdqEhsx
iMscCi0LXfGGmelJzqmtu1VEq1QItN8gUBx+SunKSY9sMEmWhAdrhig1gcwn75xamwuPQLkQFXBU
0+CY05sNvvpWcMlhfSUiV5XXW7Ujy2wWZKq0DDSkfVVXco66UdgANE8bxMRPVfsK27hcBc6b9NTK
ULuDgFme6leqGqu0D1sKreig+5sLt8kdl1FDIDt9o1egNaJXUu9Ghg8Ezoh6df4JL+yhu3nb5z0i
p+gxEw+a1V/fGnao1lHqKNEdjq6acYQOzBDfvu8Nd2DcVKYdg6d6/r/Hv1xJbS6bMYWM5B8PEBTr
3bj6FHXZ0cxdpp/KrvaFbd+Oc5xrH7U4WwGrXSEF9nND3pCba8p82PEJlDja0cCFrZMNAaQ/YtJJ
edSR9pp3/UTViCE798+j9Hth6NDuUPR1NHXnz2Su5YoCMDy4RD7yGJnLEamvJI9zkFwDiy2ZrZ/r
xDzJ8eFKhxeoQt26M0IeAKGatKJ1jl/g+bv/bY34oNd14eeZDErUNXwmoUrOtw7uaHb2Flx5SHW0
MfO4aq8rVhB3vXq8qVbSkNwmxSbgdhFIyFCYAKvyu2CKyyi+N1ssHDmsCHBFfrIYnZE6WWYC5Vdv
fDctn0nANhiA1fjylJ8zn/J+zsIeEFP2115gWdkEUoyCkQXX7RE9huC2xi7WlH8tYq6zOUisF0mc
7hMnC4qA+qvRl5LXvKJQ1V2gig9KMULkx0D9d2rY6E4+a04jZIvACRcJRRZpo6kAOnK8o05/yVuK
w8QWT5uB/9A96RDHxqa8/Li2KSxbdY+bYYuBd/yaHtf7/nI/X57L6WPFY+zCYbEAlhxcu8yyo08i
0S/qBzrQKEhRbjEFkvcIfAwob2Z4MThHpnwAVTF2ne+7aHB2mGQXkXTu9AoNKrsnjl5TFGa1+qjQ
8tuAbIKC9qUKSTV0HyycEGYfl7h4LZ5wwyxCJ1q23jD1qdmadppOr8cTr1HRwtyqDXjJCnc9pw6Q
CmEeY72umsUU64Lz8ekGmsBmvwUpIDOohBAEXC29GOpM4QlUT5pa+MGs4g/zEPSGKitzV7dtoCuO
4jKFX3U9bpSDCxUUaEsuBIrKUT/sLh58rSI1s/XOyJOYJ5nvqJw+bLGPmVAMtWZcdblmYNFzNS6s
41gyse8ApMsZV9g7EiNt49uksa+1qA/Bk7/yZVA4Jgq/wVLUHigLGj1aa8aalyU1xC0rh3UhCwLb
s2fS6xqSFQTJVn283GQXXeP/iMwwArmzHBmk6nSIGHPgl7zDrala4bw8BKEC0SpVAY+xFWyJuSBK
mvhujtHZNWbMEEYcnPC82cbRTjSkSWgR2xCY2wT9PfVaAVW0ukImHDspzQds3wSjU+Gv69LesBH8
zIpMdQRdN0gXjtIjmFNX27Wkm7cf3islKDSM+NQuM6wBFPITs6RGh37y0NR16sm3IwUjG8JYt5xM
6ZELnpfOYTow5CDdyIYc4o4RbaX8owKp7L6CYPn5dA3mUYG3jXOV9G4LeyUuZwdF9YKnj7mSxAkL
YgCBwEIC7rXXwZEAlMv7TeqidOOoQDt1xhXmONyX4M8mEr2SKAff/OtAgpRc4FBUrzuAC1m824As
YtL4J1qUJOdEbj/8G/UPCbnODrem7itlgcPvY4kKIbttxvrAvcHm9lFI/4nc9uujvtOq02Y0Tin1
6hFqykgi4shouQVf4UIc+WzNAdJIWZDZA5AOFKJFW7V/5ZLAIKKl4bVyvs6NOIvrHtwiwArVJcIr
hGX2o9+7NlZsUE/BD2ujMEk9h9qPFxu6+kvBH/bvWuBpEs1IEJEnPhdEDQDCZx1/nd+9KrT4lqgW
aEO7gmFqLcLBUH5XLALhxdaI5q+1VCuzNzD60HBJ8n/tineYaGkz2zxBQFlmHxcctFfItMf5CnR6
JOulzpKdtgvEfKyUg7u2ycYgWfIliUG1jICCdPrpy+wkAC9U/PIAt2Jpc8Ny8Vt+Lc5kD0yyrNs2
FwP4+WDaZkYx9SyuDqyABX3UtCsvHy8bgBch+pnMI5pXfgU0TWKfN7gNfJxuFjfNV7spgbkGUcqn
LjM6d5AiCLauV0hx+oZ2KQBO3372PWxZxAWVmNgn8fVbdD2gWIzY2uuykPUNoqJsau4L3ndLZr4+
ylhJuR81wnCLLtmJjM0uTtmbtu/SRL6k1+bZ4V8QbYjx+7YjwSGRmpJWaW5M2aCH46XGrkwhhlbt
Dh22vdehnGpe8O9OATNoMik5zo2LdJ98FYKkWSDAagJFaSCg8/DfPTGYT2QD/PtJs0rL3y/Obq8c
SeUWif/N9nnMiE07C7X0EeOZdY3Vtq69rAUdW6jTSVQEIoLk2bZsp7gUkxsRYLuVMJ/EX4iIuHA3
jJe0fbzCLnT07iA00qb0DRVCFb00rfcyjgunBZp2YqtGUrvGZ1y+fmWIsVDMHPiXYL0Rf+W4hARR
+Xt+rAee9kB9WAK6u1OvsuCnUrqnNGahHd3Ae8GOfsbJI7Jhow4kox4ZRsOLZTkb8M5JbiIFPEpJ
MOIZ3VvLY3zCVfXVvN0UGjKi42zMLXVfLxgDPZcuki/Xh7tEBlgFQoVUYGFb06fDFI53tih3eltW
o7V6j2HLCPNQoJkT/YhuRAq9XFTlgNoKdkbIUsKh94on8cEXlOAUgdjWrFD1l+at/DPf37mPGU7B
lzAYUAz2wvughjRp+59iib1AYbB5NESRScendvZ2tnWzv3m/RGmsG69xHxyVv8coruiYrN7bGdTn
i1gUEig3/2yuHbYW1uslnK+15wWvSXYi+o9rUsZCOATsT9AP637AVq6NBQfzoWpqBPuhbCCFqP3U
3/JTaFp1etQbscLW2VJc+fsOkXpb1hpJNWDeOiJCfUODtBI7PB1mh6xTqNOsoOd2PERkg+fwTpwn
A27J6XP+cB/Vd+ROV1fRQ/c3kSeAjjIaCKa+T5NeObx6ude8JMINl2GU24jYPE54FV2yAg0BEuzT
9d9BcVRhKJKCBjLo4lh8Qo4es+ZulFdKdiJWS9fBSHlSNNiS+s0A4We5weyH2GD3p6Ux23yGzJ5Y
XjJCQ7DOZnAKE+Ff8zG7kjXjkI1QthNWZDJJ4qHe4F0uHrY+96dANDxd5m1zZ2KU76At5yeVHP7n
XrFm4khbzVwkQ+86l6BCKwMi04JrYZIeKjz1PhDFYBGYK2rLQfPR4KE01JOIqLTyQWzUEgFtdeKP
yDNQiK6IxiK6QbNC2DvkUwrxQPxGM16Vr7EUT2FLfV51wNIwHIjLpnGaqgfuUAnPZP2yUqm7iQHM
ZXkWToHhgbSy8J9KNdD/UNBP6YgPxR0vp0eKzwmtOtdJyU9LfjSLsEDAR4E+yEZQemLyOH3AtD5n
Va7igt2sm8ilFNrwQ7p3xwGymLPX//5O7fzMivLavNG2Pbv9mVxLOeLJlTgiUI2/NsXaqyBcH4Rl
rdiGbjH9ZGm8TG6U0DRQJT/8ub4ynjFR3FsSf/BQ3TFgZ6f9inVbZ1sgexHChpLBCW3HtBNV2Ees
eWRjQN8natgkU/lwNwdzK9U32d0xpTAG1G0lNZ7bgEWh8gK6otHI+TKZy/kMKCHa9N838SC9l8yR
3I5g9KuqxAwoaHElW28VAynKBCEXAi5ti8wX7B8sK4IYcHmOrPoROpdRtnvVFk+CXm0Al6XBl/YM
+ZqPKQseozWiWh5VZhGcn42dDGqd4TOUgf05eRZdbGpLG1QFi5Ef3NMScu18lbnLd+w+lEPwJuTl
AN3hpTbi2Y3VscoueZfOfrWHxu9EzgzxF3jNM2Rgh4Vc0Hkn7hV2lmlZTt+m1624MHJsyo8mP02E
xedgOaY/IjAPgsZqBTMD156z/eAbfK+bX8P5mYB2OkM0nNel5WTtogjl5T0cRU/Rv+J+/R+y2tQR
KNQz/ht7Xwj21Rl82+yQOaZVXSr1DBCqTZl4syytKIqTFjZOaUjVlVwejycUiOrh5hqT78vacM64
AMUVjqPgBnYKZFVsb2hR3d4pmvLBn3UVcSiOj8V/oR/b2g5tg5x8qXHzd2wBpDMXDudyOLF5n5ne
z9auOQggXU/dikQwyn+V4uTn3rnAYjbyx5mYqw5tyrjEtMHGyfXZ0NQbj8BW/9VlzKV8ibACe0/q
dbWuML5RtjOwa2TchbOUPY+Vp6+CSBmljZ+AEYLOo/xTxsboC8vI5Ooo502/7HZt4gHOq3X0MiaM
xGUUu9qp+YFF5TCUQukWUbFbTCvtO7u/P37wJ5rTHq4lZer2HrNEs/6ZjRptxtxPDzL4rDSUjQ/O
KuSMQ6bjSjQnGc6zr4gae2J/Tdap47ZMRlkxNJWMcc4uM23y/QqOepidNIld7lXLRIl1wyJMj0Es
sSOWU/O9vuZlOkuSWC/4fuJxAkYDJxJSG+L9B0tJjRzYjTcaInfZh8ENOXDJLyDaR4ms+ku4HeEQ
VrDr/8FEO0N4iEf1j/foLtjbd84zsalJJFdbM7dDWNlFid5hJaQLUVBXmL6B+4E6WVcAaT+v8RuQ
XAtaz4gzfarRYXlT6bzLIO+Xw/jbtb18EENnrJNwsHNN3rLm1kiEMO+f75E0c90nxyNr9oxuzMz+
6QtyPf2beMmk4NhDP6+/UEUb6M6mlnXJXZs4GNH7jeupWk/wmp74UaNjgifH3wPQlRU+JBFP4T8D
d5wcBd3uBLUO8siZaEREIranGPtXBSCI3i7orhrYwbEdh+25KJITIYtS9ZxmGf14qFaHT7lb2bnA
7IBC+arRk3iBWcx0Sa83msyDAFPsknyGh0z3JQDDG6A6AKLPllXiOfz6ZvaVDO3V8v5ydjoB040t
xmT3JWav/0E3T/PayTWIvTAfID9cP4oTqtu0ydgKxtQYKAaCcCfKtJqGXzDWlmQ5lEED/+hO6ssB
pxR61PAL7Y9DpA/5sO8ww8R+9ZVGasVZzUVatwQT8TxwOel1AE75b5Ky1BzYJgHVKkFESBiPK38y
Mjg5NOWWtR/xwUWxESMbQVGkf7Tz2L2O6gfjSbf7GGUXRetzFKRdQxgezqjsXduuF6XSZNarqZqa
6OZBvSvJJhOk5xleOa5g22l4AAAUmRoUqPcsy+10kkWff2Rxc0GIypKVS0yZUvmqgh9sq+tBboQ5
SK+0HdZZUhWPYiJzLV1s3O8Vet8D/CWeN1HA1VXDc6MOSK7DXjomCMeBqGb0Y6/h9RFMMPd82Ya7
btjzhL+aZRpPeVgpDvdE7GI63T8vx90AARszvmavwYGH0tD6cpnnYhGvP6OxMj8NNAsu8IpmmhfM
NbaRaH/b4WspYghLAVrdlziBGxU9/2nQDSKasDeLQM/ViMG3Ee3AsIz6wRTj9FKHJ/yPxb3ALizL
nL3g+BvcOi/CWq1JK943DX2JtIV+YjFnx9Tiz+Pz2CIu0uGE+l+pja4AiBiRjVtpd47AW67J7jeh
eiYXiQ1bqKLw5sIuUP1a+x5hdQ9ONiVDpJVdlrjOndSHOnUVHgiuOofvASfUmXLhQQdUJvn0avvV
uhKhHQ9mN2wMa8igAHfEYPFG3R2nm1jVRqu7303F3BDmgA0kn77f7FZXk+7cBDrOzR8AQ/ScO7Y1
dzaTRjvuxN1CANtOPSey5xkoNPW5uhsBSN73WqRVYZlF2njPpXy67nU50GfnCZaTDfu49169Q686
h3kjw/9+S3UhRHcWVgsJYqjkn7ckaiaxS+nLQ5aUIWsTTAMFQE9XizSHISya/Gc5Dgvoy2+3B90T
XTHpx09r0djVAVVVHKBZV8nmkDNWjrxEx3/awuCkvn718E2k+VDIFT2pm/Eoc5QcPIX3He55BAXe
YjO9Vwin5PU7rVPiH0sYqmt06zHCIu5PZBi8eLkPeP8VMOu0E+Ge36nsNS+VphDK2I4kZwGQ2Pco
jlx+SeVs3k52ZZZGrvc5KTiV1Ls+bAEylSHOI0sxKGVnv8f36mktbvQYIcyzDbj9BktRANKaulEl
gBi2SWdyo8/tnHy+qo0zqBJv6yClVRfl1nlQGn1bULGXSiWvG0Ta2LSa274l7lXYfKntkmGhgRMR
IYTdosNLt8plNtxEZ7nwCrXi/EWmopPZ4PvYJe5GHXczMfEZzqzlnJqBRUrTEHz511yXYpNszdlH
q8rRYRUvRLuKk6I7gTXIUcKVAyXcsF27fZbX0BGLZYGaumEYvL6g9ENTLcNIPxsnQ5V3vGKEv/30
IDcbOrJe5ODMQQ7xSy6DpLfUlbODc222a1njD2GQ/Km4WES9P4++oHfK5NoSLbTM+z2y1Sf7QSwK
FrwQSFe8D2o9t0DOifi2YzWIbQF1HbC8Jj52LGh7mANMW97hZ+fg9e+DZa6VIgArQMl3HYfz9LX3
BOq83ZES/rymPYYxx4lAslnYiAt5USv0J7uqr5KZHZMpN6OWZ98Mc01lQJbfvi6YdTQJ/H+oiZlP
ZrSkXPZnyRRTvap5Xk4wRpVDSn3iCHNxmId1HgoNlx2uadCLaG3CdIphevTgicxrjPCac27+E+NU
9myUnB8PyWQVsU5brzjmK6Uf6/B8PFtElVLIn4cjwUMOO67CUI9CaGBCuLvFTZUkfDDw/jNfACYF
cg0XLvY/evx46XDNxKnsQXGzu+8afy8AzPMCJ4F/3bKNd3jDMWSeUaYS2WUEKfFjEoKBR8EdiI7h
81Wtj2DiqSDKcEXzKDFHO9wuibYGmr5zCU026A3M7xk1mraj5DAhe9JdCVRfTIKOViU1TnYNUz4z
oidPdhEBnugJqri1L8kHxlKAiktcYdOubI1TW+0cMvpKN6KOJ0Ad+gBJGy+iCYNMfgSBDgMy12zQ
nZcaNrjd6D7RP3JTKj3E8km7l5HlvFTwbhfP9ahY+KuMdW2Qr6oZLzzK/NEhQv9tOi/+KxHQa6vv
oMMUDYcNnwqrVWVqRwjBi8LTaYpRJ45OR6H2lWGvZhxg92EunU3XrheBI6lbHCRff4Xq/5uoKe1Q
JEt5iPwfM2UE2x7j7XQO53jAuDVMTy98b8HT9TipVSOFHacuWxTq/9aXshYpSdWByABqTXgdEC5w
TMUbXDWLUqSJLsTbwzJqSDE6vHkjxWZr2nKsYx8m1tLrKrYBrjMu2VfANJM3NWc0AjoeZevSnp93
J2c1cMe6HgmwhyCQPUg3XqcQQ0kOyD3jxgg5EFqp/MgBjOI7Bk4yrsdsm9lUrh31V2pEWNM/7M2g
3uUvqFPOF21xZ2oIeuKcaTvxT9/RirqCzn24YDqeOlwTQoO4f3ePdT+rCclfihZ6+bkaM92y+KG0
K5LCNKstXiVGrCOFH3Yf+F97g6Tu/3aPt0UAxg7C3eyQqbfjFZBbYZ4gJVmHGySONE/EkuXIFLVc
zz1sDCqYR9MEgBpWyB+qc6DzxArijiJ4ehdiS4vZZhPhAnfvTT2Npth2OxYgHYSlWwwCbHicsyiW
afWvwZvjNO+L6DKUiOwAiQDTB9Z0TVnbKdFNBd2QHbovY+me/8CQp5vcUwy6q2lgruUjJ3uXFLG2
QvZhIhvcPGY6b0z7BxUFYyLP8yhZ/eCgsE66LFvgfVS83PypkGxM4px14dpSLg7fstih/zLXwQmp
iFOYilF7w/+muDksD0L4mkxd+7UmHMs5P0coK+IM18nTbKn/w60gOGCIxQ19G1N1MplVW2uwZVOY
8X5gwrXiqUMZDaRXHctM3gvPsdKHPQvTojsMaeDchbVecnDDdjIVke/sN8F+06MqnXq+wf54taZ7
obBweRkNnVRug4fBm04rb3+ndLl1RvJDNQ/iA6jIM1sp5tj6jaaa6MwHTXzWYi3qPNffmdeZEm+p
jx+1RXg4/ZZ0lWasJ6wCsKBiHP5Tz8dU6AGJeZxMl4EfSD2JE2U77CF/j1pO7CoOil3aSsXs2n4G
+lByqeFDsqHZsyRG1jv6/b5wBp7dQkCc1mwCPsHmOCAWHXOb+xPxmyII/IjTjpBvirsDqh/M6pmT
LY/uPEcr3+nXBzHvIiWZ7oD3yq5wh/nqQ5QOGIpObKCByWsXdk8qb/0OhjT44ut+zEgbR2+Er7bs
nJ1B2PenEBO3yg5lxMKLp5wzz+GMjARXYVPdXzL3XWjzuWE0gN2DRvlcOtK/6POUW6u7/UkMHoNy
E0/NyQu8GaANpS2M8W70BUE1gRLT4ToXhNNQSwzpVnG9aR2klwW63xaH4twRVXs85E8JNfPpDFoS
Snv+/tqPW02WhAlbW3lX+CgSYQjgryezKAwlKtlSdcwcDHxIPbeq0W5MuGDPPAtefA4ah/i61bQZ
zMNC1tGrwiGCRryt1W/00DO8aYbCDpIybyfqFLV2IMWrLYsKbdKhMm4q/EzZss7fsD4kZ1F+kpu/
CIeMHeH37NQxIycqhu+lQ0d+61TFo6ey41MD1o+msIcTTXBcUC3pa8v+a+j59QJrDVjaynSr6eTF
aH/G9PoMx4lT9+eyc9agVxhAAZMfkabmoa1Asd1bYcefyyrCoFy1y/y5H8y6Bsk1oA8phc2n+h/a
kcsTRumccjoDzj9KGZsKjW/2tAjcRTb+Z+V12RhPpITaPxLvpK5PZYpnn2/j6aYzjWRAxdZ7zUgg
fEIHpja8rVTEUNVD/LynIq8gmstCCNRfvVyoXdx3X9luZOET4ah3ZQdev+aNslPZcikNhp4zQZa1
3nDACrJNGyBNI1z1s32zKpc/9VCMaH38Gq9HzPd++lE1HTYd63su18Hq7hs3pzqjR8Xizclt92Sm
eR3/KaFR8QEXhNscDqp0JQ80Og0zq+iqcaE7GqitO2UrPtWqLj5SSy84doFHxoIq5O7PtgXYU+cn
+iV+dNNuex9nUbcCVMykqjKeir2QCgmMYIw4bv/EX1fKsdN6q8SE0FVzblHr/pGx+V10P/yM0zpj
RaIVrAWTWZFubuKlGBVrtT5ZVF9sAYIvbezYIn7J6OVY8QYPB74bS80stECTH0qJEmdkddwCFLZG
aZZdvnMrOynr2h2QvGb2dhghg20iqa9+w78zRxAryk2UZfcGcx0Bz387z0M6izO6n+Pw9nuhnYXg
u6TmE8iDC3Jn09Zi6RG7r85MAzVeKLZGXQnnQZiawB1XV7XSBvpT8GwyXlweg1PDOOjebpXUGCNt
D3r3NrScUsifM8jJtn2xRymx6W5Zs7683rXDoCNOmatTS97pwkm89uHtDjclaSGJDyZeC98vXkyA
qHoY7/+GTsknTLazbTra+Jc8EouKxUMrkdaIcztWDN3q0xJoq2yiKyFGcY3w9gZQ69fwdyLeJR49
vpabJU9q9rE6OUrRx5IZepykJcQOJxQntOuwA3L7cdjdfqW9dQPmShXxue3rYtyZgiPzUaSVPxHo
RR9VwdBuOeOeBUjGtmVWJF2H7uzmnOeLtN2FJjgZ8qTSmeqKkOHJ076Oo6BU+5A7D1sAJRDnhbj3
EwDM+kqe1BgFulYvaejgrpADxcR1V9Bky6bpgivJOVwoPNUy7813oGNGYgzE80CcQjgkCFi8cSNP
asSZwgnnaA2M/iOZXoYTPTVbg0e6q736VcWsTP8DA5zdwSkTsChCV1dFZDi5Kgp9b+AJaGkjpGsx
X/7BI/9EMt3GoVwxKgoHUvmOoR4hjgKD9rDaCkkWDuP734Co/aIMzjV6CkA5lVBAnHWDOgHaC1OV
rI6MhagOQU+Tooue50yeG5aY92QhrDMdCWXnsnuwfZwD9tFMxvKxfp9vAIV/buQddXrcNYvGsMim
CzEW9+TnckWi7c5Gcpu93Lp2mEys1vjyCcMGIFcK6imURAtTrzO+87yBZimbrXC3txw2rKOq70RQ
MGPmCrV91sVadNC8cLlpEo/KFVrLEhiL5zdeSEWBfwT05bk1ppfBgIGR3DNzyoHdj0Jzs+ZJfZyK
uOOfaa/0G0Qtez1HPDtU/lqcnXbPubWb+b7+daVOrLM/LyWtwyji08f55jmPRHbCH1QEQs2GfUDy
qcVnJud/k++4MD+1khIvhTvbxJeeMSoNMAmmGgZwIsr5muTnUevHlWOikfVjJoa/B3xR63K5eK1R
W3Ml/yGFp44F3WJgTTaTydoF+t6U4M14mNx/WnWkJxNH6DYg3ayQn0jaMaSNQzNErLqUq1UVqZTJ
6S0oIyR6b0x0SEe3BSHLUc1+msEqW0wogG/bJV7Wwxaxp6h/4wKk8rOhqxrASFUdIvktBY2GaRnt
zkuEqJRFOJINJqaWG5QdNC5xuZiK81NDIrZVebDpWseSvpjcfxpk+MjPMt7G+8EmOctR+LPmtSj0
qOXCYUnz+oMyA/BMEN3BneeUR6V3HC7TEb64Ub8rn7/Z7AkHo7BsJsK08HJJHo7EZpA6yDm9ATFf
pMf/WMYbHjXyPCI7l4USXpwGQF9ZhvBE54oGb98BbA3V7VA+wGxMjy4Z19wZHo9InU7Z9QwmjIQN
ck2zqYTmnpOl7Sbmb0BPKod8qAGbOIcYkIzaWwVdideWYCH29tURk4VMaGZsUxP4/DeM5PV/GeNz
S6s5Z36AV5atfi1U4NktCRupcq2Qh5VT168Gl6F6Dk6MoGRckXBWyJOSVOTfgjfTswEvGHqokYXy
NMuueSH4WpHvNyFPogHQ98tlfwTs4w/WhYpSrVoT0jrNqjUHsOZBsF06Rdevii7ihyipZHs7/bzc
3wEbTzyZxQWE/wHVuP2h4ZewrAoeG7ibDMWpJ9z7HaMS/sZST4pFQTaRzghlP+IC/UsuxptlNCw3
Tr20mAPHWYjXoP8kZQH29UiR+EcP0x84THTscQOZLK8ksuw1rnJZ40E05EHRNIW0DmnKdB83Hn9A
6HBZB0AGmArw5JWP1T9a0BfxlKkj/mziaCgXS7t+UVR8nhkG4Q6+KnS0KCLUlRT9+hvS/PrQVDWV
z3loc28kFjtetNo/6tyI8M8HhDJzY1ORJmHnjPWb1+Vl0DoRmhtxwDIhLe183xfWwbPF7sJf0+BL
KDdgeLtzXq4If97e6tEllyvXuTf7UEsSWbFX6GkKfuz1Dmrt9ZpxFQXnn2653pxyo9P+CIbKReOT
0YTLPQFqdFt+2u4uew29UDme2he3fgCdgYmvByQqhUpCnFOtSYhbhE9qfakTNPBZULrMCOp8AtJS
sj+v+9mhrC9em/Vt4CUtA8k1RZj0/C00QAK1FTouC9whbz/trg5f5Feed0owwDvhZwSVjAlrB/ZG
YzvKZG8y6BSNUpHZijYY+jaqw7QXO+/ST4/QqrcYDgiJECttCmB+0p8IMcUSU44kktantaooiDjL
XuGLqlQD7IDoa+bK0obxW9obCr1kM3zOxMMkg1cXwpLtIcq+wbFvoceF/b5thCqOKfRGfy0rQPxu
1/6tOBlnbL92jJ4zIWP4bvJU/b8M1s5bFFvoEkbKG2SrdtofHhdzh3mYKnTAmIGUViE3eABpAM8k
XUgYOu5Nzva9sUW+8rZkDAcg4qw+0Euuqmaw1g+JqbMNy8T7wJZP5hCkb6WHiXpr8C+GPFWNoBza
6TC1zFc1WxMgMgJ78U5bupgWenNEDEBZUR5JqrkCLJl5xM8pfZ4QL8Qc43n8qIimrdCfMdjCH3Ov
yaGHerqgLiOrhPG8XQ/dPwR8L+3EqNkOh1ikSDR+h12621ee3KsWdZoOc5p8tXSYcOCJ1IztTsFn
h2FDMuPhFwxi3oRC2C6oHrG4oj+Ge4F0tnu3XPJDejMqm9XMXiezrHbWoW3PnmtOTZuKPLUPR26m
c2SiiGk0ziyeETqC0/to43WC3ucQ4sNXV15WGOMNGyY9Tuw3ixqXuXi00FhkGUlzOZVgmRxAuf1B
NAPq3tOKgOUfsWL5Uo4JtcB44gLno/YEFzAgnb7aoqiMFtJrnS6XQm8Q+G42wQeAh84q7ylAYQxq
SkyxqcmG/osAWD/czRKnvyCRz10pWpzJi18ilHVwBq9u+zt7dYbi+IvFQizw2PqcNuDudhJ5Q3/U
I0tfN6EnS6lksDYaFDEEmuU8ycnKFSg/8OeKM7zsby6TRPuA3AHoKp5wZFgy1PUaOvqJsQ02FNOR
iwoUEqz6Fm/cDYBKPHSrJ0jlEjwZVBVaJjEgTrmvU+3U6zA9q8/bYh62As6hwy3c5BfeiBLKgAsj
xysb49EywlDKyroJRhOsM1UVyt4N5l3BapBFbEQtwMwwrKrWZ2JEzmL4uLNUzoVgGtUmPjSeHE0T
Kf6O8woFjasB7nsRaycVVDeFMJwQoWTU5QpsPmJ5q/hhK1MXFtXejljO+Oz5JKww3qdpwGFejt7e
RufMXsPW48AtM7itr+HAvVwW9BrdZMMC/px4K5TgB0Rh+pv4lrGjYgBgEwonxr59WnRCO7HjJwFd
ms7/fCglET3Kd7U38H7UwVBTG17eWLkaUedNKBb68h1Ky5u1TfWukheieS3T8gARwK/qcwLd8dH/
dbTe8QnWauyOGfD8CRqet89vM1GNddktSo4GxtNq20SEayLD+OMF3Fi9URtFD36BNGTcxkNSchAK
YSh1ODwHRNnrwzDwCZRUmSlLD5cXXbIMFOIVmb7lCwLrUDjuccE+jQ5Fs72ntXwvTcYv80jmTmkT
y6bqP5tu21XOOvPhW3JsgndlyUguIG0XedQcAuiq9vqSgkTC2ZLlqMCSHjFMCdmbmgEE1lKTBUrn
As19wvOSgRxHffXBvBtPkBqV/4cgA0ycqU31aF6Z0yXzuC+5hRpK+E29YKUPvAOUyuI/PpwOVXBA
mYJHACdE0PFKuR89GCjB4Wy0+1dcYAvc5ltXuRg4SnwxscClGH5MzkpWXgfbIyt4w5B2vWjbduaX
5Gz4xZ5OCzwujtNk0UtOLiLgL0NEM/DLFwXJ/JeQzUi7bEFNmGJrn8tXjY6aX+5c1qoLh/cZnRn+
RvqNF5XgVSGuh9ezqD2ICftDFPZtDmEYLybB3zzo3+ygQJUirUlybtJ4PepFOYwBCEPBheM2qADW
V2H5W/+A7/nW4Ec52M1KjVTnJYgnf1icd2HUvIz1JaM117EImMBcnV9viOp3I231a19CelOdPypD
/H7E7z4AlkZM8tiw/uDZt3WiDWOAFEwl1UiC526U03xRFTFCrPLpt3WZOsiB7SGvAu7GehucvMmO
mFPOilmTR1BEDrDReHpe1sKTRmt7Jmghr+cNCZ0v6/JcbAl31KFChMu5+aAxV0nj6euNt3RtMzVI
DqwdtHfA5nbAmhiXdIIxtLl2MHKnT+Om+RDhZkU4hEvsEih8w8fr0tLrndltzJxSvNyrYv8m5KQ9
IDyHd0dnA2bs0PJIJ0hxbd2pcE2VGwQRzIxwJYPdfVHa7YI+QItaIi5UbEqVw88AHCkyjt2f/hDt
0vd7CzgyPjxQYz/I1DWBKZ/iPij5j5QJhsjPTncpZFIWty20YeZlXooI+vfJkm8TyZT7/AkKpeWM
94MisejbTaV/eZam5oEsSqLi8xOSWay3Cw5xoQE8rYv3ViqW3HUizEAG2eCrknY3bHO7ACs0mOce
kcDSGgPE2tCX0FXWRynOb/4GmUVA5TPKFdA+/enR2G90Y1eni84Jmwb3vUt7y3BqsMot/QPaPu5K
IvRlXccX8SkN5ZK9FfEmEjPI4dwqnKRYmCurwSanQZFMVDer4USYM9vnVSn7eSLmIc17CR1/BwTM
BWHVJEtHpvy/AefJnE7LdxRM8lAmS/33vBBsRrCRY2YzHD/8KGPlKJKNZ/yXE0ZHu3htVKAPcjf7
1oiUW44USuJ5C/VSlmkSf/muLjuD33vAskEfP4JDPPyPWvBnhslSFGga9wKSNvQ78pIfvNKvY48m
Zd8HiWNJQw5njSOdwoOGjubVHDlP7sJhECHc3UyxZO7tBZShkq5Nj29pFG85icng1IYN3+zlsWCo
3bjCWFZxC5JbLKI3So13skg/d1vuF4dmvLVlEaGxCZ169g4Vq/7cCysr7GyMfQNfk7/ipjFW8Jhw
upgQXuiyETyPEb8d5t0pMDOtRG3YFoouFad5gIsG3KiVLbjurxmFP6vszGDOfmy/zhW7FFUYlfaN
xKIa4FKxfTgLiPzeg03YdbMR1wM4x6rThHPufx9LEbwXcNkF+SpCUNyjXF7jTK52hhlE2cA/Rlm0
cN1MLtq/YJ6nNRLGdIuez8jI+Ww25S3Fry1Fm6BIHTLRPUOt9c5pd/zodEAGlAGEJDAlzqZxGA9g
7Ot+wKUz1jDoT5MyjKXtkH23eU7Df6uHb5nqGTSuPk7TDKB6TM0Vu1bw/d/ZGYCqtDs2i2XeD6rx
Elf2Z+TnpDlSllGhXobscfCdVg8eqIdLamd23plD6FmPRz65Ry1QTnZf9fLZhEhTT0qD/P7nR5pD
911mBt2iNp34zVOBaDef/QnPTK2Y+hqjHTqHITgSvmsiSXZ4YSABtNm83bmx/t4MCiHfyUAR+F64
LfVHc3Cz1zbVPf14ILo/Sp0JKaGH6mnlD2YrVLEkMdG9C4gRLuSHScQUUSpSuFq8SWh+fvZbmbJE
imWL0/c/+V4ijzQSOYpuaCiQWdkMKtiy/htijg2byjwl58nuRhyVtiYAs36VolTlG3k3EUY5HHNe
vhKSKNSDtUpCpqkaKEFnjS5qcPFAZ4YihNFBz/nVgix1346yGBDHsMwrCKiOTkpchLkDdAtbZONB
eCbKs1uS+8625gEH/n6pzE320aOG1jK4leVl5szOhUUhm1s1uvvUAX3NB40cDvJ8NfvrvXZreqSm
fLvAmjxh4sqBT6yEvxnXAN5+QpbJ2HsYy4v5Ur1ukKH1IYLVeEemqfZMLPFGE7p4PvLYu8ucSz4W
ykgLU6+k0kNQoL+aRX8gvo2U3bsM9QknhCukxYnTwivtVcZESxyBQJMAHGufLk0VzXTv+pimji6I
eH8RlhPtm1oocSqqh/RiSfzz5WVLM4JFFGbdnhzBmEDntW/pcAZBHP2m4T/GdMVuYlh1l4+ZJisA
klQgUG5EYia9kItmyJOa7txSDgATgmFRtv5G6wcODLeQSNwXylCZ/qWHSLg6wYqG9OvAhjeahvMN
HbwdmJrMRJEnfLtzX9OgbTOqa8uAwUFlYxle8y3PDjKPGb73AR1j75rYOcGPecuIq2hdZaLCwh0S
e77LoqEmqg943YBmuKhzVkdvWhm163hljhcvyRMpG4R4xypaxIy198UiAmWNJTQZOUHdbb3NgGxq
FeTcLTRAF1ZKZEJEvVWThRBpYWigJSVtxofMR4yULCe3XQ6sPgw8CuH5kN2poXxeu+rHmCvKQ1oK
CNB0083AYIlx0vEXGMfEdFJlzx4m5U7JknNLyryITNZb0c2hfaKYYd4atLbCNwaeHaGPc42EYxHw
bumqHJPkLgH/xjIrquCKROW+oBSooGxiuL9LCam00+AUs+p0QW4wIIrxBJ4KkjIyvmyd8On8jFim
PaeJeKj7vffXiOrKWBl0QAo2+XE2YF1hezbVB9KtRsl7VP1UcUeqEpfpq4BuEfDk0oYiPkBmvope
1qYPcQKsnUdgyqbKj2V9nwDnxbPJiZw9hddxM6HKXsxF6bHbMAuiWwByzTng0c9WRZVRmaa3mkni
U9F70sQ9NDwvrwnaSHLSg6nl/QjqfCWWONnP7bJR/y6kj2gagLWzp1FLYrjiawhyMlfogbo6Xhw5
+xKblUWojhmk5LhOSn1V1ttrUze0otOAQBckoVz7tbiLgn2BvQyqvEAuiK+DRCb8FQ4bH73vqCXj
dsKySj5KAUrCQ8dEDQ/JDvyAwKw5XfklXZohh8jkZK2j9rzAlO+DN8NAGNExoPB3lkRl6ABIpOls
4g0BiSsVCnRXN71cXitAjR37AJBnx9H/JrtRfU1ssZxifXWH+yhpvvwYci4vKRVSJVmR8Kx8cCRH
cZuF4Q2W9Lg9dXLONR9R/9xf915xVoNr2ti0zDUZylu26wdVr7xe4x6ALYmXRT04deHxRqTzbj3f
dIP7jlhbh5gNMygO2dPWEoo9byOQdggKWKMc9MgOZ33NW34GmcxhH6hPP4WuO9m6S9h338/C18+X
412IXg3HCHDgzwrQvGNIlBOvJ218Aetv66GngDG6BLGrpTfmXBQ/QG7CZ/FrbTXmcwoiAFCRCbiL
eLmVN2/Zz+R45ZL6rSDvALd8a4PCWFEAdP1mzh5diBDpwJDvQFgptiy/55dUl/56nfe1KWpKYhf3
oZcNJ+pheNkNsqlu4kZAttRefv2ZpOCLMESFbyXZm61GyGC/iVGlfX2xS/OqcxUUIxvNRN0zFc6e
iEZAC4h46m6NAk7yxTDBiD5PFkOzVEzEop9nqirHF1u1VkvTI9qhLFDtSWP3mOfJHPshu81KNyRL
H+8fBI5yDkBs6rsdfm6DYZxGSmoY73MiL+ECVn1dg5X1ijEb0e5iEz2JdhrFSwGTpOJa8AdLOEO6
CHoHlvgtSdStmgHOPL0vaf8ThAhHi9K45ocqIHYcv5gjr/WoD7j22sNtw7tdHh/cy+8AXoW1yAxM
LZydM55a3zpNWsiDWlWZaeVDtovOzutNUX5Wb/z4avY1fclPlVFHzx5NtURC6aqUofrXha90sO+M
XkUCOWV0sDMHcmIUBrEKxWsSLqs9i/aY9v4HA3mS4q1Gu5Pq1NgczWxgdWOv/x+UrEdgh3fN1UlV
jpKnGqsj8Emnimafj60ZkTvabSW6dhCsKmVillQLtV8Njmijvx3aTglOCSrJinQCafqH+nhlmXgF
KsI31E2Dq0NWjxCfYBgSz7nh0KMZ1t/luotC78Zit4Ej2eJUa4x+t1ALE8wzcc/xJt8Va8Yh9CXq
Z8iN1N0p8VhKGYg8cmbkrj4GawH53sq/Bqtm/2hDZCD7w1gBcmxP0fG+q9ki3CO9NGQW4oVD8YP1
HgqlFH8C6LisuhmEFTxhuJ3/AsNsaWhwRwzwLjHwxyRgCeAvjaXldgVsBsiDWbE0P68aZ+Sa+jKY
O8zlktGsZ5pr3ShfTlTQxBi7GKHwFhZTdrt1pgxe3hn+M5cAGwHoUiRMZRjPjoqwAK13/CeL8Z14
rq9vCAREMk1qdQTA8N++Bp68mf62mWoCP3M+/5vp7bWd1RnxNloveWtAlppU0IwY5NU3dRHf1kkD
L6Z17tDVuS8xKf98wy462IyeiXNJmlmSOAJYIH41rcjKH39D/tIaMo5ZYe6KitGHjvlwE99JxzyY
ni5RG3l81bT/GQXpmKY2MpLt7VO4oLQC76/xrQy5ifgYi5WQrcuR09/3Zpi4/yQeAzmslm+UGOz2
rGzBk4gA4kQgJkOTNphzzOFIuc/7A+m/okH0gRqfbl6sE/pQo0cfBLLl/HR7SM/ycXJfv5Cc2ThD
WoZ4WVckmUaaee1hsCqLPlrl44vnEYKRpSRJEx+jkLFQnL5HMMGNJtC3a3+tJN1eS1/xM5cegxkO
0Ni1HKgHVZ+TYDgMruGQWtSG7ouU9Etz4d6ZONV9o0XsTJq5hvVf0PR1Qi3jEMlSqzudEC5zp4TH
ihYt8Ch35X07JVYNsloThLIIcFDbP9/mtHIZ7vjozf0/ljEO5JjvjQwC26HthSIalqg1ayPVf2J+
KrOoD+Bke7nfi/YHDwyou70IZPblZZsGgOz4yGRF1wt62gAERH8xXAcIIswr8R/hnif8t7SFf4K8
2wsdNeFTEWdkWagO+jKIp7rzyezeQpk2p7lczUEBhMxFY1rDpjcLCS67+oAtf5u5nkXMBs0n5hu5
wyn40ng7sPcSegcicMznS8Q+WM6BoqLq3y0WFi5r2kd/bpnFQpDvJpnNwZfrh1mOu+t2/cL6vFie
sjVFRRivzx8BXVyYj88Ok2/vTnLpmCXJgsgtDVsOFtmZpI7Vi6mjFM9wfgpFldlppDxkCrlEGdt9
BE3SwF8O/o8YnttLvCWEqRSddxaCAf31rV3KsYhSD8mvxgEct8o1dpXKbY8QANOMOpG9YCxlXv1+
Uq2XAkLUGASrcrK+0+NkXZ0Jk4UGYjpuIDnE9iFEeG+9tTK7LZEXZ6RPMsDzSaAv4CochfbDvgKY
A52G7GRmGhFVx68q1BlizgZ4NO1krpXd40stZrLn6+ow04Fpv7PC+EsD64vTfQfWOrpP6wNE17XA
QzUmfj9DiOuQEYuHPTlk+FaAk7Zq806qzbb3oBNJ2/bPwaA03hVOjiJYEugw+TLFyfQ3HiyNlMrH
lGvkg8ga94J3Nq84aTrLGjOa2/xe7xq6zk5rqb8qXRKZWCAe9B5ZqxqXQRg1GeRvWz99eoaFtOYW
V2H8nX5U3uoUKP7bpBBiClr2ACWXvv4Nnd5s/j0hOxApR2A+HgrfMm4HoGB1liIZchdyE+L3xXMm
CZniX6ogTqfjP0J5oTwQnpFQwk6zmH0A+v5LyP5n9P1hTM2LVAxEskaFsx73Bj3k5hb8A/sCtZZp
lj4hvAv/eEVn5O+DFkziVsfGrAjdxX3oqDQNre5xAfkLGWLCfG3hvZ/GUVw+Vey5lFUXUAnyl511
+xxeunZXSCXvnmZ6aQLy8NLQt0IFF+XKpx6ziELiEchxaO2g94VCdWwmtFI33VSKP+ykjxR1W0+i
vDD8M8LKFz21S0BcVMNq3q0aHnp4JzzOxNrhUd9z7cxVQwleQOmbFM1+IjmPsmyrW9a7Tew54K5K
vrGJEyoJZQDfIh6Hi+AKW9DPeqJpWOuUmGsemOMZElne6QZ6k17iE7q/Wyaa3io/rJA+c0b3Nhr6
O3jl/q7dWKTIcOl32DZxMA4dg83zp79k1z6auzqa2hpe89R/uVWSbjiK6N9So4G6D7Qc6CNaiF8e
bLy8vknmQIOQ+0uPZ6LgVM+hY2Kx2Qe/XeDW+I738QLBT/QT+QZNsgwVGx8iKhbaAD/xfG719NbD
FI5UCIE5Ttmm7lVsCgieyoeNeVPbL2/6y1EXammuXlzqQefuwBrVc7Kz89OCKgiHdyRxp5cTgOdk
zGa7dMEmplJvwYbsPyYbxX6K9qY0VcDwzGjdQChpdVDOS+q6MR6UdEJfwVZ35Q6oHd00NxMWgec8
0fzWLth2naWjmIf7sBWDDgYis34vICD82f+6ZRE5SVO96ahP8E02rHlxfwVnu4TtIIUbLoD6IXj/
poyIXayDw9aAwmWZPrp3nxtw9A+RPkxEo/hJWoPD/FAB7+r50kcehSGCcEsUm3cw2KD7Hm8iJWOo
jjXpsUD5kXA4/yr6JVSbV0OzGhBjPASOKhR8zzvUt8WiYgCCCOoDaKv2x73ikUXhhj5HMkN8G80G
Z1NaWbr/kNRuNgLqBQRNhYTB8siB0MJ2wOwe8Byp3Qjop8dhBvkfqUhDVn53tYndIuLjT9Qv9zZN
YyzaC4hCt7S0yG9Y9fHQCYQRdXb68iJV/awIltWcMcYl1WYduls0ZgWTT/IiHB9SuEHmkChzQ5UO
ul5yNJna2/7qUsIx7dB8L11zYvGjgElzxczPWjjQoChoWtbKMGtsTqw/fqiyvw8pmOhyt7EKTjgb
gNrjEaA/49OjgKDXIEsoOegPmYIBm4FX+CqOhurlvp3ldri5a/yxsLJbUM52GqzzFwg2zp3kAhc6
4X5GDOTT/CS3hSg3IC6jKyc1qAhaVZnl/SmTPNIXSJjaoBDwhzluPNoqcs1/TO+L7Cp1DlJaSv5a
M6Pcel03Wrkob2VsiHIS/gVgfoScQJtmUvHSWPnv3Zd2ULN90rQUWYsX26QreYwKHfGLB2/4NqkU
+mLksNJjc0YulbWVICwdyh9jFJvKj5SKVH0w2UJ3LVaa18o2m5cSnZ7bby2ra+bELsLGvSTOwRyy
5bUK9BLxdCC3WJo0q1Snw2c7x5jkTP5apPNxDlz3iOdVygpZQKfF6SK0ayZWKR4/kGy0bXyfWLoq
3gYaz6soTkyc6k9Bh4nhwzksU/Kfk05UKKt/vbWsH4g3Pp79lSYs2EL+K+zAxv8HnggEFzZGrfrl
ZVpOXLtl5aoM5Ou+EzaxAnX9lQltElMfeGZgMZJUOKdImnQPXim0lBTHpjTnrh3MPwLDsP3+e6Ri
8GXB+QJ7Fbdfiu70cmIUaEpWi0/gUnxOp2Hi7T/0XI59SpY1B1Sw2u0VAn/lRCv+PyG8lHxomYP3
OW0S888jsdNiJANuWmWhQVf1omPXVEBdc+tz0OZLoZGeYakpi76f7I7u18Esw9upqSk/8990t6RQ
vilHSbn6Bi6Z014e6Cmo21DJS+zwiYuGyrEWtpHz9Vpes8oU4HwJrOCt6g3XIVG6qauXGvob3MQU
7HcrLVM1FaW65RYrldPgvLY7p6ODwsTYtY6r3KruqhHBHGW9wwWIFUcW1ZfGjghEFw1tGpCc7G41
0hnQ0KVzn3gB+8Bb7/3GwEVzzNvoJZAPLXnu0bTKqmN9xvxExy9TFdb+FaaCGY4wo+z8WhxUDrp0
nqUfrkE9q53vW991saZgMvTOfaa+C3mqtn6FbsFjJe8MRnOfpr5Li+IV95SV364cb0Im8fSxS+X6
rOAw+FfWfFYFyxhs+pPmURxQG/6yEuiKgqvcx5GGRL+Wtcq4cId5koRs0U5QKYqtLKBJoSzkcC1z
xEU+16bnc+Qq6bYGeWXDtiLJIVWUU1detIRrU6o3LGDdE7+7WnTpJURp2NpNZ0LnNGraZERbYuzz
bnfOzf2uhEYb00WEsH3QlA7jlQpwdcdS/RDY+6Px7orOqiDwNSIUDeqbDMG9jqGdtewCtQdR2yIM
odrCSG24W8Mhtn+H0GbtAgJlXNTRdcG+nlLYmgBMhegAjlbP+7YIXCVLm8iEwoShx6ZNvlcttcuu
VxK27zuyQbwcDpVHB7W+ZVoh1up0P1kWjgSubSAgBcxzy5pO8WYUyJH4bFhievvv+VNsWjw49skQ
FJ1PMGC6gkqMazIyqhb51qadCjC0biMOgEEeBhopKOKU9eC69BKCq3kynGmIrJLzQqMVP98fBK3i
EBh2f4EIHE3wTD+p1x/psVvoOkFW3B/NgQ8Vyi59LUP78R0re55fRy4BCuNFkEgyjKxO++3qsvPT
Ht2Hh2HgmrtS81aabl5tOFYCknETklhCJqHNU5UH3n+0KIWx4suIP3atVPPAR5xMMTgNWERh+REP
hmc3jke8ySnYwA9XjNeNo8JYnM1fy61hH/wzPT21In/DmmCw9ASiGgiP2CCK5H0swsy3MUu/OnYg
En5yqsJ10zOPqyouQJQ8RJyo6xusSa4rMeeRsKO3Fe+IPMH6s+I/UwJ3PNxONK5UgD9uBdESi9jJ
n06pOs++4PQwieGGm0IoCMSbAk/93bxsSUq3MLjKozZKs0Pj6wswTi48qrR0CwHXdvklrxFTN6yH
06mjL5jXF2jc2UQXZL2a8QC8YJqbCWTuiAc691PT7ROzBlwXwwSVh2nx8JVaofS5s0yMxzQlKN2Y
1RXOU17AvWf6jvgEs8MXP04K9k5x2kd3MVUedxXKkIoy23Yf/DeoyPOMtIOE7j2oM4nSCokq2aXT
4BSpmgPjfcFOvIrR6SQo8LUC0nDq45cswg3cER9Ju7rMolRjZPB2/XOwdXf0jZ/JOGLXWio9Ue/L
w6xPaOaWePF7nBYQxu6c6pbpZ4+hzOvMXYcAZaGc0FzNx3e1Xas2GgwGeaPsrgkFJfjFUNATvghh
zSM5gELYzRkDa2RicctlZlNb66QbD41L15Ab555eJo8DA6TAy64dq28Ntgn3KSHppxUwbZQljX5R
17TYlfaSY9cd5RyUz3uoL0odUU42qU5b+od4h+4cberXkFOrczWphddIMcylfVwVlAtkqlJKsk/g
fweHQhawPRW5Tr8eHSwpTp5OPCviU3fivGI7G66BUYI7+6n7tVYPDOBdrXn6aOjLpaaD5eOdbbkx
MRNBIbeRzjDgtzxhTZrdecECG8otFeI82oHIwg2ipvXZ2lkH8XBOXkXeIYe43wPz++uNHLVBnL35
PPhosuBjyGZxKayF79i2Ro7kh4XSYSYSZaKLYtwE+zATjBkE0V1rbgEbX5iFEjePjqJm04EmyLEw
aw+556xVQYK3EnX0nIRnYboKAtES6grWQ7hslDAY+tY/yaWJ6HTkqOCG5iIDMWw+9I17FPbZt3S6
1YBO7holSlQ8+Wbv2x9GKpKJTfbRTX6MpOBcLKb1HS1IfXtt57UoIuDAMOlBtiCRQcsfltKcb8/k
TKF9q/PLog32yQQQCWk9lRsrb8aTsbm9ocue5hLsHulJn2su2upQNnWaCk4eCTRwTwWTebLD++Cd
tp85t6N5Ejqd7uNJNvI9QijruogGyraRB+DHiMMPILfqkeg0QeVLWp84PSlvwiPJh3q3XPZnavdf
pCzK6fwRRf8xpWSIu/sAi0XshsVO3QcsKEAxcpL1p+EPDX/sgLjgBF0eSNNlvMldthQc7/4U5M4Z
wM2ewKf4no+rQR0HMa584wWM5Pmwy1tzcwNbiepY7BeWsJcrfaWqS29YPev3DsqVTPXq/rAZfSw4
oK8wyPc80X3zj7od7ki5hkhmeL7wQs6+JL8nr0X2+DMqKsVhziKI4jR953Mb7+cmlI2DnyaAQtvG
wFhzSZz8QpCP519UvFuWm68n34qGpHOE7iNNX76sndTtLndkxOOh+/R6L5nWyNgQ0nBbDWyn/Kzc
baAzS0+l/1+tryf6wJy0FCrCcBq99yAt/blZn0t54qSoy9h4vYYd0lnYD+uX2DFvBGbqKCEcr/SY
otgN8ohU76xGrOP3xHXmcTKtPoMJt2HM5v195wmXUev1t9IrWo6ZyuZVy8wunH+RW9qZhaKUQ3yf
lOmf7we5HOoBxW68NmYFovrht3Kdnutsbxr3ohsu8RqTRwXhpAbIHPK8pRpJ8TnbsnmBSHzxI3Is
lrR/JG8kSn0vQ2sPCLNp/TBUfygWutmWavq9KmiTnnC+ei4fwYOKTCEk98s+SNIJM54EMo11kjwV
2FnFoG7TYX8BKt2LVVQLk3YIMl1A6rYcjRSxnEKhV28ZKWqTYVB5zqvyWQrLQYKrm7B+8BVBcmW7
rVq5gb6FewZqYYvcLYTPvd/w8XESQhreWnv7tVvOt0YaDTIydDusII/oz0UxdfJsdvG2vQ10tDkf
QtxwM8J2qql0DnuBZMnRwt60UCrmNL4XJsyiiQ+mlf4HQLrael/KUMO7QaY4hjcWhRFaaWyReceo
E0o1A5cgpBXIrurfkHMXftiSGtvN2TQDX7glf76tL2QhK/UmuKYihNHuaLEKR+QBFCl1aZ8taqUt
1nV2ceNrxgxaPA0IGpYnoDSzzZKOVPdE+qouMk4xc7UMOfMp7emWhcAnQUn3L0rPq3ZvaBiQnqCf
0bPrwTa08n1DgQXYNMnGhA3OxJThTe4UPt2gPbmhb++zlo5tXucDtytIBk5CvgTKRATza1Luq/kM
orBKhhyYMIUEdR8De2wQdpPYDMUQId3J7mB7Imda6Q1WcvFmFJR3P8X3AqxKWgNGl1j7bGsLxsym
E0Iyv4E3vYgebCVmwOt8VLAITqQTH2BojS9f+gk5s0WKhV2pkMveo+E4DQcBiM/qX+iGTKUxMmEj
CJ3LZ6Yy4t5SSakxjsTgVK+WeveU4T6HScuMCC3akZy6WIo7DtShrmFd3Ir9ovbzkcLvsyTW/uEh
VRt5sjeJrNpTpFXTrlBTMbwc7cEHjTuQFsGnbAq7LZoEgoVzNHQEPbMfELHsbTU2NSQIqP2OjHyk
JJsLEZBIGmqku3pXdP5rBoByLziAbTHWC4JIaeYujJJlvTLpBmWMv/PKqI6o3dPmPe6742K8hIzK
pt9IU7KX2hD3v4ZqAI0RJ/TzX+E+7f7mb6+6V1dtSrSNv4cb2PzNlKovKkcyEFzIRdfxLaVn0+H5
N6/YCBcjR5dcnjhyHARcyd6aTByf1hOdzzWkh6Y+y23LAF9JeG/YCeg4RnbED3DjHOrqydufPsST
iTHzSFNbMMzJdK795sJzdiqyoP+X2WlIy6OFZ63pq67LT9PGp6FVHxMy7Fxhs5vRCrzGq/MMgBNY
1838ANtbFF8Hd0lxTD/3ZZZZldV/hZyYtDSfCPcVrm/qo2AmAyfEs0TSsn/V6ThEYq+VUJc9Q+kx
h4eTb6osv/8DKWC1oOUQx28m4Fk3dknZL/yXTbTaAi/zHNiOGTSjBcwpV+ehBJRCF/VAx4DjGg26
AVaAit60F8Gq77nylHkZED7LFWpeuRSDdCXMEi4WpUbf+0c/LYmI5k3YcruCHi9hpZF62MpqVVS2
Ex5PzrEi6aWgOv0XwnF+P+jTJ7BO7ScTyhhC08r1i8UAjVv7XmaQo7BleRyFn+ADwXdzN53whPHY
pkhAeEj/G5JANrORQw0aBAEZAz3MVXeSQ9V92yBaLNAHf6gARwbsMNBX996LYPqPggPzDJ7G723r
dmD6Hac2joRVSckoWWP4BNPzQiwiy+YhzuTp5WOfHizILW/9fJdDXJgqRSLM8a58n28ZTDe5Q8mt
NgWjeazGBeDXJIFvHFiNmcjeCMLI7aeKY7VcjkO+c0SwymAU30XM8micfpsYSjA+bZv+RDAVET71
/DaM/xS06xMl9V68D9xMfKRbdVIdv6RDvIH/U0TKQnHC+RpqpNHxvcreXhdMPwnfJe4z9vyqPmru
XPikemnnrtw58vYafxc52Qc06jCnX6vr0DGU53BmGY0JmBEUudNsAlUt823YhPXM5j1DXy1Gjkxi
gVFS4v+hJnyLyZUIhnandmJm9AipSJI1jEe7B2yC6zOYHjZmE2/wIAIVi6JQ0kd1NhhThV2SFC1X
6xt7aiQLILdA5fH4qiiH0fQAW9ullQTIP+CibnLIFSI6Ev5CC0HLovATQ71cXqCK0PeihZWIvhMG
rin12+pmX38WfuMpReThK91wJtTU33UUVl1TMOUSXEhKX6I3ACF8wkHkznDtyc8s32pdDrFZYEHY
d1ikOmISv57RbOInT4d76fSItmOaAV6pcPj2nLE1yH5+H6J6ivJvVt1FJwUTSi5EU39lwdBC9vYB
CAfpBcDOMuZsNavhKwR5mi5Adxu7+mePPFwk0zkWCm1tF+UbhlS8DneHiiS/C8qvRPAfknOBu0xd
ncjyFY5Y+Tq0R/+wVb6zD1mmQlYu1EzDKcsqdTCf1INK8Ew8kKR78eP3tigyZoOfqfavxJbUKDqv
SriKJtR7ysY7cC0d5QbHx7d3+EzHrs2HfctPh4HX8H53XYIbCYLPsvG1GFepW4RybacL1b3TAjzh
S6VJIHv4roDdxlVWFlWPxHRBD+iqeLrNANXsEU+T6iBWO4oO4mLYDomrFLPlIqjWO+3nyrS9MDSb
0Plz4Jz832+nWNFMYv6CB3cYbA2dxYAiLBz9CqHNgAmzzhzhv4JOaE2znFYvbstOQOHxCeV6UEYx
iFx4a668HkazUGAtV6zEeQHmx9cJV+cHVUXBrEAHqWoHc9xKbY6cb7+8k5FtRfnLiBzmlI+Few/X
nUe2O5ALXTo62q5nyucFANuu38s3RZuf9rQtBOdPne/VomR+DI76hnJxn0JRwE7CCbt8D/s2HU5q
iVRTJqqxD2eUOiWSsqIbzK8ujy4qwLgOEdriIrBtRk8Np3B9EfYfMI1eFXEGaMnDUpBFVMcB0A+Z
VaSwQETZyp/hqaBxtSUJH/zQpYdwlsc0nFn/S8aylUGantaUKSxaeHmwmZKGxQkRtQBoQ7u72PzK
IYMGsgs+k01ippX1YAOMaQ+isJMM4hItjxUA+KBdM0/K2kwBL/xGRd/a7+oIAF5ApOKNkTd7V13+
5qi+F1i1I/QhF6gnEy7AhR4AZajLgQNVzts8M2P922K/eJxjBaUBvXXUBGCFXfGoV67nybAOPYc0
JgibXj3xvV+be16qqPdG+uLG0rXm69RTJ7kAHdSf1ibjFW281cE9uFCxobTW7nAPDmTyLJTGxBWp
Yq83Ms+pTUtZwcgilsikq9KGIujjdFCivAaR8h8SCOa++ZyzP89zBhGSOYDPIPPMXzHXQXCuPS6d
8cOLuBmQXVCNmhcv1TQT27EDA1nTgGX/Y593rh0jxKGe+wT4u7Xo95DV6XozHBtIhui+fm5O3lkt
Im81QC30OtaTDLUPYaoG757+zSQJKAJdHMfj3lAxk6EDSMQJ0MyfbF+l2CJxDqmrv7ToiXDOTTdp
ix94AePPPO7fMfv2dSCZKpQtRZ7Qh8h9OXYxeaPkL+mrYjJRFr8yJ7AJqIP5Hx5F31KjHAzf19sW
TtDl/WQxckGewGtAICti2YqPn/XVeRWvjH2mES5H1S6pzF4qQ9CuqsVpHlrsUkU3pfcgP/hLNSY8
CAqQZzmRqT+ey/Xw2S5aDWu0HDXUgnOADpzroFmsgtodBxDVz3cXxaRc1RFdtR5sAjxSt6Aa2vPH
I4cQ6Rfm1XIC2ZpB4YRqsehJ6ZN536pCEtH1xwo4JZPZ1R3ihu9UaLCS38EzoQmRvCTK70tzaDfV
csy0/XeTaCi1kCecoGXroZYtPNhGbazonOmairoAc3Hbkx+2IhD+hLOARRts1hh0QKbb1HrwYR8n
4H1yAN1BgvtmjlEr6qI/wgawRfDhY2arMjn1a3S7j+LdFrVLV7nqkEL01qoNHkxkS/PcQolw+hvD
3aBAZab0eFNLueZAiTDFuE/rVwOMXitlaG6kj9zfuPRRuuZxy2QkiOz30DxiCawni4XBjKhNZLBs
VnFomukuE0b4K+kDfqqwfSUaNJRQaaBornYhXOdRDFmf9syEcuewQe5Bnp4FTArbPkjt+zqrOEBY
5eXXtUWd4D1F0uEChtYmEAaSp/TGaXVKjJuC1O9lELYWo5AMLk8wq4m4ret8C8yIcJ/HM1SHLGTY
mjJ+zIjp0GI+CqUgaR8jMKKTBWkMJi7d7Vf+h4V8lKk1dTB08DH3SbCVibabu1rFuB1mDu9byznJ
wGv3YnZXk2aY9FMg+sur4HL7XtYH2/G5rGQGHk3B1CS+EC6+DixBZ7UJ6YcT3JAozuKc1xRxkfHy
u87vqaWdbHWxBsdgxZhtNoyBvGA51qMbxz42WsMlrAS+LugHEC2kgoha5O+5IksBKsWSBAaRZmMe
KMTvsEWib5Mw0lCav0OH8kj53DcNkSs16HCgizZl2KdTDU/HpedzATL/6RQ4kNcMhkRZ3P+h+Lta
jONSGekXw8qIoRg0I/KiMp/RLdKrncr2Gpobq2g4Wu7+4M6jADU5lcwlyghgtuuzMtgh9Uts1KwN
4IrjsESJawTD1uLUHTHSQacsw6JH3PZ6UzkYGmyyI84wo3qLKbB6vs0vkkw+UHgLYIWk6VvajkxG
GrRq/iusaNFIZnzAwwj2qevGjF1wiALVXAaiJ4FHwJjA+0DSQlyO7Y0AZa/zlvqd5TYUFuyAy8mx
pft/FMV8VE9v07njPnY7ptXr6dnaWkJemdCigUrFswhpOS0478emiYHOpI8FdnhrJbMahgCtToka
Lx20/P89or8Fgn7KFE1c+NKZoOJQiqbENw4tD1gHvJgCW5T93+1kY1XSqDfJSBodOIJsIgf5Yc1J
rtWaXmH+WUhgLNx3r08173z7mgsEh6FXYf6uTqXLkyesmM+P8um/uHbXpKG4SdM1iaHA+7XvNta2
Avqo66CQTqfwmpG8Fwsl7gTVprU+5c23YlTLierD+KyYR66shcuD8MnBUgMHfMOKKEEjUu+u1J07
GDQrsicwGeBfL9RCSncoM7vLGwssGL48BG0q2YCVOdPvf+TKm5IVxg8p7pchdNTRJN7/zfg+TBRJ
/rLgjwRkeujHVx4cZoDc1+YNLXuqjOnFEpbq5q98ZnJT3UGO6wiBQ4kNqEspTD8OC6V7zppzZtiS
UjtL1Da9BsMR6r7gc3sDvmGsbfw5ip3EqMuGGENk2ZL4J22mASyxJng7yGi0Z3LIYGHuiTt0IQ1J
Bza05li51axHreOC4fUnYVwNsS+RA25fNf6lNB3nHLljuaIGMimFl4FPUA2iYy8Pq5jDY+U/uszY
+XOf/Hdt9tVictbILYow/+VUWlK52H6nwTW+FUcMDzaescEUYy9rnxBN7Xgh8f62gavHgAqbZKWX
es6pKqnrqgCqKyQeQ467sqZy4pjCjRQBY6JWhpEvJK3UMfiSkZW9VqMPeXDVF6rJGsZrXByJKmBZ
fR6+l/Dggs0oc8ELqhB8xRNOMB59joszIBdlCeG9KNhoFbvubu8TaX6Qw3+GXQja86+LUc0oo99v
pLo2R5SxmkoUzkQGaMMtAUWb+k6Z6L1FwkuH3C0Mmr1hqVbzmWYvlx8rwDTv/Eusvk1oPTj7ExeA
YTVTIKQi/gN++WaB+ETO3w7Ypt2VAoSfv5HgFuu0Sx/64pSvR2mP6MPv1ZP1OV2uHez4038qBYWL
HoLcJ2tegDSvMxUY4Rcu1nM2pmE5giCJkFJvTqgdN07DEl6KHYV3f4YvyLFnM8egzx6tTBo2gWje
j5g5BOZ6qHO6lpBSu3N5ntsEf0wkz0Kcda6STcRpaBQkdSTtxDips5NFGJCZGuki33CAJqiFIBBE
2fN3wCKsTnxbZCFi/NI/ke8xLs9zpRafjN6H1Pj4+4/lvB8qbzTc7Ev5O555gU7SaU2bnw4oflCC
nDDeBVEjF0vkTwjentB8TkpjPamXjz2c9EqicQYr18lOAUNSXsCwOg3eCBdt2VB1l4P1Ax+D4Plx
+yM/BmwYYrB7xmFLBDdVKVrrclJIG124QcqIsgNCp7nM7FfW9Sjgq8ydIymxUpwtFP5WZofLpv1b
QLAb1sBI80i/6Xol3HmMosZLwbZWtZMiE9ta5vTu+V3a+UyD1HNo0bb11YV3W5yLQ7T2Xml5JJRz
p+x7dtwJmK8c4wSEyqLGPiePO9H+ZQ8OSuaZCs5gyo9Y8qIQJDw1VYCGj0J9KNo2i+A5MXqvTpl0
3+IT5/gPNX3ff04DcfWdvSjOVq19a3IVsuURvJHu7CNPZVBLJpkR1n7mhwhv096527HqSHkV7hB9
Vl9BQjK3YZtWqVOVdU4Xg985rYfOUky4i5l4BZkxpMYHucQatwttAsbU7YpiMGe9u3/l5lxLjpW2
z0B6pZu3FLR3f/o7l68QwNl0VYb8MZNUgNGUj/hAd4duOP+ZfR+cEZkPmlK5WHXkn+dzgazQUhga
TO9pBd2s5HxaXPXA/Qv74+Tzkh8H2dC/eyqgT3kwegLdhIqclMweXxwNkfVlpGL83cjXiZ718WM2
URSbyWNpC3hV+0xXqfmXCi/jh31G6fF+34Pyb6LpryMSeYA8tV73bxuH8Jjk9PSkJQZOZEs1BGxD
iqBfF6kvGhusoLlEXKzOgPkwhe4lhST8hMeSZrqopEDXZkm6vWTLLAPb1nbJ2QHVV42o6jxNm9qS
AIDjw+NoYOt/+zJSDT/+jGPI1PNCcSbsxMMO3WhA0yGmc16bs5/Om+4OiGCYIlyLLdylRo5WUA3Z
GjtL0izPnexLKwArMhDHDvlP8lF+0UTXm0ZPfsRJhUxI4VDpWb7CfAL+Mw7uZE2EZEw6/6HIkBWJ
HKLkvnLDrTXiBsdki4QIf7Z+jwT7gQQTtbKjhVPwFQJQr9j0qlbxRyc7APejBtuZXN7fCO+Fl+y0
w3cLTSjVHj8vXQfK+uQzIawDQgmRKC6eA9l1Do3eWRum/c/jUu24Ajvkv0952PfM6piFhmJabLVJ
m4YHHAiwfKHBms1w7JDeGCQHpuIoLFBPRLOAF0lSv52JWE3FU1+7VVHfCe6n3ETH0FjwWC7mHwKs
SqeVCyTiQ+YyjYM740dD8QY1lgX1M2kLbMeZ8xXs5+XF/obbN4mpdueg3FQ57jhjnI8LhjKrCUeA
XFYRqL+soFpH1nc46frfbEy/Niq0IGbr1tgXfY2IgcMHTw5h/RWtj4szbkobVnZx7TwzqjGoUMpP
+n4QZKbrZFhJVTlaqhFuZWa5BuU8dUH88VPcob84qG24EZRQDn0TcynVDWlkaBA4MKRVjqZFqle6
YTXWsPSoWGNgOFSpbTZuKju+PwCpFjZlCMiSZju5aQJa/V4msdGbeciCKl8yFf73vf4UGm9mFuQk
t5qqVZN3MHJXoTN/la99ACmN2v9U4L3SOGJrL7T7Hjx4YH7neImoK2wOJxX4ul6V4KEiIetZ03p7
LXKorSl1Jf6oz1lNgMjghSlLj1Uk4B3pB8jDMR1tC/a+1G47u3UoyTojvfCdqdKAJKDol7k4Yxgd
yic+KbMxHpkeNPwuzzByaHfAZ5G9Q7GYbZyn8S8WGaat6x7Qi76pjy+HNlhkvo+FcSQkcrx0DLjF
MtNrXqHQ545U2iR1JjaaakcTlk37TmFHwh2ldR+MtIJioQwjLDuC50baOdULQosWeJwR3NRx8mmc
nvU6weaeTu8rflWhWVB7dXOG9DR9IyQAlnezSS4HhiQ8kndPk0IUPywNlN168sxsLnzQim0maq/N
DzyS+L84O1Rv71w0wTPBXZYYuRuLRx28ulYowMh4GVV9pEZIaz+2aDunwOSd1l4LWK5mOf+h8M0p
4/eCa8pR4QAuMN+G6i/OueeXEUwVmXkYmc8dAsLNCjcHI+Opeaoia8uh1h39B90T3f3++LQ9dqWS
1xjzVerOxhC5tUceFEoQ/yJVn+hVNKvIIqFlGAD/whMItduE3vpBegFNGkW8WPGSRmyPirhbyKpz
qjCmKAs37393A43pKrapZoUTq20MxanbMZtOmRbXT/3pOrXycI3GjdMuQQH1Rs6EAn85BoAJh15W
cziztBXO/8JB99vWm17OxSgrm5gmoJ9edLs+OYL9B+fEumtRhopaZQ2Rf6XB4kl0fSGPTAQH3iX9
WhPSY9tVMsgd6wdETUEoNKHCKB0hCeyeIH7kDWHzL8zf4ggUW2JyS6euqi4+xo9MLvc6HJyB+pcX
JbkUEPmjhzAIR5QEmFGElt7baRxxFSifgS1vI6KVVZvVJ43ISn9JBSxrYkxR7LtfOhm4yAk7QZHM
RDqPBW35D52zNJLbmkqWBhnoX569MXQv4S8Z19/1qeYTuhuapctC8gTsR7j58hIBjCg6sj3D8Pyt
QC4iqgy9KGKcuoNllCLYXvJx1PDQ/w66oAy6hIzKOmJhhm5xM3oUgom4UAqcgUYd3vYFd6q3rWn4
gUl3bIkCPVCOni7vF9BpqENyZk1jU9hjbobBiEjnAbHlONn/vQHb7oCR2RX+JZ8gPBEGnJ45UK43
UN5BGK4D5XxzY4k8i7T51j0DdvtQcHgkHtI0avyvibJZkoC1E7BNBN4vHd+l9c9keQgBLNQs51op
qATUrD5Q9c8QFs6o/aY+7+fUNSl8aOpBV2//K4qd7nkV6dx4i/2dNfPgsCXRGqOlrm3FEzj1onO9
0IAxpJZQZss+aS9YQxAmX65nt6oukHlUUkrtyNmHBWa/AUvvp+3nnGXNikqey2p4QokfumjIc/5Q
ot8sTdaYNT9jIYstLtmB5dbz9tVCGVZSUedJPSdqNXoEaf6DULNz50ofHvibD3725yLh/UlRZXMZ
pHFUrh4MpMmfhJ733ksCehXYo1yQiIeAQiGWnp75lDF69YlKmZRq2CnAltxNxvlRYGRT0RxFhFVq
sUp9OcEWVn3s2GYI+FaCDdtGo3yaBmXkE754YCAicZ7hSLvqhY4LchqlXjjNlRBX4S/cOZNteJ3n
hcE4ZOs0JNpF/DYWHOXvirZL+cDdybF3sgbAxT5tVBNUhtOh8SHmkhGqYHKxMdvqVIWFEsuOqoQ8
6aW9oSBtyFwPLwBLldLDItqnQifY+h4zdRPweez0AyenTxxs1mhiEmj6ppMxz1kODVUQUom1/KQs
qahLpAdT2GJVLlnekuaKBJsj0NpPiHORY7pr3+fKOK2AY9FLEp1FLpe027sm7BFTJZg+mRxcOUqh
FYK5xZx2XjWVkj7U/i2/bEDNHRRI3ATmQOOSEjNAfU4nh02VF7MQNEV+F+PV5wwgRdFnufBQtdgW
xKNLk9mqMLtc45w4eCsdTZWtV+5Nqhw9JEXcOcqDlQUEsWhWwLa6argTdb/ad0VNzIk3aM7MJzff
jGcAviim+oSdRFG0xTINf1fuWdhG2aN3bCpij4zh4KR+hfuCOGeUZKVnXXy9z+5DIrSzS9vzUKBH
SzFXORdLkr959zR5pFAKWjYbq92hdmj+o2zOTCorMUp8ptkv0NzgqASUUGJQf6EoS4/dWP7ciSsO
rltQ79ymge4yiHdmEubZelcfu505vhk3nr8uVXJEmMGNBU2Heer6OCVe2k5XYEKi/pnSliPnlEp7
BdDg0RP10rrlfcfg/lTS0NH+RJN2QCKbKJg7s7buQ6onXsslmRBn0AoRKJ+KUdA0AmB1BbVTyQ3L
gS0iYfmV5kZOQXpSYBwo+v1V5G8D/HNwC40bqA4MGQEpKaupKfH7rb5BRV03Bcht+P0GT2/spl20
yLgB+voC1J3IY6ZqROJmoyTfs8WalFCnB6cGQ2CXeZd6CU1cDyQkpJGoIFzN0eSTOEwX9Whc1ybg
eAMQ0fzLyBTkFZNKLMlJguL2pYZJshDBoovLoJuK89LMXKGanWm3DiEq+IE6zM5jxpSUjtqIe1Py
gm13gFipgqXKhVGZGQde3HbFnySTEhDq+amS3xKVX+IZTdBqJarRxZ/RRI7L72f+kulQRCQZ0asK
XCtYIJq6Or0Xb+vJHW19vbB4O862lnkNtSux3hShYe72dVwsTc78IiIleYUV+xfkyvUzG3xzPput
r0NKryekOdY2TaQcJ3AV3eLOYjscFkZ6e9eKJoL9yjhDLhdlDS98eaMtzZOStMmg3g0hLxP0tA8w
f1d1CjyeMRC/s1LTzSb0Yt5XeJGpK3Wl9JaPZydKxhYrwCbwgDaqVfo5GgrnLQPmn4Qqc4uY6H3f
NjWFcmxdyN8wW1izMsvvbkVpQzyIfgc1tPOuNNe1AQL0tUgzGfRPJlk8Wx+4DI5TlPWCOD95xLeO
W6vk3AI7EeSJHnvLPQEIY7APR8RRkTmKQaY5ay7LSWTDNcKfbwQ1mDEQsF4k405HGxlYl9G1ZX8l
vrZDJzfc2RgZxbJmlov8VXkvY9y8/g/ly7MnNoXGo2a7CItT4Y2gwk/CYW2s44kRKV665uQPBBRb
PEBPUku3Bx7/YWlAM8mlMzpw81hVTY9OgSydL0wrNtDyGYZKDWVj4lmfMnCeoYDZGZpuks1Lvf7Z
qVFgAKt0wIFVbc1dhXmYDDTFrP5pHtgpTMpW+koz0lv2Jeqb6LqbabMFAzRYCRrizEEmkOUliJjH
6llYV8lvQ7fIsAdS2oP58z9y727mZQw8TIhNvPPLiyvtnXRAK5lKh1BGpAsOJAi47MZJZy1sevpO
dGmZxSFUqnMlUKA+hMJ4U9Yah+zGf4a+27BuQIEYyUetYXX1lUgT4ieRLPPs0+DyiZvBZWdKJAHO
g3dpq5syirwNWd17EUNTq4FOFxOy+k88DU3csxkqHgyaz7B6gz2E5zbsxPxkcUtzx7nr9cJi0DV3
RXNvem5KEgeelSRInlIikh8zpb/pR5+pdNHsjQgqWJRkHUmFZKbGFe6UWRbnKs0cBeebfDRsb5Nj
RMfZ5HgsE44rOYbUd8S1Rhw31PomFwEL8zcJ092+y2BY/lse7Lj6JkID1RbWdc02jJaqaUwWrPi+
YRRyusk1d/qQ6h0pzBxt+pX/w3Rm3dsIzVsFV3ODqY2bJnZAGuSqz9+gAH5+LqLgio1wAtUwxj/1
lshnzLAL3D3fOHx7/lxaZQ/5qM2wJojXAg1IR4unfuMMZr1wu9HYTN04Y325mTrYBRborWGSF7ix
WyN1ERnSv6xLvFVfnd3g83FuNR61AUNqxDXJY0Y6K/4ocnee+IZw9p6DuHLCrOMjJmUe/8TSRcZW
5f955DnxxkcoWI+LTsT5oA5A6f8RHcLd2UBVOuKIXsufCA7Vm8yW66qCy7DpUYsPzSc7mgIiWKjl
v3g5WMTfTjFV43psOe9k3/ckJOv+NqmHcBq4wCkdIbnr1vdWo9b8H4I7mtio/BeuiSP+mKRAJVGn
aqrfEBXaS3wDic3ybm5r0t67HwKwi/s5J/ZDxSejMgu6yr9P2A2Uqmq66GGbLZ6FjCMu75qwVzz0
hFCbqmiLoqvnLNObrnvsjp3M4P6tfqprOg+Vx8gQ7Dye0HJRLIhfAvJ6jHMXb3tQVrSc+z/DNaKl
14gpe+SjT/WThQ5R33QpE9QAnmHIzmPX9X021osqKV//g8AhEQp97dKL2b9cHMwig58M89QdPlYu
b3Z4mTxnL/BN+Ic+TrnBpdjTOuRjC+tl35TWhT5HeBZVpfS/XRwPJOQd1kdFq7HqZtGLt4g8tsmJ
ApoaBEjLCsK19PireyADVpZu9lLf1uZUfeUIgpJ1tyGKLr+Lh0rgnHeSVXEcjKLsdQMwYuQBH+MZ
pMOlifObhREo4tl5bVIqn7+1tNNXfmH9nrUwP5QvLs24nai/bt7BA6Y6/mMxkn4O6il1OMXRCqKv
kbT40sm3qIMl/LAXSHYdU9WiTzO+aBSodQS8e8OYi3kKVCo59/agSKxC9v+DV/rT/O4H7cp1QHa5
uVg8nV10nbIz2OnQGx1K/GD+pQ5QB2jD3GekiPHZKDzwVPZa4Aak3Oq/3ogEO8C+hTa3d6HChqU9
wQRB2HaSqTTM1R2NtQwkVmdi2P4tsR1AXQWm3YlcyDS8P5Ntu/TB5ME3GoqRkhiJla3R6zOBUq/F
awsA/x8wnpudvKLVbPPJ/UYms7YyfTZ9Bg8bfz7twFY7dbMNoSdBtMP82bvAJ9mhPkMNEjtFkqAe
ZJbqQwHFOH2w57UNG8ALgj0BMRu/PUdbr4d/pTFTF6xcIGeUYQWgfLWdGmMGJYcz7ObCSwHoqdRp
nHN9oFrukLoD4rkkSoSldQ1B8bxXEAZI1xXC+y1u2hg0x+hyycKF/MRtviTAWKtX+ul7ksfgqc4E
zsTLymiLSkM0DZIyniVkNjdzZM2asjW3i9Out8Rs7fxofKGplSZUuTLGuxLXT43NuUjoZIxRwepJ
sbZ3T4T5YzgKxXD94lhAprUtzTO+t1jWvcsdB6Jya+V5nTtJMkAjL5hw9w6MN66A49yTzCqTkZQz
xik6rVRCL7cPERnOWIoOY1DsOcZKajnZVHdTQn5smiiyvou+wMDPZGVdUa7cLoVPksoFFSULsLmE
iZSPWkAzdRGlf1UQOwM8IUMk8h7Nq0RBj2RjpI1hC70SXSD0WmUl/gOtabcpzr+zTEXIPbHh0UwX
ituKuwgeMq9dmKWdIEmxA/3Ywt2MoqBjDguyOQuHtXOtW3SfaOzelGiu7qXvJKPNBW4tiRcYLYwf
/W3kg/X391o1l4ixHZLEzyJK5eI/DPg1wwNSHlmoO0l3oFFyZajLT8gUrA5KVneDMeMGPd13GcG6
LS4AMX0pTMOI/t68tEwPZKM/uN5LXMV44bb66epFDlcDieQjxyLkNYtABAJev4b9gm0c7b/K3coZ
RbZNRGuQ6yck3uyvexAXsT/WDAE0nLwqAlPSi4Ehw6ADjXuIhvAdOPSxtoL0j3PNlab2HFIHARkG
j8tajHqCYfoyEB8MtF5KeZ4Zhh5So6bdSal32lajFriMeGlpgICBqJXCLi/96IwXq7H9wbeQGT/e
/t8LoR+VNsdnN5ejxl2U1KCoPcN1XGc20FpPLLHFfryfEYPLgs86DyEAsE1FkUDHoIXhjSwQdrg5
o/AFy+JmdiIqlSqqTSz5CMfDf2cYDlvF7ajOIUL6EFzQY8mYjmAHXzA0mJ17sHiMR5zNNtAsWE/o
agb3oETGi8gIhlKgxmz7LcJ/YM8Rozp8z3L9J8n6Lr3qNK7YoLdtH1HRdYgXIA9oTLigJGn0A1GQ
5jqqVCxwborxFawDSPwPZL4lAUUSyWpRMz18TObdWzaMan3O8tozge+TDidJgRCbvbt6kdDX2GW9
Qwx0vHVP1oN+V4fmtqyRg0z6QzOfUI6S+O481GFI1joPVl+kJl1QWDZXusQuXMDLiT8ohrZjRkxB
YIZmP6DtsunQJplG4G/0wT5hBtDjUYP3OGAx8j+mx4GBtJpcnAxExgGBxN6PMM8/58HqUrMEs612
Ba7BOURlbNVg1I0kv9Z+mNxgHiO8FUzlECIj0RG1Nw5dWrgKPaLFegN/2Dksy77Tew+I97LeHqyW
fZU1qZ8CwHYdGtJoJOoZwkxHfyXmjh07qqyF3432rXO03tplLXWlNC7Qtm63AxR/+/BeUYQb93a1
qBOTylgRjBQmjnII4w3eNx/IoOxwQJXOaB4JY7y91P/TkUqoGnHATlmqfxBks9rjtEbqSEqh+zPB
Bw3hg8yaz+zjZOVKxPyTA5i02a89HSFFh+hB5CuPlCDvtHosYI5Og+gnEm/XAON/e9XrQvkS7fOm
u78elDyFsVlO0s3fetKsUXvJoLNDzZxuoT6KuVgR0jjJuMdkkIrlaZ0PM7oGnEOcajH0kZXNP5pv
jS313BiVQnb2292j2g5+vjI6kGxsF/nf3wXVNB3bht7MO+WEiQZxl28JIDSN93QHL2XT/aN4j1lI
A00pFOv8GOzLSRrMUnqBU04zZ3Hky7vAqAKkufI85Z3FVN7TeARgF0nPC3cmc7gBwZWOXySgaodu
vrU8Vvw52CK6G+cMisozIUrzbr827XvNS9/GM+vry/RcXa0m7Jus4+xPzHtgk1/Qv9zqzRtVsM6/
8JqIHGrAV3jyVVEN3sOclv9VCyKHuGgXTKRNvoEkErVw6AXajO7RB/Uwc7OpiZlEod7p3gG8dZZR
8Q/MtgOFxzAAw5y1NAoSUwe2qZ4s/Ii0fI3jYTdSHo2YFYpiJW/4sR/BU2cpnkE6R546eOjw44h2
Xu5jncOI/2EJRbAlZdE0dEoTGXpKyz74LvIDUXTige90piW0tJNMcNCgUlXm8MS5SacnM1WKJ8wo
8KwP71eZmABu04yfpe15+ARTKX9shfXL/K+hs0Ptax03rzFpSKHp88hUWXKI+/zz4cz9SiuP1Aeb
j/qO7wefCqMDO2IBl63iNhS74LQsGPmwDtxzXtVrM2dM6ZYxjssPsa6Xb4eGguUE2ipizd4MKG04
/xlzc/T9VCOx7X3TQ12O3fjOZB6bLnxmsZhQUE1xXlpMwju1yfDeHPtJXrnx27nq6l0wUOSDmuVV
IsAHe5pXheC90xPUms4JryCCXC0GLN/ayVdpA9WEa8MSHEcK/UV6pXE5RWfrgItgo46LbB3n9Qzy
rEV2I4OdNXo7JGGoZt6h34OeURtoxm+Wp7X1sFoixu7qTMVTUFKWbB6vHR715LRGOhz0jlG+NOnP
XYUhNAaaD9vbwt0WRCIeGHz98jsL195WftMW6WeE4qx1BQU1a4+gyBUPhHYNmMzETcY9Je4N862t
Y6E1/Doi8wfopZK1fjzqrs+LIOKwXB/icdkcAgb+6k842BCyaUVk9JnZEKfP3s30aS9yzPCS9s7k
OYh4GHZhKDac42RVZ+SeapNZ+9XKX7fPbBZpJ+Pi3/DM7uEK5HMkhdsTtuB7cb2/CrC2kIx4jd94
SAvLVXswEV6dOsEws+gyS8k4i6/TE3wBbiqOM1pMBCpZ0rTgX+g6Xhuss5cBvambKho+5mc8pfCr
OlIyplPHqwwpgkyib6JgntyzA4P4ihv9UG4REm7M3JbG9to3TyWUMDLT+ABsuitV/nhlztzua6AT
MTAcFQQmcPPM0r1xOaOg2ivH9v186PaC275b8SWTewoV836lFgWBxNVlJn5l0F1D9FyusUQgTVjb
RvexJswmKVfnQ2dIclY96ZRZYt7ZVBMoFpw/X4A2N1AODxu9DVJ/kiZvhW5d37mXRYOaLOhEuKON
zCi3FAR1qwpyo2tjZLu6H5QD7iQ+aoZL/d2RJyV504iD1eGSynoEC2TUxj+L1B/Spl88fvRC/T8m
ap/pufWCJRz3ZJsRIGY8nkBYKHFa26WVDL5Jdc0mA1HJClGIJFnKTMC87n4I6RuXrX9P0wdD9wkc
yXROnN6hR8Pi1rQU/0Yj7c5Zv3Qqz0+DijVj8BUva7rP/b4NnH+Rem/872nPDqGEDG0T/o/Cpgb4
CBinq3BaNsDDgRHl5V86ZGLtNU+OIdoGwb6xfkwiwV69FLw8FgLofG0HZk2/NmjFLyrj+9rXShi+
sz/Hv8M/5fm2S80O1NNCDI/bqL3fat7WCVeFFVHNnZKk6E8KELS/tldiy7yqghH2n3N9tyJJELhL
8AS/9eZA1FBGQtHRbfxIdAPye10dPwA027IQoKGyEMZx85bJpljq/ryQupblb8iQ4CDNWO7/W8Ay
4+i75Op2jGcO1x241UBEcobAB8PsEgb5kmSrjttcioAhzQ4P6soQomcpgELhtATKyl73INenbwMM
xo1nmzLC7xj4abckvXZwzBSLodRFhxPvrY6V11uzjgyWrVwTz+t/OyYi9NthimRTjFce5CKCDUc+
lM4f0hcGxovtrM51X62IRblcp+bVF9rilMU0bG7F7mu2wOLTEozyOsnCrZElLNEHzmZ+tA+lCFme
U79iVlQNKW5oewmdt98q9GyWRe/QktKBiyuoBpGq0Q49bNX7IDRzw45gX9k6pudHjYMROvZz+yeW
LimfG0ejxfbiYkHpinDrp2agM+dnkLUugIL+fXPI3mjzmNw6N2eokv6DzQSltoZF3Ubhwr5hE1kY
N8ocvWVFEA450tyWvJRj5r3XFyUbN3iajbLrMzWSxV+gj6TRJX9xSJzLa2DadQI0N1MlNM7IL4GX
n/Wu0LCoc8eAORUZ8gWWxciWAN7bIfEP8ah+r0aHm5Sqxh0Kot8TH7j+Zg7BMumhzn8lHwxtrll1
lTx+dAuG0COe3CrD2SXqYF4GIGAaijkHsniBC64DXO5rnDwFEcdf0tB2v0DityqocFmN4I9W0HXo
CZb/0kV6emJP3CmyoZ5qaKdYBSSJ7UUYn48CUPCQr/U2szPdUqkGv8+NgR3zRHGV7nhOMddP570j
5tnOmba0LF2A0IGwHtVxhHUycbxlM9j5gEmwa/2g6ijOajXQUP9RH4oSpwrXd0bujV40K8a7flf2
VJhVaSSnAAgSTUUHmQBsQpBwPDljhR1Xb5W00t7ANZGNEq5jF72mCCPO/DYLdRMtKz6FlL0zwlXl
q+R3DEH4bjqJltIYONWkXBodxF/ZrdVc/+45M40yPTB/GPeUgzvDkpoLTRflMsOvXlVhfRPv5MmT
a3GNID+7qw+2+OKxmEvsw8sdEv22sJuSCl+R9Rxao3b4BI/U2FFG5VPProCnGuq3HvhcLYRte1sT
gVxmIx/H09WX/JBNYiaZLH3/0dDKDDvpJym0g3ZloO/i65oZkStlDvyGnJF2diYx7opxL3/+tatB
dfEbBmvXtxAWV9pqdlUlwvUeDPCzeNe5IsZ0meS+aH7lVHByO0BS/GDmCn11l3WoKG0TYxjodVBD
qSxGLCLJmz7AuthNGbkdEa17GbVRDFwHCSHqgHO3sd08fe1rT57fQ0xljg8BKtNoDHUrjEHBc2I1
nOLwfB88Bpp3+OSZFQOeAJOQwIR6bHz9X8wbP3qFkBtxW6FAGoKIsvt2F8gqjhOXq28wP+JpxLao
ppue0zh9q8tULiYh/JPHqgtZ2sySUGEQ3oqQB6PwD7xyAc34JXD/+N5a56/Wieotb8L+OEIwth6E
uNT8SXkaDjta7UQyZ9j7dMNKv1HYtpbXIOZHYZwYTA47opR3EWzjqIH43LrIrmFkSs/v0lxRrFjS
UzRVlxACHVvQYa87DiDmO1tuEMZHIFrFYyFNkJiEu1JSYkyVPPeTiJeOYvDy0xBIWXyIKD8CbpfQ
354BDXoJPq80cMLCuEorRCLwrl5aFwbEdLul8GPSmi74wg8TV+dCKbECmPrGuHIh5StFg2nqX1F0
nR399S0fcBpgbCPmSkWtbbm+PkIgPWMijaw9uCk5NZKB08CuZzc0k8hvWJ6q5GibNNYxQuePjwpt
L+03D0Y278QJUtRG6yZKCSolsZPDOLyihXW86uiDjNOi3ptNRCbmbjkrqg20Xd5QCXtjOtUeo1M8
mrvRVgV/PUN55hYk+2w4U8L7CUTWKSW6kLmZu/N8/++/gbRTcQmDw10WohrviG3CgT6XMMfdoMV0
cqAtnfwj4//7BQrp0vzGW91VCxnhKcHCpdk4UTwCwsgKrvfDeQANHTiygu2mbbSudv61+Nc5Y4ki
7nJhptxbJTmAm8e2wVvGq27rre69UEFuNuPcpnXZpadcLSNnpMdolia2B8UWQOmwJWcy2s6PRTk4
cW73oxR3k6P68kIq8hwKt9LjBXHLMy90n7frQJb/qlMKb5ge8J3tz3kq7fatwpOdYCmftjBmRBCn
g+pZM3Rt5q0RRhF6pR3VdPCpBbKjUXgrWmWdABZm0fa3MyaZDr5LfdOvQDdSaH/kl2ZRTJRdObcb
HqWFZfc6d2+we2Vc1iAcq9kDL99tthHIHtzaKjc7tHMz6meL/NFLp5nthICJY0G8AYnD519mn8Ar
FSHsjrqlNpLaMf+VtWhLXomBdX1MFnuGEouLrSGPKWutbtV3kobP8ppF/E66YT4SYN1JgkofDOsm
5u+Q+8m4IVldE1StaWT6+UWtuvA+IPgmKqbuK5CfPGbC1XWfPJ7gFKZBjPa6f7a4GgNExES9Zjd3
SotOnkVMXDD0Uo8SSLIpI9ZpWiQGx/iEBjOXXyy2/Z4wTgXjO/bhqnJn5feXhzEfO4UrLie7C7h1
KA5+Qz15qPTAWqFZS8qNrwDRYp7L6N1dF7nHhAzT3qazom8Y5UqFeiVWmnI6uDRuQ0Pr8BKr/JaE
eS1NWtU6r4mrkR/OfouDp8ZhTsKjbuxG4kZ6m8mYNztmqo6a2j2thoWR2jCANduofj7gSW9TSFqa
XlCjam9PdIoqt+BD0hiRZhHAd/9u3gkBVijnQNNAkwkl4fuydWt7OwgOYLqw+kuOfhcCl/icsrvj
d7pzO9ZKPQuHC64ayDZPenTfBQBip1tYtIYZApTaLzLJXj/xeuq9Dgo9wHQ09pNCzk4nHAa3lvmF
qIscIVwZOOlbA4k7KGFW+zPMt4RPI5/kRzfeMNd3CCxcsPTSbf/g1JCCdt7jITQcQ9QbPdGKpuxk
Gu8rf78/vkDarx67nNAjK7z4p8IwDL/SYFknlgFszONpR/HzsQM6U51qIsOBPCkI/rUQwruRrmtC
FROb7B7CuwgocTOEs5RYmiiXFPj4k2k+J4g1j9ANACL8TT2EDyLEGtsGSbilpGP4bggfjnpoTybr
J3T9GWB8ikxdRkY7RGDtoz6vVMfrJ4JGcuzcnNqYh2PeCpikt/mKvGiZDbg6/nlwcoRdUtER62jn
VsNHDDZZQTBVz1bnDrdG8xOJYnvyzAh+Jr5/1ws6MtVqxbTq4c5apk2CU/haIWez6PRfykemKJkj
KfheCRE0+uoAWasGIttSdvlGCx05RmN3ZNqmJiaNSX1T+z+7I0wPGsc8i72caxaEGt5q99vQnLY4
lCxXP8ukA8+/3mdse0uFhoDLgg5kAnUGvhS+9GEo+E15jEvoYEgBYEiCT9YxucIsbmNHypWMCknF
kAmypQ5kFMVmIeBKYQnfAWJDT5B0k2T6Hn5IuDIVQiMr2eViXvRZtWCcRdiqPekVKCpgvYXptHAd
X3pelW86JM6OXNhIkkA6r0zCDZKPnrxWeyk4rpX2rHZIbm38dD4o8ibOwr+F+MenlxyYEnBVSqPR
UlNP06Y4VVaJ9IbcSUoexmF+h6E442iK3xs+kDj2G7WRLfnRkID4ApFnSEvFCwebajanwtk+atwP
VvQ/EaA6e8/gBzVGJzf4NnA0W2oPgNSH4ptrCyXv7YxkCQsdDiXQ6EoxRIz+knTtQkvLcTQ7S4kO
JdALPOrKHuUJTqybC8XU4ojSFmC+A7AJEgjnsR17Bw1+oZ4I2KQ28W9r6CP7tz6iqSozd5uO2v1N
wqw9fsoFmmVMM3CnOVqdfeUoqiLeZZ+mdhDXK9iLV4Y91PaaOaUjXL5OryCYdFPy25pU2o++Ir++
oW0kxd6lGabCsyOPF1yWMegV6j3aBWulo49rKZa5d/IfNkzKlsPZZR8wU4uPY+HrmQ+2m8nOATQo
t6A8CjuMy6nky10CZbt5wyf8Kw+qQo96Ctr50JryS+EvRqlbF+pvuQe7iHKEdzVt0v3j7J3dYay1
RNoQIXfVQcHruJfliU4VSJUAIbFqYLp38Bnpg5fxV6xiHHZKmJCQC4++BkeEEU30kY/4KFTEPBiP
PohwPLZwef1FF+/e/TBMVa65O7OvAv99wXhAAbgrwnteXi8jUQMfhQ15AYCqvzARnWBxaiL/Smja
G9rN8Rei+Q4VOG/pZX8mzVV5BqZRRVeDBGJPozBqXUHaLS8TTbe/2GjBftqTDMptmUO2H88MLVVd
re02VEZw6bsxD88ycO+Mf49cZqmXw41zTQR03b/xfB5R1vtNRJrafOWEOq3lNvkPVVx83X+LD7/r
YAuaaecRjS7PmQkh0N/WxoHkDCsvOFf7qy/a4AAOHLD41k9rG3dAzUFA5fG4adQ3DJ3Uw3kEgx9H
9U0Z8590xLNZZLz/L3cm67tf74B0JvE5RPf78l1ltpkM8auU+joKlIGud2CjKerGtUv0K7HuvGrs
KvrHX0GyoqSn+024ivO4Eefgii5DJlsnIRluw0zxZ9ceHs6pa3QxqcemFhalbY9B8Iv548XCTVZK
dasAFopc+p4kDX9Mj9TY9l4mquh6crUqfyzwqbsMo6Q5y7IRGHUHSE95yK4jBXyLezb55cNtX/pe
AzsD4o5F0UrFC2zX6TPABvJFz9SHi8wDZmXFNxKdiVORDkJi74cJ5aXgZ9F6xJZnPLqliSUz6Ohw
Phc33oR0085KFK2ivtwUfwEmKiLCtRbJp/XUpf8nhXcIXhRwV44XNipxNcI3qvbD3peeqOxlTeek
zCTq/zAZXeCmVrNARfZaSTcb+qEu9BaPL+sxneTGMm4TEyb1pTJlKhEuj5y2VY2kleRNpzSh3MzG
HVqp+yQ6DRzhhSZP9kClCcHrkOVzJ7/Q+RXwCtHN9xzK3PQ9cd2u6bN/YmGiPm7FYHf3GujmO2bW
gLJ37E9f3FraOZ2uMsR2vkn3vbbB1q6AA2z3mUVUaKXvgbM9JaiwoVdkf5xeL6fJy+3XieycdB3u
C/Fg7+bnP2BIeZ0dW/b/ufwy3o5DbF8U5AUujY0tuMvKrZqdkrpLm1NJmhXtYTExxDmV9S4X+N5W
i4ai7CjfEOcAeW1dYHLWea/PX3yNRdlZxxsd9sYL13OyF8zX8huaEhjAEfGbmttTMqQM2j71DbXr
NBjEsIwCLutwWdDCXORVG+3Zn3MEOwTyqwZL935B5JdKXpdMZY2LfTAo1qTJIaQPthLcuawmA8M4
6tme0RfmH0vk+Zp41f8Dh0X2XdCdE1zn02MPKa7cwCo99G/Nmu/VH66xWvX4DdOklell2/8I08Te
ES7jXmF37kSyWCNDwQ2kpnbP8uDnCSGuLMXvcFrP8TZqJso8jEkKJs/BTPZRVL6zLl/5LkrZjM39
Bq5UGd6qufE/Uq3J4Z3Ok8/zxdvggKbIJflRTMvdc7teS1k8jhe+9DE+L5ML3QKyyJgG5yCiOep5
ExB+Cr8bkWaFtnT4jeuwKL7B66fnLeyYGCVfIiBu39Upht5mGJ0dgL6sPFqIrMs15+RAn9VUhbVm
uFxXXGsnflAj1dcr83fQ2jAOtNmhWlmHyGi9iiHIKDI51h73JjewW6mh8CVFeOFraPw6fKVD/lD5
M+QAM3XTKnyoStqiY4mUb2hUrdnMpu/kZljS3E7pZbAJXt6fqLTpYOrVSxBHDzm1QmrMYWjI1eZW
HihWkxKCf51x+58hgeUlB3Lw2S0hKU5s9WAbZNqOaBib0LnT+Hz6BmzlBTLWa3nJo71qg2DJSGaG
lqFrV+7lfU1d3Q2TVPgPl6zuu5TC1c8h5VR9xMR+1PxipiskEFdbyu3R0IPTKzJ8/IOe7ONE+LoP
gzuz2AgaRWDLjZuluE3/OxCEGlZ8ibjSqUH1g2KHYaN4JA0hwAf5HlxC263q94XnUw7L324bLYiH
pHwaF9wy0Kw2qFxg2If6pvk8La2wobDNrekriZaLWBIEOJijSpSa4iJnUTKZZJeOCF8XioMx8sla
qe/chVDxrddQI+IcnDvey0hUaiPbGoFzE00wGxefp+Ky09dzvVDw2tCKHty/alEFH+U3PUWOUdE9
6L00WHBVgNr7RuOCHJhkao1h/qAxYxkdx/rgrq7mD5+W34xWdIB5QVFgM+DEvCdQbBF2vT/7VXjx
uyjBsmsUwkklnhr8BR8zGvc03C4ZKrBemqFfE4PRm138RWuqdb2el4vu5OolqQceD56md5TiXbsn
MhY0NADk3AJYg8j8ZWvnzQ3ml49c1SDc3pu2gnu1q6Sv+g6DoyUDWHEJpd5j7xaQyv0Wgrr7OnXr
PsX4kU0irVshfHMzZAcQp68z5N6nVIdsvnshrN9Wvl7jWYls7OJI8sADukdW3RPDTkbrN7oA9TfD
WILlZRBLfmGOe//z5L4LRDt/+/SvxJ5Y/7rN30Z+SBOGK1Tl/pnxpIIu6pHCkpx3aw/WDOWTqi9S
bdmababzJUgKYz8eGwYM49flK4+StPTHWctDcwrNho2PshVmKSvjoycSIjpaSJA4vgJ+8fKoS3Vs
9mrDPviBXA+EUnt4eaiZn0NhFviZLlCIc24an7fIbM6ZqMUtqpYG89aaw0sFId/pwAXO3rFjG4Jo
cr9e/SuielCouDpjP7i9LMpZXQgn9SPYcnt5dCPKBeuAzwNhG89sUDL4nug59ypJo5vUbk5NOctO
rE8aWRLOgqWZij2D4edzYQgHuhEEOXwvm/Xu30SdMbJEloFI/yeDPnH74eBZx5M1lEoFkk3Aosjd
y43j3k26KcFBfwLrNQpaKUkx28o0RJWcUv/n8+3Hz+o2f+Ugjx7z1I6S8MwXPqKGbHnpZIKgfjS3
12Ui9+69xRk50rh1GjfkJEIq+O5FZt+Yy6iW+bXG0azeQfe/tDvudSVuEfnpE4yp+2OLViSGiEsB
rz/AEiHvv38wXGOd5wCJEui1Z/opD4MBs7TqVwfmZ1bm6KJPob6HEBRIcGBGKOlujd+eu8mMum+E
tJCfCVHDkaQ7jOzCzjcqAXeOKQOtZhnQF74nUHczpfmZvIQVAQoeBPdX835nhwJ74N8AzYdM9bDp
/ppvjEihja1lXaj/s8aOsbMklQ9MQE8v3SnGKybwi09fdloFX3POi4aLIPdhIrcFZob8LO9ogtye
auWN5zR37zCMqvvkvSXGCU/fA0bymGUaOKMUqHbDJPBeMkNdHZS/cX7QBPpqlzl4AptjxPLAHj+p
Mj+gk5WIUSONfoIR4X5oYF8ZFxwsD91GlSURMuq6M6+fTZzAGZqeB3umvvQW0wGYOEiPLPAD776h
fjPONTNXD9w09SzdSVKm474XKUwL0fez6V7x1ef/rrvb2PK6Z92x0Jtx4yVDcu+xS1jgcDZ6cswE
0PmmIk4Z87xFdRFGDUx1arQHjOilftEpv2gTSprf3OR6oxmMqeXbd573VYQGlo2THBZGYRBJ4Fpd
8aEoozOMEdIZzr1YuAERcb1lp0q9Q/0NxfDuJvsFfFzKppYE4CUvQjqwBu+0dW4VwKhAVXMCFjAz
KxYFlm8x98HNTFcAg35Ocoauz30Om4hSLbbPdKn323qiOGrfT+DrdUerOT4X9rvTM0Jp7c7jkgYK
IcaglepP0LKEy1hxhC0ZxY89KmnrcPCpuip0h7zEhsTIEbOLDC1TV4lM6aBczI2fF6itcSg1lo3S
ejJ7eBa+zhpQtDJs5Gh3PWZhIfXSh0H8R2tbUuTLSHL/6tdLB9EjpIX6H+aINSMQgfdU0PmRzFTU
2Bs18OWHE8l1Uqz8csplCD5ibwbiMAAJyH2TBy+aWb5OtwQ0Aj0pfucLpx68dic/B83iSblRbqQx
mIpAvlTZmwtbvsOmaOS2JCDnV1eFiqy99Q86YLvSssdr2IKXVaeQZ8NhmbzKqNVuibp7rMh9HQ42
i5L5U9dVCuehKPYRmfqVmgcPmvat652NmAA5sA2/iIjUwQCSf5q9cuJn2VoXkVGZxswigbK2T1Hn
Cqbeevlqns0icXUSwrWAxKvsfqS4ZBKOG6KlAJtyNWQrpns2qFqfiUdGdbl7kXnR4vESeN+jMAsq
UvQ38fcmi14eWaXq0Tn3DwC/Rien+tZvyip5qvFxgjNHC5cw8DOmU2LbTun/1RXan2L8f7PEHUJz
oGi7crnW5HQYab6jXBSBD/B1v0s1OQdcj22sSe+S5rwxaqoYVXfWeLp8Wha4gPQdwrMCplWN5TLr
CYloy77YYdvUDENk3IeCHzJk2+wVVQWc5/e+jpr7cuV1FYZd8CMmqXcpqQre6s+99094bkKdu/jv
uBK63MAvlIVxwsVGMMeSb+YftTUbO+xzyq5BnlXnNPaQJWiVO/E2mFn6K8xATJEgk607YvqmmTSy
RcEYpPcDs/hxaGNwMl9SH9qJ4kPpPJfvgnl0txgTSLDsxXb+bF9iV4KjFQ3KGri62gkYAIUakXLy
F8zLyZRFojIgDbOnN9S2ZsD0P6VzTPyWSJ3VHR/t7qU/7pd/wzWXGN9nKCUp5lCodvchokf/dk6F
VQ7g+8hrCBJrC2tdz8t354EPPPSxLRN9GGg+XTGu8tQO2Ltxo8dJijVVsgzWLnbYywxgq5vIBNGa
H00mmMNAWwN1WkmeOi4WnB3daZ/Vts9I7MIB2dqUymQ07u/Jo2qnooGEmQFxwRxQlgKjp2cWGhFp
S3/h1wfdbkdpVVgMlUMl7goqvSHdnJFbezgRl4eToEgk2ywc47/K8udnGu4RODYSVXOieFYVCbDB
VNehRC9Irw+waRr2moT4QMn6En0PVswqIFejsxBuOWOKt2+ZUilc3tg9N/YXnQVPCdCShCiHQwoA
DNZO4b9U4XJeVUH95XvpsSo6/4amwTpE76kSsDgKETWL+lGVfcw1ypn1wuRQ7+shw8hREhiTYuhd
J79OBLvo4/d+34ynMlH5VekWMSNHpHOvhvsmUs3HxMyqb/ygnWF/JR7aAya/s2gViT762DSJtsHP
c7Hq1k1k1BpaLHj9sf0dnuLJWJAT3opJytoKcGAKoDfLbPBZny43zlPjzb+6OCC//CT9+B23f4gI
k/pAlRYDMhyFVymE1n9Wdw1n5PjQtCdZCEBOdJBMQWM2WXOcaczJWIiWrAwPTwDjmYMtHnNKHpnA
dfAQHC19wV9BnJhMchu20GR9ON7B4b80DLbdKYZVuhTzm/d6iGanngOkHSqhICJG8IZpKG6G8nZ2
pO0ZhZjStAk0cbJ6moYA5BkdmYvEn9fF5TgUhCUxhWW9pTL3XOG4AIo8+Y5yg4E9NKrcc2ihQkiu
P1z+cpAIw0nhFRaQPD1uZi1AiYz6BvZy9uLCb4AvdHlfryJ9aYOQwLibOdZQ2uV4udUNYluaYRKk
+YOs5aRE+n28gBh37GswlOBn3PG06RwUTRwCE5VulHT/MPwb02W8PRoQVfa0WQar6o94VjACa1L3
ZIqI6hYXOlHiaGdua//NblZrdRWe64tk9C6Resj1D5rl4tyFck52Fa/PugZy2+LCNeVekPMgktT0
0GuifSvguru0qDSCCKayrrTIgTQcB6fFhj2I1p+Wjvgisr46oIexFfJzqejCPRbG5P9EwVk4v588
n9eVCXd48k3Q32Mp8rVOHX5eiKfY2wGpKFHyFCmMThIzpjB6t8vNVTTJ/i2PN9QEGmpDjzKI+GBm
eGrAk6mRyK4fAmG52bM/2RzCEGKVFon1VI5Q1EtFY4+NZjHcnAzUqXM9qDd80BMrpBetQikou4hR
++MWXZkuR1MPLcAcLbCiVpvXNT0fV9r9DcvEHrcP6bof+VJtv1zOZEes0Dz0x6O+3WFqW0YmPAr3
oS3Ww7PncxVzWH7YUHniSM7dA5uh0elD2fUQ75oydjiXd7LPUVv968p3NrZAT0i/WTxa1l0vtQmE
wgig6BWcGVpMGEk9qqxSY2SZMVRm08N1/VwaE6QisBtNDG9nmJ0K07VKVFarjooPXozn++/MqbFE
j1wqmhFBbGu96J09wmxUSTLMWsu8GAuNJHYNxP1/9pP6Lo/E/v6be9ioYlo3wWczkNteVrGnhuDL
6M5mBJTP+FhAAerq2QdXVuUpZGRtHa/fruCKE7DHdwCpiClH3hsYckqjSavnYRvcIs3XqqIf7KsB
kxJMxyaD2a7MEB9VBwRAzfRx88Uyr0q6hZfGVC3PZObGH8nDNxK3R4/nVqMCcXklcOzyfaaqacwH
Bw5L0hUmMHouGV+AW2Au7iKDBdTWWidcknBwR4307DMo2vMKO3+YwzVORnDRQBHP+qjRk+NN86Sz
XPeRVJdMTQ/aDS4C1QtURNcLK2CEEFAG55NVBHfYfI2o0jtSIZoevS4A4BGNRCOTEcPLnZo4M9Y9
A4LkUXKCc73psf0Q5QTT4Zabc4c8KES0xsuJUh6dKT3SIiABHxtHsxRe9ll3vj3q1D6pv8q+bIZx
/fYyKGWMP1O1hdkGBfhlXYkhJDh/PZaD3QEkqVh+XxVrRjMEeWcZlUOh+mFsmvW+JQrr1RNFFORa
isggDCh+WAudmDf55Fg4p40gI++zGYLAgTW7fEU+gwCretCMR3nUFWCIrn+KQEE954h8ofSKguUl
9v7D3TRL2dh+VSZd1Cz7GkWecWQJTEuvjNf5iUlsizIvZtLpHGAMxWffyofk38rr2KsaY9JSOUf+
kLHPFNsnnJw3f7KNrj5yve838pbdZpx7vyqolCbr9Y1sVa5jqOXK4GJhawfuPrnMMpo2+4JlDaI0
nk6A2RAHM3C9ww+6sc0Q+hlshowa24dquYeH76A4e6hayjLGSoo6gjeOyfqoqeCF/BNcuh23jdi4
U+CwKJAElxrGqbfuGqPF2Kn0zXHc33gs44bs5/uxPlFHN1MaqBt3YRyMGpnLnjoXT34heMA+VK/d
bcOdjdaVcmx6vvPAGEtXgpK7J92Qq//jKRi33kvwBeknH+9q1ZvVM/dUvAeU9TmumjZa5Q3VFbQC
RzL/DxVMv4zZh/upO4g+VG6Y6JBWdyZqB96j3/1RYij29aoAciMh891KuLz7YV1XMsD6IrfQYLAO
GfU1vGzh0Fz+d/KT9iXJ5tMiKJ9LbvQI4OPzOUftAYIbPDk8fHJSPdBvjxuhuIomBMdx8zSakrHb
/X1kKEeCM5CFcZ4uW1/Uy6PobnO2R+tzgMdegNrqj7Rb15RMiqCVneGThxIYCNXiQKqvkbKyn9Uh
uOFnJ8ydSGIIb8Gs30ZwyQmEAP+41tYTp9Q0ZFCl5cOWtVW0pEL/wWwJPQuXfbvBBftyZa8rjAmB
Tsf9BIA46xbIxasr4uRQ/TBhi4PA7yA3ytd/FxohEVUc6zCJddagjNw0NunZpCU9s/x1fuAp2HDe
BNx42M0/5yP6UupFZCW0bH6n15Nx11I9uYAw5cbcrZx1opkMmYJfq4hn5V1Dc2NowqULX7023B/n
ClfkJl0ZFSipscuazPxJkg9o42EzmVeAjXfNo21XopWINel1aLncBKazhHLARzn7AnIBGe6iX85Y
cDShU8oy30jJQ7bVYl6CUUQ4LtBN5TlVoTOMa2A5omW3KX4K/lVr4vKrZo7AZVksrwtP9IZrFQ32
f52BIEFS7tbLjJ5dX9b4AgwHJTaEtECgTKl4Q7KrA0P+q1HyDGeuVuUryDSejlN5WEHc8vSh0V3K
vzXdTyPJgd+DpndWao3A2OaLOZh3jgTwm6vs9coSojaqnYRBel5JsfZPRFMLLCwAYkC262MPZKRd
fZPNpn6pUOOiBWHUO6EDMfmGNvxDRQEqphDnKM90GEFNUFfHFTlW/UN0UtXM3z5sfBxDZAqyxZgU
ydrcwEBiLPYpKUy6O1/cPtZiwz9je1mJ9cXeMwpctnoksYgbZb6qhqJduYmWzL8EZpIiVlLyGlgw
BENq7U1vShnmzqqqFRLK/Wbh+Kcmx9mJAUIXJL3BCPA6gtY2zVcBAANR/S4rwou9WpxSx1dZF8eI
nDCQ7eHKcZRjtzkYwDOXJc4DXe7XeaPoAN6933eOsVRkZl7u2vZe0k/T4GXTUL3pzK446S6Try6k
CLTNF4Su8pEK2dxu7b9SasYIhh0H07zp5LXNEghKUUEQbwK4aP0aQ1/fT5vtetv3PpCqZdQ7lktE
Yij+Sr0VaJqdfx/WsKUs6ut+4tLxiG/Z4AE5g0bXcPkArBQxRMAV2rK0YAI3waXHV/7Y1d3UQh5r
NoFZUH5XyV2ZOCjcScMKOky5o1ufPIF500sJh9tErlDg3Suz75/O1Q/JWK7+SM0J8ILrwlf6JBjk
9IEqqFQ6oS+obkd7WFuo50LMcPQazptPOwywlNxkuKL221FC4Bm3rEa2fMXxAytHLTSW55MzebIz
zOYhf/ukrvGrzJecV30MyoL+hBdirnWZLUgiKu3pJpK/9gzzEaNrQeDk4Kk6Bt9VBNJa2fo29nR4
c+jSmSml3T7ZsATcj18PaV1w/f0EsEvbcbyFy25H3XOusXgtZxVCPs+7PFnYxNxVcxoAWqVhKa3z
MOFQrkgPkTo1jtGkba3qOHakyCq3jSyhrTDB9F/oEL2Z1mE/FUn7mqj8M3N0e0r4hgt8VS5Ms0bW
2AwEICfsaXnTQ1lFojCB4LyDrb4t+3Jddl9zsL4TlbUxNyur4+GLm3/DFJd6d6u+dQFf28U+ZjWg
zywou17/PvSfs3S8ZaIMUV+9q4KFH8CitToQbsqk4Kd2Ohb2fML1biQwYR/q6xkrDJ1yZOgmWt/x
WPxFicgZpDH9Ascy8Zb9AHmPdPlQ4k1J5rXBcJeMu+awCPun0mLpN9m7Rfd0X8VWUTroYpUKI52k
unCpwxa8St36gpalEuAal6vnmUK217sebfFuQxtlzZYgv1EZluJNDB40CMRzBG+6fwDeHPPQkMWp
msV1Xfu0X7z0ccp3YOnrbfO1eNCsl7NIthh6oapDZP0XAA7A6RcmQuFLUQN10hwcaGWjMiIj44GP
vFM69jG4KcBKNDBVIAgbFKRw8fxRo5/BvNgte/SgZIknJO1s2MoYZu7Hcjd6KXPpCJiEzTEn/0qe
cSU7SG6JVtlC6U5CpCoznnlWqbnQEf0mGDKiAKYZZkIp78oezrLpmyW2QbyzCNPmTqPNNvfaAsOk
ysjbmZdUv20c1WVG9Tj1HRKYq8SRo4F8SPxMYiiaGeZ/WMES1obRsUpF2jhyUEXE4UBu3MLJI3c3
4dJ1by3PFxw0qG9I1nFAcuo/cd7agszfaiVe0ypWVKg1qgw5jb7SOOndq6cAdh74P6rCYq0mDUYp
x4bJpvYAv9b0iOdjQvF03loF1i/Ca5VA9T7J+hYvL6PCpxdo/853R4OTghvVyBdzgUim+pc7+eHK
y8sjeUq/6HNy+74yXI/d3aDzYJXqRUe68uAuPqvEbjMRou6/RfdvKcGVCTvWHImL4UQVJvkCyg1j
08bFzuxD0bJ1/2OOYX14SpNegvni8nZ1M8N0A31fH52LaMJm8tohVL2pHJQ78qy1B/kazLK14ppd
ozR1W+KTKG7ienVYbFncPOCmZeblFdsDJoeOahvJYaV639o7I81c7zDF9VQ8am2LatJ1Kpl+AzpF
QV6iPTRdgW4RVs1gijMRtgb+yWdusNVdB+/TNV5Zom7GOl+m7V2SdSO1FyOC+onNJ7tXLOTDWGKw
xkKTVIp7Wl02hZZGkIZfkFYAdj0+9r5jn6EeWF/0B6dhkINCKFuS4ho0M5ZlUtKMj7S65ITzs7to
XcZe9m7u59bYuTJ7fr+PZUpc5PgubMw7icn3COzltCp8fImna2YYw6vcjsx1OFkmmX3s3tIsixjX
5RjlZLvQ/zXQkMsAPQWUoZ+zHD/hVYjelh+zUqLmEbd3Ic4UVZX5J59tkA63SunC7TQ1rQ954HrJ
o7QW6DebhEC00/ysm9FS8K6GZ1Btoz9G6of8N9sCbMRb2WgaDKT4bP8Mw3pn7k3+G+EKnW3T56Jn
DsWr2njKXopHFwAxmQEwo1FO2o1zKgP3HxRj5O5Ijr+pQBMZmBy5m6lpbEKiiaWvyQm61i0NZEXQ
1IvsLSVFccA/em6zXRbbaYgjHTJKZeZL6OBDWX68T9WJZ9dejbSwcdM6fjc8RPu+BT9z42/VKlxz
1JyLXvmcyyC0CRjzhIzvccONpUYry9VJzgg76ybbXJxchhWpTmfW6GUUWN0PH8hf4JtvxPz+d41A
klXMlZicMLPNhL1u4AMRrAWuXaOCjJLb7gIf/M+truu7EVlZ23WWcsak2uaxiGW8JSg+CpRkDlXl
/NXw3dqjHovE/WoFiWGYrWuZWDLyfzzIXviKPecz8TiVnSHcOUf1BGvX81phcMP4AuGtT9loLvwm
itkqvwShcrBEah9DlTTQLGxdL9/z+ZJw+AhskwRMSLUHWJuGWdtXn/Vj4WQiptC8S5bBtWl7ax6+
13SqjUAVoea0J53S8ToMYx9CV6EGI9Hmnybc1yJpOmxZZI/TMtNAE89umNc82XQG2Qb9uM56pZV4
Dxm6Dk823j5cAe08zr0UBnGtntd2GZTXMLLjxcvkNeP4fGb9yXj5l93wiWcduEm0SmrIBZx8rZpS
PIyb4jrmf20G4x9HT32MWOvSiOArZCXgj4Aey9+sBUZ53iLXeb7VhMQgpQSt0Ul05bpr2pM6moWQ
fOIFs0LNtivbFsOkhSVCjMYGReDzBgZyTOrQ/uxowmX1Rbtu5G42GrodR1mngrZxYFVhN3yggJgx
6aLTIvRI7Ay9LJtiG7kM3BQpTilBE9l/gX9hDejJXPg4NNLSGjtKI5d+SVMkUY4YccjH9bwO1UvG
t0UFUXGjxTLSECj6bfRDkL+Q99/ASBO9EBaUcQ5NFBuo1Z70GeDpKp4bBPoLH5wlVEKns+H1Qe4n
MIQTkttbE8w8qkmFxpqAknThzZcD01qUzBu4Mfzm/H1649dYUdV8Z0VG9fJjn7OkyP8EtTN/eVRk
zCDPtiADzD7YuIAtfHzJ7d64hphR/xu/2CZP6poeKItcnxgSfB7SMSJ1is2Twc0Bq4FO7v2IiCPT
98ihBuZhW94Ti4iUHSifPzZCUqeWDLCzeJb7rhrr06tKN6UBhjtBKcZ+CAv+kdaQpmgf6PFCGRrK
GV//A+lhxfWqyZX5bBMRozW9GHb3KRI+jjKtUCDIigYUp7BXfRVtZX4Z4kTMPOcoR/JqGDxaGmtl
D1gbi8YY3ZeU2fuYEoGoPvhXMoSaleT1BJRobLHTpiYg4cyAOZXcAKtDm80gIpdaq7xW9yMb2EEe
Tfawt3OArEMmotfAMYQsDffRxQuWhgtTKVW7kMkAowlh96jXwW+4EzD6yx8Dn84VeBjOMD8fBIDE
kkvGO0gbpZCyRMmsL0dureuGL/jx/cnNs4hcZWq2G068B62B+jTKmqApmKNDaQUvylrAh5NsmY6m
3dPvvQbNSmksc66XJYTkiMDeNeVR0qpUAZF/cGRlMaa/5h9JgO6s/ObToUksR1AUO6j9+MuU3k1r
Mk4b7U50hMgTNPSAoxhUDKtaONcRdXzDFJ0MwWpNOm6fyGG+nmK2r8z4KswOpzqxbPoFQnpqSYTX
fPO5snQwiuv2jCetH9iZOSwVy7BZkp9LfSwCFS3w6Y8fPLV2+vLMA2o7LYI4XW0+UthrSs2OTu4y
z0kNRcheAhSg8ycLRJuVkJN+aCGuu+gV9rDsQmDDqbnErtM9AAcP0pLpBNZDJSvcrbqszEXZSfq2
q7VNVRzy8h2WABgCdfQ66iAWDf26TZ8grjUtTewTUcwczvZnvH6NYf9zr6Y18t3bl4mjbt7DQggd
WhJO0G4wEEofUADpTfLAMlZ4oySka3JPBiEDzxfe3FBwaM3Ti7zl0+m8UpQ7QsjXT+y3VPUG6i8P
cpeR33/p4peznMhMh50s+mEEKa4dpeFIncti5kFVvh/32LrJ50f1h8l/kj3EriG6DQ6GspxQLlv6
Ih8CgnU9FMtVo7pg0QGft2pBRpmQJgCijPtnZFY1iEduaGEwCjKLod3X7YmJdH5PvgmJ4KRE2Mqn
xcpYt3BaXI64c3wM2gIbzzPo5FqmDtvMJnEw18c4I8atELFLqIPjt6kk777ypnR8PruNOHCyjIYP
dmsLLs5DoJTqrwTKOyNHwTw/BWPpPlHmI4EIWIf1OCfjSCMiSNYU0eKu4beYz7em5l4H8z7RZ0nX
r28eDUGETHBPMhfiC7cBhJ2x862I4FiZuuv5dJdiscaSEtKOMxVrfl9utR9JX9pFWVUTsuI8rtqw
YgODDL5hRHeJNJv1UvMk3PdCpT3qPK4wnXywirD6EKI7PA8e0Z38WEcqjHv5k3bRtrJInNPWXPmX
CbKB3u0hzgf/a/H4UQtdi5WYhaBB2kqEpsGjkhc14BdYmDl4sXzljYerY/F+Ty6sCEAfhyIfeWKr
CWw7Fy3x1YK1tb31HxcKT8WL7Pj7cdCCHurJZY8tizfP8Sc0X/hJJSkE7JmMC3PLS6H8SWMzJCjS
Jy0lMEGYrf63PAMGKPM4T2FImPh3ZFnnKcE8IBrL43RpFuzNx6pFmQuIbS/Tpi6mbg2qnA32JX4Q
xOLc7dvIuTSQ3FzorTI0e/iOv+jshnfrYqCIWsQbrYfp43DNkZtbipnKRDdwVwygdX5mIH8iS5IB
MnjLUZcda4cfwuvv/IARCH2BjWI6O+/JRXmfysGmbVSmBlU3h5XsixWRaM6K2YkvBwhgHpPtpU0p
W9dqr9vmGKs3GXsbrfCY8jtGYDU4l/5+ueluckOEDc2rco23xODOOHqBUxM69DKuDQjkQBETSe+c
P2ZtJNOeUZE6pYD7gXyF9QOafV2M0OrceTOoB273plEwsJ9wHCR9NFWphuMqYcpdik3qvsnJC70N
5H1pd4Wf4owH32ezrhvObtqXIRfO4EUr5DMlphR+UmqLdjD9Fj/eEDBk41W8MLl8hQK3Jr64zyfS
7Dt544eg+GHV14v12hByVvQeOiNDLgD7X6026tBtX5IFOALz6XPcI231hrZ61DIpI5thY69lTzJ7
YXIxPnhXMNoQiUSF/ul2eTBNVScfPPxeskGnJiowcGtkdqg3LLbn28nW4Tu7DhzIJfHvA17L8Yms
C625dlNzxLg+SEr0lX/+nvzRW87zBfAFuC+x7cP8MiXFLSannyOTswyBlqEoO6vo5kG/jsrO4fjf
v+4Py9EJ75SxwZXm7PF1JVkltSzMBLChIAMJwl54MMUP1oPpUza207L4XHpEqNQnEoWy2Tode2Dm
Qb+Bg2ltICPjSQE9ZB7snF8D6xY9cQRL4ClYSIjOQyjOKuCq6IUwHba7CaMp2C6JUiXzHKfM4OgZ
mG8CkrfYiQb4acYF5vbBgdGVhUIYwp3TjGbO0+nWTt3+HPrZkEDWr/S2PQlVy1b/9+/X366mhDHn
d/gmP4oHZy0Is0JRBzzyEguXRXdhZ2h/Y7xktzGa+vhfszFm603Yk+Exq2ZhNYZzMx1mz884/zNZ
H0BL9pnmaYaz/0YjN4O5C+9J6MCmqrULS/U3jDYsQvKQOtVjd1FZ7M1C+81tr5iD+Nk1cOE+i75b
OlYl0TmigYTYLB5+pa3MsQnryfK7WMh08xSqCKotAeMkCwiypTBYG6he7lmTi/xv2HLyOpAySFsz
+2KLcLjphaCHAdWU/Kmk3jWTbZBz4AeAGP7khHu5VS0UZjzcl9CPP9KZ8+sTW0QA+4Yjb33NoY+2
o70yGL7JotOuE8Hbyogmu1S4EeehkJZlDqtnBw5WYRQ6YGMqAVFZJUkKZobZAvIsElUVZw55MQq5
n0zn74CDyaewNBy+YUFKp+YtfIfHE1amFiWJ/3ugdqEZwroy85A77g2ywxGqNO+M7kF4jozcB1Gx
ZRg/HXMMQTE1FNmUo9C8HAblvpXtUroKi2yn2eOsf909fcnhQvuUzl6lBe1Nsnfb0mBsOgPrg9H/
toMSeif61YbekNVHKYZrkzln1fD9lTRMeStqXjKNdJ422RxHUmusC2CfwOUY++Lcl8PyUYs5U8ZW
WEApBoJ8guzroSN7jQa0UYtawXX+MElRnYxhtRn//XTUW3xV+YKAIjUdxdcghmFVfdFOpBHkLl3Z
zo/4qQJ4Q7HtdYJ3Rk32Sei4C/c6oXWxFB46xKbZwhuBw/J/Gbu7Bx+Hw5h35nkEoHXGxhxHANfe
wm/XTuPpq23MCuf36dmByo3VZwBJf9FCgi2CxubDisCSq7Wvftpk6WfehzhkscsSYmoPT6IcgYep
1G77tcGQnwS0eJDCQ737YQjCDIy8PjJbcJORaxFzTpXLSlV7wYI2ulmc9mqCLt+/IezZXXfVo2gu
EeD14yQ7kmeffWSb7vaPnjZm0uZoEAu2f6UioPXI5GBOWCfqoLOhhY0Up67O49dJzheWmTB67761
3RLtiaPTSw1HDqtbgpKmTWz2VmL/CPXuGc/JkIuryPozhDwGElPxTnrDniRU9DTpmtyy0ckEYeyo
8oowvYQ143hW/lrJP8tyWZRWsTVvsk/Q/6HW10VXlIazOFpK3Umn9oSWuc8pwK4ZosGOzGW+bE4/
HET0BVSEOaVMuXQ2X8CT6BKfVTZ2fSTbac6BSR5/kIGR8iCnZaj7twFH27CH2fzoSneGf+hJE9v7
vWDV/VtB/WF4JwxPGJMREXEgAYot+bbn6sDv7RITeneywbCBKc+petJ66ZHtYvHqT/vs4ObKd1Ki
8/Bly/T75JJoo2WupQ4Ul2dpaKqBglLB0zRk3yhdCX5qxmkqXpgIlJbgEm9q8exgeRuM1QDO/Waq
ySDwjrDEsmBJLRBUcMKndZOVJzCMG4Hu7RzWuG4+Racl4NHCyY7YdozDS30hsS0D0Cei7fV/wLjf
USHtqucaSm2FJZcS7oz//PcXGme17812OwfjuT/FEy1yCINZaqTWKEu81ab3poaLmgchEnvjx/8q
CZ/FPhz9FTvJXjNHb+lo59AYXaiem5+KgFYDMDSBkvPMt7DgrEkm16gYbpKyRObaDS91dV07NX1k
wmPODA9mjgpnQ7ytqUQ2Isg4mcT0NIZhlfDYGKjA+awLzWjQJGYwO7EzAe2n/y/0Lfc0M1F1vK6K
I23kHcozysKSS5amhQwFLybUHJ7gTuL6EyuPnWPAnO6su+UfwBqFk80A19Q1L5Jw0q9uZVIVG6Hj
dhS5/PSEX9WvI4M7i0GIVXO88Sb5B/+ZziRb6EpYuOGEMw4Bpmw03C62atoDXrnbV6yAdZxCgts3
pmfjjkg1nFHQxKP9LY0Z2J5vdTP6N6MLyQqNV522BuXQMPge+K7RomlAJUQCWv+pK+nGHifHWxUD
Ag/VzYYQoBdL68IrH1seWgK1B/Ni0ihh/pf+bVhK6I46Ikl/IwQqZd29OfxlBe14MDCCmQ3y4Gxr
xKRBpawE3pVubrJUF5bDfTaMeS0xo8jHrThoqQ+kvPT1Zz8f+m/K3u442FQJEqoVP/xkN3MSnPQS
RN6HaalWTlpn9GbrEuHQoD70fVAZzCXZeGpwZYVEPfvRuAeed/rZdmi6qSYU/IpvI8CZJISB6hPd
sJ0fZd5bLSBpgOeEGxhqooxCBWwXs1Keu3IZv1abUHe2X4sM8EYYm1dZOySF4IlMhKSTsdnKSzea
w5Fe7+IGH826klKpVErR2BWJamL25tt6LUGm1Dv4Rw7GqUMk41ioU/0XsMoVNaiBsTKPtCEGuRmM
oTOtk7sEiHHaSn9SmSuc77trfaQ1W0cGO/NVPCVMVRkOSIBbnUVLB2DttIfbtUy+qoHPIjg1Nu0W
jo1Wf7RMUun8vUJnqkLMfQc3e761g6o0AsYK2dO/KgQ147RJ1RAvVkxTEZ8kSWKAkGftksPCTncp
YZPV+hxgnAFkY2nHjdBJA/dwCRyNbcgPMPyiVzDLyg0IYIBX5SwtIISc2DjIvtoOa5R0Ag6LUkrt
sDBv2Giu/077WzDeD32nOwphf4UXWaHHB8JCow+FbCAo9aqcab4fG+FQfh3ZqX/KQiwaXkxgSCvU
sI6I43uwCagUBJy7FrET4nAAiJYiLm0ThuNzC+oLNqmn/ZIPF3CiXTEvQRGjpjtF74m3nT+Hr8FR
pd23IUQds/MzdePEeQJ59VRANmRbQZZJVPdi+C3OzEOEkomxSqeZ+F4UcVEFcyN+ItFl7nolZ3X4
rav2QvK1vEwni+hhSf+2GKhJyh3mVRN2nCKfs0dMNhQpmweibOW92jpaNf2Jxw5GAwiLJZrtpSMT
JETEnktR497+GAOrOvoOWoq8TAMUPIkp0gqXR9FBSRDrUpV+j//VTCSieVID7hOur+KjoITaSiGj
fBVjv37gJKVQGR9a/wgBrU2zR83/kbBwaSJiMXBiLpZBihqikGzdQmmwV9R+9knSeaZqC8n1JhI3
kshQgquQTlaqS+bzP6WwdbolkSJcZ2US2ktTB0J7iYg4aBJAMbgWvT7oLEAD9e/kYQrqzK6SQbwG
cipW7+tImwzLFbNL30JKtIPLrAGeOidFdBB7jSo9c1Obw3mBlJMipsx5Mb8X7px/PKkn9YaP8x+q
PRQ/uXj2vwIJSaMo0vI6YtrzbkSuuj2LGgexlU0Cu/AuytSC9SU494Ju9zMoO8XJ6IMZaeVdWQkp
AYxXx+lhNyXiRIHCxafbLx5ia3vrbqlKRfGIxMOsR6fDEiKDZSifSxK1EyyChPEJZgJru0kRegx0
o5dQWF3CKJIxj1dzp3ULnKMMtcJvnCr+7hoRG1B1LqM9rTymeJl3O2M2BqfBCceg/yh4Ovg/LH++
LC8ztqeqfxY+MUCthfSWYsI6wyfWeEFegolS3mR81qOSeS2KeMSTis+z23vL1oZeL0OsAB3t5J53
58jghGP3ynzVzC6Wu9dBRZ/4u9mIXE2OSLhL76qGW+oVzVkOZnjwRZxD/ns1M+wXPCkAQkx/YbVQ
vSGyJjWEwasgQHMPiup2YWvzgOIhr7cqtTjrtzjFGT+r8/uJd7cg/97S+6cmJikQ/fExG9OEqgBw
hNWNaFChGi7Q3dCLestWRbTyQ6e/1KztQu/Ic29QkqHUjeUqwece6E8dqBPj/L8Xh3mA8onM6X5q
zd618Q54llcHnzIL4aRRPfn4Slb69BPpo/9mWGrpdAfGCOA5u1O35uvtq7LQ97v8ngMljA/m9HrF
Zf8wB7i68bFe0SvizOFz1FiEvEv4vJQvtYne+hS6N/vkp4oMW9fSIR2L2ZpwPqZ0yU+Dj8KSwGdp
Uu4Ckkh93xinYPThUhmkBZfR0mKsiaFcn5WY8XRouIp2IY/CTVcSFdPgKXFplRx23HLauReFmlXv
7x01xEQoewG/DyMzHoxQabb+qhE0wPQGY1Fzi6L+e6aRlQuNIlciyi7rBzRmQFq69GeSAHc+Vtol
LUGuWW3H94cJVTAO+BjruTJLU3SeSxTefd3vaIt1MXQ3Zif3ehp6UQFkaSa7c5YmvJAuE/BxnAMf
4b3Pn7jikIOEGjcxEC8wXqfwB2d8fKcwGwM7WFh7Bh7pNdoKBnf7Tp/SqUcIEjtvQSCP142APhjD
e++OPvVkvSPBSur/a/AKikL54FGeOm+r6oIknY6gL5P+IS+A48gB/ZvGoZ4up4N6ODSNu/Ncupcp
8O55uWD/Lbwl76RHT9bqb2q0nlszYUoaeoszM6EQ5+qiv9EmXyYtvCtCuGW/+fJCmDBsIp2EJptS
6vX1zGMt43+YeQCuqPO2Pv1Mpqjm0Q5r+t0uYNPzGLd63CngM+DckDSd/eNLdV2+Nj6L/jKs79ZC
496zZp5m6IYcqpac4HFYjMsqcIK5S/pYCZH2mqAFmwwQPDjZTKVV9fom5Xl947pCqU1Yh3uWyYOl
fMWlw0NeI7/F1Jum2LNRduUUZxIdSoutzJB6NS28w53iz0AbTu6KACcXt4WR8RxQ0gtRY4OAqE6c
GNofEvirjHZfi9qwUcwkVNqwUHMkdEboPKbnko8jVcvnEZYAqpthK6AdMk3697fMetglbl9g/pN2
FOCWUY3cUWUaL9C4wgiC8w3xvjM/X05a0tBROUSzYs82q//0y9EWrKKuYfWju6bOAyFsDfwPCluA
Bzd7W1CegswqLnpTtZxakmkZs1EznQdvqmyc4oa+0lIf7a4kVL8lkDvWjnTjidsGVLZITsQHvid9
Y7jwuefMspQS7fvgoSmIYkp9Hc8pxr4SKIxDS2daIXjGu4rIS1ZfBEVzbG75qfx8MLiRRV2+Dpwr
hl+uOxYQuCf6WNyHl7r1zx068b82um9FLqbCaZUO6VwtWEoHXgyEJDkcSd6mFpcXb4d4NngJw+54
oncAEHb2tepKI/4T9yqqURXW7QOXAb5Qq4+s6Ullk+SkzCsQLNCiT89KAJ6tbcyI3IbucFbBXOp4
spRrUWMGkXZv5oMOnOYOR59U9CH4JxEAgG+jTI8SYztplSaqNdCwsQx0deVWGJnQBg9NVUFc7aw4
4jTV8rBMbn7fw7lm42xam0KZ3MRtKlIPpmjJYptMQDiusLebpFNTkyVo16jfhh2A+JMSrFIlso8o
dSkzQEx5r/ZX1lHoWDcnY8ZK2oHJl2rhEqMRMu0Avlin/2T5awzDmv9ackKCJ6iPHsznEG2whpxU
zINAXp+UO7wIsTgjmeVVE5VF6Z21Rj/O02OKuS58ZQPg+Ba3vreYz+dBu+bP76iEzCFtW889mf1F
99sCuc987fW6B73yRuZ58RziK5TNlEmuL7T4OMczt/sC+RUMVkMoS9s6f7MYue4yZZmjCsJxnqkK
FFUNZJiMUbE/imf4e3apEiP5I2iNdOSIe7bHsFzthwkpwwt8HBt8+L6BF9JHAuhxshmr7Uijs58z
XzpZ1h5PU7bvprGkmM6AZVUto08twU/PHbT1Ww4UdBcrkuLOcqt9WzH4ZWAET6oxeCKnv5ZbRlAf
OZ+mo1xMvtpU37VR9AvEBf8vN/lcjz3KOXhTMVTWq3D36GLZ9/AAH3wPU1j+7Ondb1xjL2ip2SwD
1mRBNFDXFE22nHaLQghqkpy6vHS2inVqlVHmgRw1XAAgGB9HjdfhIA2oIwrRyHB6+pY5d2hUjcoe
hMEn8ARIMULLP5u1r1QBL+IpILeOi8XnXKOJKYGMiEywxz7gvYR1nFO28vnCNdUBtIAlMzvr6rcu
DBY1SHX84dsz/OQQChODiNJroJQUX5cG9dfDRflgA+xnhHn0FfXux6hVg7SvH3Y0SBU/Xeh0Hfct
iJ2STyp+8hOSmIPLqzQOT5NkB9BM4koQ9sZwOASi36pIikxCWEnqHgVasfGWi9cE3iBYg7Bft3ID
1/coOmApT6PLnV9KcY0eAbEcN3gK9PV9hV8qfrZSH/8m+t91D3B7htJ2Ml3qi25TQ59JIclVXXf6
jhmynAfOipecKXQtL4pTFVxeto/OgpXU+SLslGUpkh7DGWY2P7yR+xaEp/K+Q9xICB2pGK90NqJ1
z7B9mR2ULjAeRq/ydKw3kjACMg+b9M/qDxnbOHePhQjZYvH7+JWzg81yiqLVMAW7R+AsC8bo4T7s
qcfivqUUvsLA2GpcUUsrkqPif7lwXXS3gCGOS9lSc3dPcc9ReIhs5DYM/XR4Y6TiIxgVU75BXAkI
Kec5hMym4tB0xHX5IvuXQRCkl/Wq6vovBZjF9cNi18uZFSxkYgswCtfGDMrGkBkUt0wfIAn8oHrk
AqixAHKeQHFvY4qKmos9ZfRdvZbwvBeiWbAN6D8+vDLMIyW+tcKFP0ROMcpZgJVCKl1fYZy43QUU
dXQ/5yRxQaYFX9jcePl8UmaU4cDk6fvEasAuVK2VtYfdBEAsshdYXEL5FC6bRBkk8hFzNZfE1NWC
58ORayp0Q7HXGiTs1ImPju8CZ7yf3aZdqA3J3qozahEHX7tymfSVymQv9PIHCKaJLgeJdAuao18R
IsP8PALmUidNVcDykNkq6QKx+XaDyUAhAQuo4MQOvc6f5D4659uMH9nFhL/EsBWWSj8uoSxnG6U0
AZwHgkswczCumbsraY1fq8AN3px6nhHC/lherk3XNx8MTsTqlGBq3rhJ6DBKwUTCSOxMnSYa9DTl
7cxpxBWAOjhD+3uLwzgEs7NwJ0A9+aVOzg4aJr7mWyCrHCuPPhh7+JaFvHS5yNEv7RRjr5SDWzfV
dNfsCJqQjiL7V3kwT773obvWReCTNx6Z3QhvBR4wN0uL1zBO0gTdcGX3oO1hybsJHxtPMg/u6XTq
65O2UGno3k54lRgZWmfpNDCTgBM5oufiQ77afrFLEY+EJMWsUX6m4W5SKgeOVMCWLRLGu5iRnK08
p6lRdzw/Q5LYO3xdJMQ9R5tb951ytQ2LpFuiploYSrmrY4o0SpTy1dr3h/kn0vDuoArAc1NXp/IB
uplEmpVDADZxemkT8KSp8RCzFCoA1fY8zlDI8ug7Wi/BmEavIcJdQwvUDqbZCXooBWxGGCr9wz1I
4deHrSiR/4DKU7SjbGdP6rNTBleNFyxUiuAsEwsffJoDZfIgePS/NX+PoeXBSWmdVMd3Md8I8wMf
hhvo6ZY8pcq5Z50Oskuh2yIIWE0GOjc1MCk1mz2UwWuJ8h3lELbdfYipozBg2sirjDPnESGCwXjp
kuxnxqsg1aTUfkN4Si+diRMTyklU2vfjIRw6TcAzcffhalWQ9rVy6gRn2VEgg8Ie65Rff89bx7k7
0LH8E37dsaEqVBLTvtCNyd8VQVJCbppiTClLErdfCQok9ZOOMhEHbHa6z7iC/+FNsJVJ/yAsaHjU
PxcghcVIslqmsTHnUZb0ZpxGM0vWp7IgQ6qQPPcCRDe/Eftd6x3jDUF33gaSdS7HVtqCy3R8rPD8
lV07AEiGCp+AaQkPD3i6I+Fgb0Vyt1oxrJT/LfhOt7WuSXbM5xhhrsmVR7c7ULdDlPL+Orl+hUhF
GR9HMqRxcw4KK8h24Mn6l0k8bdU4wXzR9k3SSZWoG1mJECecg7YbJrXxAmZ+oGV9RZUHU6JrtMbX
BQ5DN55ElPFsB/OJKCQVCxwniVmM2ODElmD+wn2tJt5qDfcF6ZMBF0/tV09YVFC44gTws3Pnu+SG
Xl/U27ULUw4KWr1+VCm9YEnZtkv3/NtsofyrE1kmw5Fr3J1257pCK66ZVK4lJTtX5KdFSzstu9q9
E+5DWDQFwzBVKhDhAXFo8+zMVtfw3eWhwmO4qmtnrOPZf3xNkN5E1ok/JUIpy8KrIWm3aB8xbKTM
sHzVcQpnsOBgiPhNY3Rdnp5d1Rb89iGdmBmdDE6PYzHkIkKiq3pBwRhesRVyXkMdBAEtsa+weUcY
r+86FIOhCgK+lShfIxLSy3IowbsiuF5hsCk5ezz6VuNE50SgOE0q5HBH0lkaakF5o4C/xbpit/WP
GUsGJ4KjFfoWHrS9ZxRAscXzPbvAyuJYyAUtEcs0sNSQ4JGwsLgUMQK9lOKqeXoWnjlOv8/Jp7OI
gqibZV6UA5dHrfTq7b5/PnwI1fE9GuGiXmA2LPWtjahubesfaWpM/hUNaSLzt6esuYZ6HrUK+Xn6
BOnGGsIhJ8tnTvga3+UkClLj2ylEEykg8FwKPt0gu8PFtA0LMmR0pO6QfbjsvFHg5jQQXHDuYgam
GDPTDjljy4cGXvn3Gh+Ag1G0f/FojYLzOy0nLdAI9Co5dClFqqSPx2sCiCHqo2gkDH2qZAygAPAJ
l/4QuAmLX9YImfM+f100TcnNdWKvBzwGnbh3EVHFonpcjrbU2yXK9Kg0OiYb3qr0f2rIpEyc1Ov5
KT0URb1aIxMDxM609vxqQfIG72xbBKuoB0YdUnZvQmQIKG2hRfwwedEfB6swCINYZzCM+NeUEbAH
r7sJSyBEJuwqRJLDXxM9xM73nzxoYuFmCJPI5OaIwClyAOXjsl7Xs2XhfP7SswWnnjx5Z3h70hw4
E6ur1Kir2NyBwtBZP4cUC6t1QSqlAIGq+y0K/YN2lXE9jjfusuFsek6E0I6a8832gH4vbTFxgCEE
fz64lSya/HMyqSr1+14ui9Kd867uvqt/Z0XaIrjyWjgApEaBIkWd0ZBbgx3sJhKLMdB+G3c8yJIB
/l2botfYHALndTDj5V92oWeWx9gx4S9WQ7GbrbFnjLBsYa1Jn44hjtw0t+un8Q4Lx7hY6GAENamV
rDP7xpDvEdoryxOm19CERQjdmwM1hOYPfejUGqw4Qce8J/LL/BngPiuCY7S9/cD8QKO6126Y8oLl
UQRRyODRdvZlsNHyIgrKDqqdRxUCK4HR1E1LHwdQEe/hvmOww6xehNcECHJJcvMmcviD+BjxCBDy
Bh8Ehy9IlskT6UTVPh4Ibmtx4kLqkwszCrrbwv9Aj/iNdSPJCImpEw4OQLZjCt3hNM0W9GI4J/Ga
LfspaZd8tfSI/o2mK3vF8pDinWojvZBqhXFhQcbY6ni4zzFQe6ueIjorbALphXIVIuiGHbUZnTOu
qgEuP4Kbok9HRJ49aThaKXTm+xoP8M1HX/KWULHc0rKyr5MLWJl7tnIGIFDwDb7eX8EW21rG1YrX
q36pg/1wQHMIGEVB9dCK23mdVu2W4pFOMOsifEHdMdm1Lv9Txg9Ivb2HVkPqkRbfXLDcZUrdn1vs
vSmaRtoqDtD3HTMN7Dc5xB1rIGJ6lVO6tIjBZ7IXiCdhRzPepvGQhw0by009r6pJE5Eb1oHEY/hk
u/HAC7iG/RLYNZ2Zv2yxjc0AEKVyYzZswrb3AVmhphUiBEsdqq2UfpzBmRMFzaw2bhWXitOuVADD
C0qRJoRzFmftbqJG2F+ajNc1rhl9FBxmz6SBgQFgwC5WO6+Rw+xwCJgrCgQH6dWUNeRn8AFV98NA
ITW8YAIgkG2vm+e+IM56d3DVO8uu0myWW9S6hYXDo4FNSyrhy28GFVIWXwLm+xKTEdHS1jvDDD79
/CUZBGiFddK0wDXTq+vVOS3dTvhgWkSag3z+Tk+CQ6/0E9IpRQS2iP2q8ugq3davMbzlc3f0TGKn
xqm4RRLAy0xhTi+Txn3qn+tcOF9FG3ENpjYpb/Yz6o3ZEu2Pml3T2id+UtCfYBnT03R2GEE4dX5L
F/WcpqVX0CXXNlFlzyfnbQJL8yMUGLGXPBSp07oDbtnSbmLfFJ0+bVrXGmZ1OOmGCDeDb+auBOJv
a98CVKcxi7DamDIiiG41BNkOVyg+OAesQ2Vfi7d8a4ji1jGvnNswGJEJIF6GAytLyR9558PuVFCI
rO3jWCFgW+22VP8H1LpvIZBoiBpIJtnPZKKJhCbSW8YXCTRZlptng8789W2zRRIbFw74WS1n+e0z
rc78wf1dNoaRyQmuo5QCWVzIc8Qpc+BSdRWtQP57wh0nzGDBFdEdTPWPuUqQM52/lzAdXkHwfBi1
xjbct09KMQNxgoScjXh/le0ShEBFEQjRFSHoyyKSJg4NEK3CCXOKPFIqwLbNA1YeGYw6xBdMkR7x
OGRLvNQNxltz+qFW5F4O51wtE5ZufHb2jK74HFgB/CwgjlJxTkL3HSHI7jCmKi9aDuAQmojgUern
YyLBV/pvvlZS8bCQen4UAzevIiqI5pZvnKaOHo5rn1L3QjZHDFXsmQVYLZpgr8ECEDzGzTGY728E
jTQiV4+8k0EvymqTfSboRuaGpe/ZBIy5Yv3KVyMGfETgmrJLx/XXXFKMHxMYmO08mA0WIT4oHo+x
LYGwWCMPCbgW7+vThAj5zIoWqdtms3j2P/rLV9QaWAo8pNTv8pTnqM34F7mFmiOy7ST5YWOs7bL5
66WVp1Qu+hQawcNH1gFe8fHXBdZLaQgI8j3PdJ1vjkpaizqDYCh/46T38xm6oDsb9VEUNZYTk1Ph
Ahi2AsJ7Ghvx+oPiNTpqgOXuFfkY1AmV2knCws7G7qvzfTK7ajTcnHZeE4JBoomuDLP7oZgblQfe
5jbkIqMlrEhDpp0taY5Qgkuf2U3vCoC7WtG/e6REr3ZRN8/SFt1yGyOhhAzqAFNIoS2A0og0Om00
4O1LZtQd5q1Se6lwazoddWJt8idlchRrosHxwtGm681se8VNfDuiubwUF0E+sPicUIPaRYcBPL8q
o/H8g/AY/2hK42NCabIWjK1BNczWx/TZcC0R2OzrreVEWZ2dIcUXi3759ORCnqsFoxSE7MmqL1r0
pV4dYhW3ppKeZ1jNmXlF6mbdrNFqa6BXK03jlznSSc+HdDYq3/lQ7+ESRJKmxsYN8RkEnQzMTnGB
1gG9EN5SWLBTN3NJO8HiAPhXuPS1Zx4ZeLG/ld2ZkPNPZ2E0oaQBpDxHmDlJ5R84DmgtFGNH6FeK
iN81cZoa9av9Odu4aP6OH21fE4VP0N7xxWTw6oQzenAjGea3pikrZ6qpGEa55zOh5SZ9HnpyUjrd
+PwNrjp4OBamhWmkf4bN1gMZ6I65sWFZjslqy4BOnEl4FFC0k7VtjSKkekzLTC6mx/tDZUAoHR9u
LXGX+7S5TRRIZf3Jtgr7D58c0SV8/xZeHB5xMM4uRH1TPISk57qt8yMgSlCOp+bV/4Bh4qG/zMf1
70PWLwFA3DLkRYBLQBesCN8qJGUBGPppYmIayXrtSxZig2Hs4BbU6y0OR7SFQlhUzqOG8FJmAZK7
DWNbW1gDXclmtr5lG6qbtNNk2lHdGjkGl1KpyXkqX3md4Mh3DyzYZenagPBpxgA4aqV6QKIeFNZ+
TiTWIz4tHY17d89d7q3rUN+malLdMxbuJfBDTBpcqbgrO3XLMeSvX8hDy1vucswrAKc/n2ClU2J2
oaDxhofM1GSYr0WRuNi9V0c0fi0wsJVJk8G/lNqPN3wAg+Hd69+F0YTWzbgkDqGsMDp8VT3I21J4
Ll4xNU+ZC2xb9rizADOxWnHeTAM4osAL21VJvPaVBNC6CMbP+VDap82EYxL8eySz2uLZLxQpeBbZ
jArn1IIv3/dsRWUFDvexH4QN3/k91W31Q33MaCzwQIUee3sROPvAdmkg9j++IJVE0Y0fj+ud8Ln8
L/WIBAe7PZc6Qg2FvswEgCIhenpRxr1xt3M/aAq1RucHh12KLDPqfvI++zJkJxSki/0357B/uRao
ug0pVARu3Ss7bmrGSuJvM4tYIyVYnyd8oD2Eelbk3oFeTIgI6p013S78TK8Tz+DuVChidEibsXra
PuhA4JfiFU/P9XfhmG5B/x7f4aXEg6yHsBnmHcg3YgkYQucwvSaNlEbU5l8LHInZleq/3yST5B9q
7BsNmHTGC4WRhM8MdtGEoo6eJYzZcmCaFmv4ZO/NovkGBUoxtGHxA5BHgEsAe39GDIpx76kzO450
ZwD0sHR35z9q7BP+SaM9DgTI0iGFmDxHnfbyGYSc+TEDWdleiMVSS10t4XJ2AFUFu4Q13AZrnp/x
EzO9QCE+3Us+FlvhZIx9HCwANFC9YLbc0Wu+tXkxuDQCnqWflPJu55/+uRBuZyvhqHKoLrEheiKZ
w8RYuGbVBWb43hbjTxuroqhsKoFipdUWbHhk5kOc1qBImTq0L1s4FANQZP9xAaxg/c8ezrFQ0NOK
lfK/Z+1Fc/DdP4G/QV83gtbjW4Z8dXNuO8UwIhXoxo4zd+2KolbyF+YHbUhSbSIDXHzZWiK2DIKk
iFbw6jwNFabexW78cHSSQ8loMJXgpdX+ZOM9y37gJ0XmW6R0xVMK2Y/WY+ve85xz9/CIO5sUHld4
/m/Y1GZvH0VF5r0yW3U5s6It8A5WNoXWnCRdWFGzG3v7hYTruOK/+QoKYL9inm0C2aZEQfXA3WhN
A9kk7jZIRT72Y+JKKYdHhfiFMJYzsJ3u61vYJ98tjMkYuQgLIilIaXvTf8D28lNBD9jSZ/e9aEpm
Gof8g3XFSlCMbjl+2hetJippoJ3VsybSpXHdr9o6KDIUEdEbMNu2Cc+hGo9eO4MlIviM9efftKnr
TvscwP5lKWyJK9W5v+H/vPoc0Q9ajW/xtVROEASNOk1sc79x0po1VJieQYF6syWSlsXnsfs1lo9l
xc018OOXOVM8aXp6+xa2vYNQG3AL05+vvO/wUWsv/02GjszjhEuWlb4VES5jBNu0oNwn2cmUugOF
YI9ZJhCW0XupcX+Wy77KLI8OVNWmACfupPedcIEMhqyJW2Tb1EH4KmZ33yF14UyKZT6K2a72UAOi
GXFTR1at/53EdMSa6XWxwTuNYr8gWKwu14InBx1TVVaB7KuKeUniAvcLbVQrs8vYepuj0CNDcvGm
7fT8JoWwvjyKJhbrSOdi5cxdZmhKLCTdq4OeQy/1uDVYSK9x/cuhxfKrOg9NlVxHE8LrYCOV1Xyo
xCCy6oj6YQzoXuHCBrUBOCWZx2QwUx9n/Qi58Tsev/7vGfn1Y74E8/QJ0P1qbZWc/OlcD149bFq0
qRZI4uZnouT5dqJjR9XbCBjCbMMrlmsq387l46WmVH/AU0C8ea2VIu+g4voCg5xe6VYiRI1DgA30
n1JUlTA7xRkQrOwAkCHIP24AeuskjAgtvL9HL++gF0cZCOUHJMxXDWcld2Yp8Iyu77p8n0xt6JSf
gqLAssFeYUbz4LfMMU1oJG3OVJinAWpPSciR8U/5PaTyWvlDmeogVaQYGzD/ogCabDmxMjyqypQN
ukh6nFVuBdctNfj2vInSgdBZIcDrtIYq0iSEvDZXWiKPXD1Ag+ug+IHyHwKozOV7/+wvk3DLD1w5
iWbp1YAcPNzEzn+Rd0S08AFwMQVj/0/4IVuFBk904JBPlO0M8zZdnyLvs5oklPIN48Ln8DwlfB97
96M/6FMkrrmEoSn2Prgh+zWcjdf7DnH4CEDzvb27E0krMWVpow1o5skI6UV6omWynMgztEE5Ucit
rfoWec6TZA6jolXaZqa3DX9GXk3RAnOKSzqP9UcaoIqusn9URGC/nRvelRh0KcI0mMT5qiS2jpes
k+BLHjln1qMHzlS5LxVKx5LN++Xwjt26jwUUr8ek2b6AE49bKEJOR4yhqGL0BZUPn09Ysif3bAoc
Pz3mozurMrmqZ8Tw2c/YMpYjfEbhP0DNM+Fx6ybE/OmuoqL7OaCBgr3b4fzIHyscrOuQ+bshCVlG
SOkAUydXb8L92XYg5GeMGODf3dkuJ+HE3tpvWoeYshzQY5DDDeq5gizE83qq9//56EORc0PxjJ3w
g8al3T/F3OxYES1M+MfI5w03Ei8yTmH/Xii2ypdEgS1TSDG80fQrFs/WrgFGqTDTv5I2PW8Bhx9S
yHwxKrl3rES+Zy7gDnGnY4wKuQw+rLITKIZnEswxq6wa7nGPiSefJskKbDpd4nwm6aZu5+ID+DEB
K9tq0RLTDtAqfgbIpAkmx7+WMLzaFIAgTcTIzRgKPpwB2M/jBBzrW7qA5rciBSm7ZJNpUFJTQaIy
7sCdIwpR5mBc7jTv9TyBJcw3koD9DTH6RG2yWmVhl6ys/dgX1CF7BfMuVISjOv7EdC6Ss6gQumST
r/44V/a0SdPdS0BlMUfDQQ5hbNlULgFj/JppwvB904JeHFqyNd76klTeHyHOgNrQ/PNIX4VSlqh8
KPOJgVmizNX5C7E7xmr9C/wNu0zfpZQjdDsFqMYXXsP0zrv0ekFpKPy5uQfPy0uXfwIFaD3JPwNm
kItUCcGvZKNK3570DM/8h2bSwlP5+6U/YP61kiUGlibmbTchyhzqO+mId7G8mNJmYapZZimMuM57
Y8AmvsPI3FRRTCA0Ldd+zErrzCruFS6WSwPqXkr8hfCNGv+9tVHN7Xzyi92+p741IUbxochrlerJ
+w5hcX6XtU5zY2JajER9ZTQmM0RvkCfelKewlOLDxNwsU7wxHg+4SD80KOAR5Ueatb0Y3iueeKXs
T55z0F6Uux/Grna0Vc+c4giudYV3RzynPB5M/AAXAw0xEHeqFCRenScQEBpJNY6fuSLRzviHHm4R
T8bi/PXWhduq5XypGFBPXRVX+FE1Mw3A7cwZtBTRyXsx/3tThVv6wpjgErjOiemsZ7kH03Iosi0g
8I806Usc03dtyTdhiCcUPzxYTC1Ooj+SgMsXgJuCParY4rfkME2j83zrz2mdA2yiKtinWlbsh2kp
ddnS18g0FBcWooXtWKKI9RpEj15xY+yR2WUw1RhLS03yJ0ZtXY3sFJVSqc0/DpgGySDl6E0DSxjs
RccTzNfiQfDl6c8KnJ+wtdCMuxAorKG4/Zgx5kLMT6+ugBi3mfBuFb4i9nD3I3jsIwKmb0R0T5Cn
uxe0zKHvPudTz7zxeysUIJojbUkdgKK5+I01p2DZXlosscORbsrKMsA4Kq3iK8RfkDJ7CB5bDkkd
PSIp6ycsFL6dKDdj+CnbG4Pc6LjBCLmP4lsPrbyAheUbM0VGzFlGI8Z1sAQ+qRe6Bi+tGktXqnpH
ALhRNXSi7EqdW05a2eYlgyzihAiLvQS41l4s+AjwCU6lkYQY+9MtI5VRDGn7AFd97dOPUfg+s3Ky
ijsYkbZxpBr3aafkiSWeJK3v8kH1vh7fpA1JJQYLnc5vr5DiovTAwWWpF4ia23WTyPNJxQCHSgFB
pO0XQqsQ/BS/XtWWaozFhPUsHmKgQ1yQIjPoN5UPaA0kIs+PfzmYcJbBlNlBK6cPwV4mSKg0WY/V
/yrg69PhSG8MGyv5Fqx8C4ZnipkLs7mLIwhdouYSoRQwAJzKnSGEYK6kW7Cfum73fa2enjx/ZYCc
PYhIrcxFGyzaxBizl/p+i/NlnQ+yAIK6T8OtynQFrrCiGJdbtcIHAOsgoN28xngExvPX2TOhyS2s
OLr4j73tQnMmgrzInNwsPtuOLuJr8YcHvTh7pQ3V8BXn7GpePfSVZxFJQ23fOGDnMqCDgGViXPla
Uc6sPanTqNfyPP38ki6R63W+sDcc61WCXYdC9hoxrb+bPUaw6UXRBmxBoBKoQ43wYO9ugj9lgfsL
H8bxNnDclCEFrZJftB3kvZkgr7KA7cABClvkFImsntJvtvJKgR7RNFNgn66CAmIXKI6XGWytMOhz
2yGNFhzkkKPqKGps4bTyN2wBjuv4YsuYcwg/Hz46mIydImJeybgeanhvknvIqCS3eJL6Yasu+ulu
7GUfjcT9hm6ksRg6UHz3scewEOUr0Q7dpBixPsJs7BVREDs7fKuQWUZEetqsqC3N1Pj+eoRR+3mX
Lp7olq1EJK+pO2P+lqAl1U0flacAjHt11AKA3RYR1Uwo9yuHO01A68wWKrU9ied598uH3DQV8D68
DmOdsrgcSoiMARgsMKoobEiS5/khGL0BMckBIGasLJ8xx97AG6guQFbU6MyyL+NmiQWfPGRSNXk4
ob7wXpVVH4lHRoICcTtCZFj6hBNntMuWvUY1xXpxvfg6000+SLVgcBhGKtVlk/nLtVYFmpi2cYrn
I8Hvk1VwgINn31Z44TdhDxp4sYf/46iSrnz0M6NF2sKZYSInC7D9aUGY2DS63hVPBM6+6L6meQeC
9GeVtENeZfONQSa0Ir9k6nmOV6Ezq+2zvJrAObul6vOMD29TYbCYBNm1HteFZ1wK/1L+P8wNWcNL
vLGPnE3StnGVoEifr78pai5EgAo2x6VgcNkR4v9HKdbbrBlmYyFvOEyQ9tl1CsdRQp5/yWlWziU4
wJGkUcqZGxbeAUgO9R8cee/QeeyTiAp7GPdu713Qp1j1XxIQVfhOf+82qx0cAKuKpcKimN+8F5mC
YlXAy+zlzr5LygztsnwVFDvL0rzDo4Pen7yVjC4mf+EaESNn+4G2XblofqFQrGVzVp2PkRVouOrE
oFEZZU5SFljXvmi8SMyFeXAAalB/stO3ZtT2sts1iARtHLA5iqusI7v1vHI/RPO0KVPKU0r6ZSi7
/L/+7PHjZDXjjBtJDkPXnhNcz3cLhli7BrXp50zkwYFWvod7+I+B6cTR0671hLkKJlvwFiu3VN2i
iDB492CSuAOtLGTJXbnDrQ7zbpTQu2CptUW2d9XIb2f2Rn2UdoIQevxxkKHd3qe9i/X5o1Hj6Jlg
10aAz2E79RXKMKEEehZ43KDtWsGHakSAwOo2JtbK2GwY145h8BPG9viNN/KEuA9emcqAY6tSF4R+
E4oWwBKC+wMst4zpx9CIpsBewOeSAr1EX+cJ3feauF2xEuqK8j9+6Dp9qIW03m9+ysWMAYXM0UuK
HHswvyNYyH5a9LlX9Bl+VMAxogU1cZ/69JKl+LBRzP2yrOgTG2q6ubPSPtqJqooNVWDqEtop5N41
3HIxc+s6KyXmcKeaUO2R45yzhIc4Pp+1oqgkjJgsYFqMG+1g4g3gJ0DMjI0tbsml3sizazt7RbAN
zkWpD0D/RUrkn6njUayKxUIaGBGxkQjLT+zKgezX2EhmkYWu0i+bIzDnxcgf+J4RzAYbmN2S1mNL
y/cySaIWQWKm0nNGwppPYXVFwzmjML4Wasug2DtHTmnJF9iht5kuka/Gv66Yj0Ol1MlIurm5sPhD
KIclha0dw4R+I4UdllJ307CXShaTznk19TL7lkqPzSFuCkzU2m4rYxH1IjVO5u+EVFno7Fy8E/Z1
Xy9sej9PKlo/Us0IWAQuagLqeB02XNn0EBOk6/p52cihIM1Z3KQCAzPjiIUUqVgaqMezkXFlQxIB
zPyxR9/R9Azbj7e6ZoKLmtbnuaVPr4htQbA2h0r+HSIgCoDW2mxNLJqmilvLvJRXZDQgP/vUsqLy
OWPgdSDyK6Yruyj67tMaYPRhAtQAF5vqauW2YGeLYUaiuj3G4JKHklOx5hKbp4WLm/Ckh0HUZG7n
XPQxhEkAVde/teTizQBDjmPJBrvZeOSGrjS7mUcvCtqoL2cgTvNhiUfbz6ZmIBIP0/OSl5g0hZiR
c6dFJ7M6RuvD7J6XQ4SPjczY62j/HsbmbRKl081Li0Ao7I8BMhLEVY7z4N+YLJDTmE71mXoUIy2l
ctHqCqBhlLJGR1JYdZsDRMxmtFEG1d5RGWsHqTkZwhSLFmRQ741bcqHeUZNVN4gz7AbfvlfooQQd
yDehBY2QsbX2Zzz5LTu0Z0/sZiX9vMqaGtNOk4Dm86WWRWtIIsOsfJi+7WhsliVFbuxLoI786TwN
K+T+CqJXvTRpgsLpFYOfJBl/hOyF1pLLyXxsDDuBI9fW9uS/3jEJanLMtqrNTFSeWebK1YagSxSX
/22v5+bS48jzs8X49WSTTPuTyGEPgF9PUbzq0d3tvMAZneZNmk/PRpkCk5o+xrtbmkgY0nhpX3/Q
aM/1ANypaBjZMrJvn8QtLNvWfMESgQoidAQDedo391CXp2BnlnxYVVs6vH0PQyqfdur/zCvgxzPj
eFJJSJrqZQREEbNqQtQGi/YgB8ed07CbB5jSv0HN/cpVEbG7x5t4UO66pDejdJ804WiSRGw73ab4
UNo7PP0tqnDwGaTyI8YU9FFwnIln+V2XfqSYoEnopoHhBE7jTYnl7AyLgqOqA8/0tDJfpavGNhWF
OjYH675hs7+OAlPQPYfpPs8s1O5kG3JvynkzRAoIZev8ULyyBOg+bVasESX/ZexzPPSdsqqSovLW
Xh6uwfXpyGD9mXH9pTymtUpCD+FLdqL75pZRgdRWRki2F+8kDmVtjqZ2TcjLD6JOiCIkLZ4rH/Tb
cbd+TR64mI1zihgrE37Urp6N+FRZmfuTLCC5nk8i8mvlSX8YuQCcWQzLKaCAL2AwKq/ADEw8asmf
FBjHRiaJwU7METmX6FMFuX9m1Kgp3k6YPtBCn4pb/ojh9T6+zYUhGShbTB/5Gu51TDbdCCfg2Bpg
7xEDnC28gTGbOA8KHKxiIbBV8UNj3U+gLQBK62w4iaVRo6n0349FBPiSV0L+B0BciEfe2dJLs0mF
03WhOMjzxxntTP5Bv8cGHUYxERO4CAavuiVHvf56zaxrK5hq3iNT17TTRm1UzOprwR+hvVfK/kWI
BkUEw4Lpmt1ZudHYL9IHs3fdl68Gw8pzzD68YxjkmQm/9xbeETeTWx3mxTFNi7pbEJ2bjV3VksJT
BDVL+tbXNF5hWC6tta5vpqRzUG8WbHLutsGFCUOIQiOtEDkOo4VKegLjBY4I3rxcjbQySKgKu5db
bpbjspxuzHpbus7V/ZfdVUPB85GjDHmvgoeql4eKBC42dHsB6hEAgt9DECuTDQFaO4BTBmw5tfQT
bPh9QQT6jKW7R5AN6V5GVSARBfZSckL0Vtxh/0s4bOZLPKpM+dlaWOzMRMvyJsPJjBAVd8rVNKy5
5bUn9wmGaJQAvUkcg/pXDcNY7DIklpwxsTZnQW483KI6jIvj8BSBCaCMH49H8a03oGbjBnDIsPSg
KngDIhlaB2PUyM4xITol67i6P+gGGe2b2+tiM5+A85xUZBKUTBL85a+8f5QF7HZIRSZ9hmo15/u9
c5GmX6ffF5UoQgUHBOOtUMQzFtqjEaaEBwKQJZ/NzXzHhqLccPW7DLV8/4Vb9BbjxKqsIUVU/fMw
lOc3LN6MiilmOJZPcCySGlPNYaH9DmhjEO8vu0mAaiCjsmvzgSkhMBUd9+QpGSFEAJkRPkKVgxQM
BxtTdMvlhVbnx69EgWH6DPwkX4iiHw7p+/sCG235SKi3voMzCjC4UUla3LEOIparMJOFqbzyNQ8D
v7Ar/zwRTdHTAtVPmbEW+rBJL7+XlGDV5rBm/0IDE2ZRio5Dp8IzfpS6sD9R+ye3HIH62EmuaH8G
rcZsruQSbUnLR1UB3jUdYgtRA1tDAdlGernZVLzHBfH8eltmY+F6r1aSc7zw5e5XbHFYb5Jx+w+/
T4Ir1yj73wrp94lOkeEr93NDqO7AvpAB5W1+9GY586OeQgg2kK8uKSo/52U+LRrNhazrgJ5N06ky
QU4FNemsYyeczSXxxv2TYaUX7UUO4NNH/OijcIABSg3+94in2X5CmpDh79LQKDE55JtfysdZIXLl
RvDgHe7jYsmUBw8re1z96zx1IV9Z/9IE6jVz65a7vlmyUfqZ7s+0mmZWYo5U27+0kcUlHJjSuXlf
lTQs7nmkBK3rI/x4iW7rRIpyhMsaXWFDkXjc9eNKuvragKDFp9YppiD+Q36AkPTqta2kfkwg+7Q+
x+xojJFbbMz+20j5q1rDyiVdInXcPlsZwEflUVKQHCjl95Sz6mwC0vwrLkTWry05ZX176d5D9wR/
ZzmnG4waZdyj7pE/gJIThLyRNyvQ3WMN65Qw0gmCp/wiR9X2LpZ3o4uE564Z9hBXV7AdxWLiUb/5
zWEuRutdWTwNGYv25AnGeUgDYpeM5m2i/994AAGalJTKm76cyhnSJUzdkX8oPdtj80PzjPOKgsfM
7UcUNwEXKCRzyEbr6yjNycjJk9kGGfqdzkAP02aFd0o6zxy7rXGX+3i8v9wjGA7ltD2fbxcj9q9G
8jb9rbhBXRUKu2bP3Yp1qJH4VcVvvounqCzjFQhOd9sFbC/CL9G8PuvM128oNFa9/lmd/GdwGh14
pVZnR0vbjCC9m0R8SGmJOgLLLw8qLABnxzP7r7H/gmdQjRUnfzZXQGpbfqwApDK8MeywpV051obD
DADpwk0tWGHdA6WqvzeNXxr3EpOIXf0TOJwKy8Nh8yo2c6hRm8YBTLRmBlJor6U94SiRTgQ/d2o3
1cxHVEj64yqSiN6e/FNlfodAp8V2MhuF0mwbUAwBnWBl1yMIkZ6M56HIRME0NEvcdjzO+Gl1PGEt
D7gGl05b4BSDW1i5Mb3EKfBXhtGj1TjG2PUjuEGfH+rUsEKDcCIwMC1nsLE/74x+DLEGuIZKmDGN
B9g1+wLleQYy2nopU3Lm/gTx4oN3MUT7Pg8rPO3x6IcaDKF97NK9H8R0HjNGL9XfZPWPjljigUNY
nifzBX8RlZD5WN8ReaXSVDhm292CCpGpMPTSIlU/+yctQDeW+cTqvCWGsisYH9Ofgxfd/Ns5ycqG
DwlUr3z2xmW2aikjXz1yAaZrlTQqJuLMLb8fc2dApkw3d+5uYikut/gevRG6nsZAC6/zgKbQ9PAk
8LeluWTwuzK4Yos2lz/je8NX89myOpu8JxK98VyLYAj0sF0Yu3ePnHD7ILJwIwf+d0ovIP+SNEDd
RJyVDh3KdZO1XTrXkMsJZGktePR9RkED5FcS+KcPYscLiXzNteRV+O5HyDxsi1tYzWmiaf8ViN7T
4yGpQmf0eQYb8Mo9d/Onu1iNuz+Jq4Rj+nVsqDnF69bR72FSVWAe59sCNnPqgxv/wL95MkpbjsLT
ktwnXvLsho+Etqh2lWW+hbEMcYwQsUyJ9BV8YUzF/IrjalpHLQrMjyZnh376/6jZKRHQtFy6wImL
drnmbVGtowOw87OkZqtModQwrdkB/HE5L3i7/Ky2DPbO90zzVJtJA8jet4HeHsjjFZKfutPtacsg
dReOJbAt/NOiB8haHmqJ7uUHjGs5TbZw9agea8Xrq6uc5/QMTvmmP7XKHj4LMl5pGv7Q6DwkHYcf
Xc/B3iy+ZPuXQOdFmS0lyJEYtDB+JI7a1KdHGcp3ArXvVPu/7CVQDMhc6iOP+9iGNCFpUTRc3wpb
8jdQ+ALculWQ1wbGu9UKbuZMs1TPubY9NeX4zoj+BqT5A9QcyRozwcAj3bdSmWWMSu29KlndR1Ti
ObqJgYPFsDmUAiiIIqBoWGv+Iw2Xm6/yhhJcJDI+cSaZ5rTv++yFksfFOoUGBwYzhOL5LrzNHLVu
Cux4M2WjabXPA3fU7ao5vU6CrbmQQg4zFHFRGbxSnsknGfifAmUXBKwxaKo55kKRIpcDYF+adjN/
WECeRG2os/Z6/1fjYbNaxwD9nJ4JkI51rs/3IQI15cFodr+CVdInSqRKAiCGkga0nqf7zgwjHCtO
zBoVhGxU4rLSAZHt0dUsp+Ji6X7FtZdNdmV5jqJFZEWHvsHbD0A4dLHJpKrnMlSVUhxFu9a46nnJ
eIA3IdQo5OPOhj1Po2i3bymQitt4Nu8NRPoyTKke+dJX4MajPQF8ljzqBJd3BgzKgr7Drp0aX2Sd
D6HNzM9FzChTOc1F4grMmt2Z3V4+eaq9nA5NHo0eUr6b5nxbCCVzYrElh0aqIGs4+3E0/ubFZOgB
6vN1uLInNU1gudo5A+EhDU/BfFCL5+i09jBv+wQu+QycueOI46s/INshH0RJygpX3gYpMJcOaYSQ
FIyeBfoKpk1WQmy+C/YDy1k3YZuz3+XZjQQ4wz9FhQuCcVIlgRtCkZFRbPifdF3Bn2hT8oltAz9t
yROwSnCCv16irLA+XEe7AKFz2+D4bDDt0QWgNdn+d1WMaiL2NWFJ4/0lZJ2gzQyAuFxbL8phpMvJ
ARVqe35xDhNhxSwyZ3QNlexbJqndg9lhruCcUHb8yCmFJr0dXpbTjkYtzEc4aDYazrUDBBSB1Izx
/nkX1iNaowMBLGghWpPVV5ktUASSzOdpqaS5O/JhB7m6TWXr8ekz+HbMfql6HWcUe2pb7NQZxp9M
bGpoSyWjX/TP81+iAkAjLqZJbp/WrDESjHeS6A8nu926G6/NBsZEVcwdBOnio7GfDLk/avmwL0KQ
Obwmb5RnlJeTyN7cEaPzlgrd163xXHYhGv50PGUvMwb5EWG/ILm+2nnVw3/Gik3YuXY6T9AflUfj
c5MvAyTWKl2B9eW4LHoF80BhhaCSmjiXynjqFYTgORhPDp/oRIEvX5Z82n9lscUEEoM6wnoccL4f
80DmS/jgeu8dBHvQ9NH9YTdn/Vtshj84IjMB0VvWMyla9NbKFi9eBFpHdDsFXfWlmoKfqT3QPP4h
jNRKOKEw8EA86r8a1FaAX59NkUihaviQTg+4Ay8hZLpRdSnG5vTkgrP+q+MDfSWvnI1attRXobio
vIuNwcgf9N+0ws52oSvJ6zGBbyLdZxyIuo3edeThavtqIrMHU3ZXiImD8e4B/zDANXrA+LwGzdFh
+z0EA5+dKWZky8ccucbgLKCuVM18FxkIRBY2JyeKJrQU6rElCSGpYMoIvtJMSUEizRV4UZvXiVFK
YYptpIpM8aNfNMYGpmZ6NnklyHr+pUcd5BCSC81HfxMiif5fet2X1eou1kNSSDZPFqiPGmZdMWir
7XkiNAXIKhLKvz23s4/GB8nNHp08nvxspzLZtnXiASB06Gb6sAdUJ8X/lcjlWKGVEMENAlrN3s3K
x42oA1HiyqCkmvz7YmiCvV4pvk87Vpt7m9lzPlsNCC5T8AZymbiW9hGO9+21oyLoWNejxzS3itn3
Cs0caxmUwaIuPKwoqUGp/hADi2u5lL0T78F95R7l4VVBCV1E/+u4JlEYGKwEI7MdTp5lb8NLUakR
KySFkHMsZYw5wvFI0nbSrfZ/5qzqyzZdLyeZqEAl0RL19j4lCaASuk+7mPfTERRg6JzJhNdDe/TL
/NurV0dEYqXn19GWLo36Qzmtd7UFUEcJYNHqDpt9qTGDaJW7fooBVHjDBlKQ5vjNuy2HgvrThefC
W8cDiiYuDwQQYVb4DtfPX5N8yJFGbXlJi2Wh+oEzYpjlFxSbpcYlh5QyfKYIq1J8GhvJbHvNz68n
2216MRm5rGbTaIgOjOlu8AXC/uH0GMgyVmdcYIIQAIIUpPEHGXdRL7BHp+qlbpnXb6aSuWtNX2PL
G12AOldgBmVz0QnW+i7MDmMR6zsje9QyHfUNbQgkd3OCc6nrzx5wtX6njo6AwevXq4om1mW237va
KPJAfEXoTlBVyAkHa/Ui+ppuVKxjNbIjQOKq1YupZacQBO6BgDCeTne0oS/jN4ikrpjdX3Wsa0uz
/xx38pygGfWe1MreguUkVHoQRCIJkerRYuDpyEqZY8khbbw5snPR9xMmGwXATtIGeyQpfvo1rNVb
D+PS7SyuhHIPct7Bin+5QqTCx3UseUc6Kfq7lnR1E+yz5aCHUhfNjm5+WgoQe9LluKH3Rqb3yEfO
FlvuXp7L4OjgbECQZf3X95cxzeLfjOFxodwvSUFeNq9SLMwsIwRuGbM+h9FuVkZFSvsZ4yzLEXRX
mBW8d4bS0eDDxF0Hkdmp8GmOws3PjVygfcM43EbNYhmXId/4cGLkc92GROZNs0o69+pwJbg4eOTx
S0K4toi7LlgOJQ+gfQ/gcsWgv19E403Ktiih2rFbhPtHG2ZMOrnTJNtt2KT91brFsVIZhgB0GOcO
4YgYkB1g9qa9TgRCxt0DIGLYnytJGLEUj3e118Ric14lWEM7EteXVUGeVrXQofylH8Pn7yJ1A1zF
Yyo4UM5gE9PX+rj3EQpKSyygvYepsqtskyXtbEY9xIHkdKRyuNYDMc1nK1cJ3WVCHQugU6aSGonj
ioVhOeihJEPxmbmEeRRjH/d51tHxg9NQXa8qiyuTU8urUzsxVkBHqqAT4JEeinx2YBKFO+dYO+RR
YYkLPfxExD6JKV0pfEM5WgJMYFS4JDHelL8e1EbWSzqpMP8ammjhzLu6im3i3orM3W3yKyH48tEL
ZLn+Ug3l1rme0ZHKPTI0WQf8oLrmtSgd4N6NE94bK0Do3NWXDO0I1KC6H+yhUjqHMDKZOgMeHXyd
hzv4WB5lazTwdypvK1ojXSCqvaIkOVmAaTaQgOdC2Z3tgWGMlIqoth+I3q2yffMEtwam6rKss984
UDOOT0oRm81akW6uidgZgC2VLeSHZMT0mK+2PfVlOs1HTLtZ6T8MX8nidyIbElxKrRg8TvoluUB2
TTh3V0QfEBjPMfKn7oHEeyEVVg7A9loUwJWchyWMlh29mQZ6DIhP8zZAqm4ayN8na1bDf1wffFgS
MgF7uRepCnJjBPw9/eme7bLsxthPUnOaZjnSU2d68TlvNuFujHnJoQO9fXo3A45pZGLX4tF0tcuq
S+Y1fAbIMen2WW12gPqskkAZtSCNRhLn1epyprNk/dSvhFYZW8pHVK+9y4AIWam7+2Lp1WwlqM42
OVt4YVfMFIEVq27yhaZ2yFQkLF5jvfZKpaq3KmaEIUXqGvTRppcocGtoylIj1IyweWAk1LVLLRJi
DG0goPvyqKRakuZVOXmeeFi02qqmXrMvQbN2OoHf3OlIP0xXNxRth2HUcJIgrI1dAmeBl5nhhJcH
OUedrEiEMpaC34+DXxecCbA7vA/TNK51OjdEPNvb+igZ4X0z1uc1HlrvhP6lfNFuTd8cAsNs6aQ6
38uX9jypxOI1h8MFI+dSxFctyU1Sq8Pu/CEzNvr5+JmjtKdfIEqpXcfFVmXiK872c9iAvo5yVaUk
VJB4mYFHWAwrV4XtaucNtRczbsPjhROcszNHdNT1mcNk2uirNNTpZekIsbCZnOkllUZEAdtIBIMt
QAp+DbVOFjCgtf5sFhHDDWbjdDyrOSsjQrlFfLQTsJ5Sq406o+TWJXCbRwoviRlaXErYTp8oLtmw
QPknzJddWMvRE1E2iPynf2CwMn4S+DJuRHsuyrgi42Gb+3rvCHOeOxGh5ulWb3NWPRauN1OnUeLU
t785jTLDUCBujmZ+v6TWI6tCBjmXJSUSEGedxioFfQiPh+6rXhQGuDorB5wC8QKsZCxLeiM3EBry
StN4PEKBJZaFYUEWZTHgVYMzj3+hKRFmAMZ9Mkj9KDMBq3CbBGzjUZ+7uDnm9GztzpHs/E9EGx6L
MSEbWOsvQz5QdL70H1fUamTvNaK9GYE2AxU3ayGQ6dnTQc7+2xQSB9GjjJTqAIx3tXQuA8VFkl0F
gYZ3cwFdKUAZ826q7nVmxNPPdJGDEs+c876iE1ZuwoBk1niDHvGSymEA9T91njN/Z7CxoyHQAga0
NcLw1Xl7gdkBIdbK+2BfcFG8lGWei3o3p1QcoO6f8NpBWBIZ39mJzddnYhFZwtINXOJIfPsRntIQ
fMxyV0oJT3B0YNkB0+lZsB9SSrf4YYZ/uihYLVeUqxTuivjEKek9n5hzPUBPMSsbqtoaiwkThLFK
3axR3d7p3WEKoHjhziFeHvbjlT8QHhU6iLi+30RLX3aQH50s4q54SimG73ZuYANyUcorGt9Q72qI
8N2Cfq4aFw11dErQdM3heIbQTk6sn9C2hShUMz5cyjK+IBt1LaXQsObprnhGtbIDg+eJPLVAHkaM
Zmg2PzK0UNj6AGDGW78Pbrm7+Bb2dWskMMTSNHG1rZ4F5/x8EXFRbFZ1LBNLYPtiQvOCAtR0qF2o
N4NaDf3F34cqX1SYskJ4G7ovl/sD1D7EhESDjww/LJLbHckql/MzgU/Baf8Qa9CGftENSJGUwlJ1
hF2zkPk7wWndECYveQTJT+92lPieTB/UmBl1EIa5gy8FXb8gqCy5CXZU/q76r3lbwJo3rLksqVU/
txxeppxIoqSl6tIxW1vvlTx7r7JzhiNux/5JOmbzdGh21lxiFI+s5TJgW9DdDaqNRjVp0u6YJd4/
vHJ0qubvm8Pelnb58wDAYtLLRxKZt3+r2JCj41hbw4g1uMExdno6b0tRszfvWptYmdRxlyDN72XX
7aaHNtaRhcIbResI/QA0LYmRIR2B78xJ19R96g5BwjFTb9NoN3AsvXffOPUfPBANrhEFapwM/Lbp
vIWQ0vdNXRx0MegYGMBEw92/01h5JFGqzJpfxofC/YkzoLlTSn1DEVMyXP8uc3CrKn3DYNNTxmbV
Yg+/gA1MWDMLETHXa9STu9pKFt2YTmlXCuIOPYvySo/lZQ36VmEZqKjip4Ktn2C0lQsoBJ+M5wCZ
4SC7cjGwX5hot2THFWIw2EtbCb8EjbGaI77HOFZfgS/KNdys153lvZO5qarE5wNd2yZum94qvtUH
KQwyGuFgRv/iVe8qhlYHktaJChDx6GS1FIPm0+Wcctb//N4BIrmT7omwnVuu7CpGbaxwMlxv/RRW
GLTDLatiEaJ0Jp7GAQRrrnQnZSvKin7AVH7BHmZn/terH2UviwLXn1zOn2Ou8cpaXc+p61n6ufMn
hNTRyWWaiHktogLYBR/dO+2oubE2BqKvBVK9D0yJLdqeaVBG1Nm0lKQ3GoqJWbbeRbxCfXdgHNJK
cswDYRojqn5IHyzzT9FwXGykLzQbJWmdtZPmn9nrizOvmXEBpD+Vf1rFTB/U8ioBnNfLXRXyKA3Q
lPGy7L5tUBbxg5jnTZL7OP7ETvqONTQzx4bMIFUmKeY+MDKEPpsJ7+uCrU/OcoH5AQ2u9unnuRvB
VWeVTwb8Y1lJZeFpyl76Bpprh97HEGSNK+9UMVnbyYsbE0Vyu72q4EMJky/uwMA1j042FBbq2q4Z
G6DtQ3i8D4JsaUennXAigOva1fFbSQNv7T5BpGwBXTZPsaCsVoT292wWOSEhb5MMmCZy/Vj2Dn+f
VMKPkyDKLBu09JHX+CDuTFOyIHcPNQTtAIcf1seFOxWk9G5qmlZlL7NrzEMIEyNTrtlbqz0o3WD5
oppFbQuVV2XxBE7vyrMjXJ02DJd7AxpXSTkre/yanRqEv+cKvJNeOCstlC9CjRJ9ix3rZHA24aoh
p6x316fDDh9bWynlSCZIiyooxwHmFwlHnrCfAD4LqwPbMYVl/KPa4GDoSvlBSOGxOO6Gc1S8pWqJ
UBTuy1BYUvri/MB4Dm42qSZSdTHerUL8+Wm4ANAHvxs6TQ2FP0I7jSDO7nGh/Mb/8ys6bX8sMowu
Wr+QIbVMSK+2p/9Gyw8xPPufEQzc+/BTtLmanqZPeZJ1lt2usD4MmuoznAbxV+4JxOHs+siTyetN
0Snb+1b+tEnse0Z5jg/BiDfG70Rzu8QhZRRb9StTXAvzgErKIdi5OLncFaJJk9a3YEaD+LyPxwuE
PZkuW99743UANd6/joHcEMOuMhwsWOE2nNgn2COW6A3X9JCUALk87JGRXWFwLifFLQFH5ZL68VvQ
EODnFzB7iS64HD8cy93fiHr+H+l8CkKLyiyUrserMDbJW+Hako9z1C6Jmb6NUY9A6tOQdLleAcCI
UfnDXuf6C5zqvwDNVyEC1V3oB6B2LS7tldutKEzG/UkCJGCnmJEPOFmi+7r1/FHkDtXdNB8KDJgW
3oInxqmjSMhUalH/Rro3HixdmVlk2o8g3vacdGDzeWSzgoZbyaLAHm80fxz58Jp7k4Kvq6HQbLIK
NvzAYEezpoSH/RBbDknHwSqIaH7yyiegGzjSxMwABoE010340DENOVo+zSwd05q14263b3EUVJDO
zqLkRILyWBAQoI/vsGBrtvyuB1nLC+pHtckmfVZ95ViWCmj1diZPGpPeIJnLKHZ8B0FGQxLcpOpY
UHfl9Pv6Dyv2J4mkwWbw/FFPyaJANumwmoieQpGNb1uFGZ62Wv3Tea/OXpatDWMb7Lh/5OHpyP7O
RrJBYV5LMjMPRR7Qo0UWmO8Jbr0iOhjS6eipdCkRdm1vARR2683GydPLVlTOYgiOc/CLtT6pjw2u
/0rKFyov+THQ3eAsBZkaUSdJW9ne/RirLHtCYV507rLRIIKdopdy9r7vfLan5CripuelAAkcttCu
9pV+knFLJteIvLZP4scj1jgjvilY0tovlcaZZA5zBOTpzhP7knuYGzbhLwR++6mT9Z6Ath6Wju50
qCMphlJZ/v5MarJT1EMJwqPPImsBs4QLdOAxMpQ0DK8ClZelGAr+rYB8CEOJatcmueqHFzagf2Ln
7FA0D9JElBa8/ubn0nY/ZQKR2fSM1mbfFDpID/GCPa0sOv0AEOSLSPuOXc7++MRlS9hU5IoTSbaD
cPj55GE+DWKXvmqch0Qc0OcWikCI67l80QZUWqVTwAHnFoIjk56MWTk3qljqD2IF2c+WMWxqSm7a
dPyCyCIQr1ufJ6Rg89Bi0w9zpL6vI3hqbCQhpHOue1WIE+spNHlTutEQ+2iy+TFFnN022YmBUABk
JKnOffEyaz2u48GyMRR4pI1hxdiHxRq8VJsWHhpMKj1yX+CXCDW1f4jnuvu2M0JJEX0disYx+7Uq
eOv7oaFvaiyK+q1za5Imqc5WvVmMMmQ/Un2fLgIXGAtzdXwmxVPI8TayvybzJvIiCpUtxWr7bT1j
+zaKJ00sSqpf1aDcyQ2LTyzcas/KdbfJp4mt6/rcrrt0ZmdLDkm2L5sRCJby2w3HtqureT3ILy6U
/DBRsCkIDUA4sB+Cqdkb/rwXHv2IqgpCX62HhjYxb4rVLr70y+Ol4r/7LaG6706MlCec/c7ZZk0i
pxmSoQLaPzRrZjw2LqLST19Aqn0rhy3ugCUl7iZ/xAeVqQaZCgeiZfusLhOdTVt2KsARrzM0ksWn
i0zfIRdz3T52d/ZW3bdrYBqsm/WGKnKFLaR8f9ucErw0zP38vIjYE6MX1jbZmpyM++SHGAXys5ca
18ptirg+FqD9Uh9U8G586RfmhWI3OSOc/knX4VvQ3e62xj9r5Uv7qvUIvs2KWRzNaAOYeMbAhlb5
zy9iGr4t1vLoIJdJcCm0Q5urGolYVON+EU4JHMPuaW6IrpmbeC4pMzk5sJMykCllLHUyW9aC5qz/
J8+JpU+r5Fia7Oof5TBUP9Inyr564iBaPUTbNTJhH5rdrp3hUQcpzWp3PEvmW/l45ufDR3rH5S3U
PhAPeoHNwayAW1zyE05W5Mq2f4DRkvo0VQ4un1Fwt2jeIMTFQtLTP7ss1hNsTY4WU3CfSodUqfdL
/CuAz/AuqGl7bl4uCLmnZYCXLN1IptAtqbuDQ3LEe/O3XQlYyqIgJktLO6t1bDXiDHgCQ1p7rCmu
2cYX7UX2tmYT3EDYsEUDHi0FCpDAw0nCHYJl+JMKX8Au6Hi/6Xk9Gqi18WUJy2YQQQ/qLr/kq/0r
phy5YLxsyt1tAvZqn9oaYUo3aqgTAZ872vRsKz/nd5uzomQ5d3IeDUIUDhU+oNpjVQ26joYP6c0b
xCl9y1ulLckm7qYudvf1m0ZiXlmWIk98MlOwSYHStsiNdnC4GgbRROxBLnG4jBjluXYOFWLFfyIK
fjShQ5gsdwFFUBg87Gp5gXcgbqwzhRzuLi9gI4GE1niQNugPCCW/fAnLLccQqnED3hExqEPcWTE5
z7LDnp0iNaqirqHvTRjclA9oH3E9F6L3h74X4RYahqgd/pcGTWv2TPYdQvkgwvzXfPF24qlOUE4n
5LMPB86GnHr228pWK8BOFq1wjc23+IKMxDMvqhsXCCV1oyCOyihvPSR/Q1vYUYegh6qhb/Xq7+yv
XstJXRhCGMSQS+y/+61DbFIEo/pm/nAFVsGhHySQom+1q9IWvHlRN2/VJEag0Z3SdqnFp3jtNdN6
1gVni3agIREkNAtcV3uKNIWNe40Q64LuplHrYa1dssUOFNU1JquRm242vb1xHembQjNpa+zb73cA
JJObEyiebpjbpZjWSwmhNMyxsPzQtfVpOCHwEfsk7sx/nEDZcJd6ltQ/GFN/KPUbNTuJeZBVNoqf
Jf+WZy5s0dwpOf7M8pB//fQk8irKbOdJ8nQFLCHmzjC4/q9ARZZVV5VjuDW1HWgewrJE0zVjCHAD
YDZEZqdt9F7QkEy6BKa+K5rZzcplUnG1itVxFbliiIMWZu/E4qFjKk0F0K4KhSXEDmOGHNdRaAuM
cREHOrflioZmSOGXhvzovLqe5XWGtO5ZUg1+ZdlJo3ThXfryg6GS7gZqW2qOk3MHbMfxoAXymy/x
3pyHcKpC1c6MBeaqZaSDScxCb5vkhPRW++/x4HLfuWoT/6XrfE9Jmx9VnzDxTOBLitxTV+8sxrzk
w30NuXlms1OsVvVU6ZmOqQtBZhl6ZSz6PjFevHq6Urtji0vr73bTYr39W774mYXjY2A9lr9rGwKT
wt2jH65QXEnF+8UF148f0Nt2EVLgUr4PBMRUcC+x6ynPnCmvypPuV1v0qXQ7+BNvX9Fp5UUQFnyz
5CIrxLyAAWLh5+AUEcCR324QAQwrLABhsH3LZrdGfANjsRDLJ8EYsG8ZEzC/7fcYf8zUM2RH5xkr
6+xwaEizTelJRyNbzWQIbEIWHmI+7Fol0H6yiOVHZroWnkH0nZqHQJ+L8cRXgLWgCvSvNE8P4gNp
l3My2DGyhYCQNlchYR0urICwvpeaRblSqixa+ll0yN2GlsU05IYCWey+/m3bspsP89/jzV/W381r
JQ65S8wr1yvlDX9Jv4E7+J/aaOTG5GOMVTB4HAi5qfDTkZ+dmHzC0ueUvSGrahRBEIL5oqHv7NcV
lbXh7JW6e+I6BIyZ1CfI2o6rucE5MD+nYAca0wOcS8niAmaZK5Pbk2v0m+wEzrGsH1PDf3xqlrIY
uKUCK3c5RItpmq6hY4DGFOX9moyMm4S64V/e08Xk//YbBfvARAYIJ1QyXpYQfnhQtnec6mUtkyGK
1kEDSb6AZhcuUxpnC8NNPXmWlli0fFTS3KEZvE3/n9pORf0dPliaiAwNc0Abyw68vX5+U2E5Rra+
2Spa7sjuUPwqoTwmKpaXtjDUDM0lx/saUY0LHdj4chpK5t2z0v8+VSbV7ThUr+zHGwfcqxEt+BFi
w2luEHoRRl9gkXHzdQ1v5Q1VQvJ7gToyWuJY1d6K0/hNmWghQfgsYymVq2gAIlw9bWkxGXYMxcgg
voUjzFTlEJ+/0+oVTw5GPkGyJ+gYIKKHUVAP5BcrPjfSytTAsTLATfWmeps/PAICNtCJ/TBF+NWd
jKWEJsyO43+GMSAwmiDjDwKb7qGL306nOcoy0fCEvzbBsjtiJ5BWLsTnJdJoEuViQazeTP86Vrzu
kHKI8v1qgoHWFub5a6d3PvxjRqNzrnDJzSHIacY2Zp7Es23TjYcA7gLZkPTweQLHwHoC/pWqq7BI
ooyG8URoy6zgcTQ+ui5MYyKiU9CgTNFMpCWQegGGuXeKElwJyLRXOhIVsvlsdfyfj6vPz91UBEL8
h6xzT4WeK17WBOyDy0frMBhX/ZjqGHiYbKiSCW+qF22lmK5ooK599s7RRhXlK83Bd9ABnTa5tjqs
u+f1pgAEkaNSIHxNSKqNQG9IzozXwtmGMb46VxRzSgA6Vvi0uAvrN6QcdbylCCLO1yF3dVWXRZEA
4Q7Xu9eTIvMaat2P1tOM6PgNj5w5sgM+5JlwxUK4TAoIspf4tFauniAIsmKaFU1I2keV0ON1XVve
SoiAJyLQHvyX7z5WcYLH6up+jVrCq/qTFarHkYqht2IwjrEXrvFJpMKH43CwrkgRuSuKxaEN5L53
vabASC7xLZzof7CzGwbQP42JBMPRtJuSdABsk6rlV1mNEw17VLHnMx4i5zEIDcQvOlX3pcHjfz+M
ekeqtWjoRzrRnuxr6NfCOcrGqxNMoDf3lrMq1sCAvuOuzl5AAD0TGE1AH+91hS8Eo4mzvlkIHyXS
V7V4uTCYbUknFhcLbMis6rpgEsN7AbRWwbB2pLv4VBL0mjycGd3Md92JiLrJgUXaytd6drZUdSWi
fIQRMFQw0t5dynjcU8euw7jxSFzXloeAZwIn0Y+RVrmLCJp07F0cntMdEc9FJjQsbLMqaWhFdapl
raWKUtsiaWAHd8sbdKmM1fhe4bdQwdNtT9o3dsKkuiB9Fw72n1VrY9z0Z8DaeojeTON74sB+VqOc
mH0d/0+73NpcGmuIk+VHkqNikuoH/j39uLNl8crbX3Ier/Bn9KVKD8vthV8kqQ+TDvNyn4oQw7Ms
6YyWqzZ6ZtjLjJn3YxX4IKfHCFFf5gadvpcw7iC94Zms4eYgO+YdTdtobB3cqgjFWm8yOFJBuSuV
B2J8k/+6SKzeK53eiD31zjE0nRa9OyAecJK04RgVfQfzHwC7Ow2e7R5RTEzeUl2sjVFXKpjVeGqV
wa23XK/Fti+7Jyt9ZCzhuSBjnzUrYaIifSlGlGHYvsG9ajw6xlxYtUJBO6Ct8zwUAKUPaf9ODQ2A
9HWJNojCyJgIdFnJXAeMtmNOzKp7N+ZdBoGLmCktig9HsNVqgJY0/OQIeV+sEPl1VW21yMu/D/o3
6QQ2Z5EUP8TIBldCAPkhmo7DS7aU2nZFN+mfbR8Z14bl/uXIVtfFNUzgow7/98JzvdGYW1B5bJNj
kaFaP2T8269AdrhYL/kJBLFvMHFmE7Hwa/LTToiev9aOY7ben5uGOIZtPXU2vpyDtnyQVX1WO7Tb
klR/g3/k28PnaBeyK7eVI9E32htJ5N1rmte5b/vWWjvEtREOylnk/HuK2lCm7Q9HwVIbMPig2B3j
EimcQWStp7f8iihm8XTZSR2PQCzZR0Ym9mwqEW5wScqZUn3XpnRTnpsXab9cpff1IHtf0NvZIkw+
KfNLhWJwGTHw7tjxCAO4NwCaioptIl+FOX0X9sT4yLuhgp4/lAl4+lav89OEbaKqyToc3ZjxnfP1
ye/uheYa92kljgkRYkCNMmDYPCmCD4faODlSjnAUOaohyVHA1O5s76lLGOh73+SaiClrrIhx3Jw1
3dO5MVtLjVA7GjThRS8C64fYecsbqQlECY1r6HmL71owraJ7fkeh38QvxpXPSpE7wrTsVcnjW48x
fB9krLc1YpeTJ6rvj8LnX5uKQL0/aV6PZajTDP7zA35+byqHNgBgbnCwxToD14/YqccjcKI/QvbH
8MReaTHB0L9L2ATAINj7V5tisSAejxJwsOwLDTF6XkRABrS99hdCaE4Aj5VAbjRG6dCKCGA3KyTf
ZOrzOZXLhsSChNrx1heeVYuqGCZmZZx4kojL6jCoyJolW00BKDUBNpZ9yf/bxLTrpCpA61W0xayt
aPUA83/va2fgtMZYYbUh4HlTgJnYDIjnZvOP87hj3sTLUiy5hjkyE+6DXRdLsfJlcVa+Mi1jgwfq
6jqZhyPrWfsQ0sFon1/OoNI/lg6osAYlzLB8rb7jPtEsncGPEvNFYxAqIVfsjJWybXlVmq3pApzj
uXkgEyW+ZAj5Mo9u9g/hMKWIPUkkmGpHhjW4JqqHyqDmNXbp2adWkQzEWt0U0z1bt2jp2OgFYZM4
Qpt5j4NBUNxIZC3BDDFhlOzDWMfNRIydnpVFtBWLW2zIilkFSCWddPyr75trim7SbT02CAleLV04
qq2jhcR1CWJxPh0jTsbyLpwWNfx8dzUUT7nCi8O66A20FrrijlB+5aFpmeSENLltwd3xtVWoAGB2
qIgUEsC7iQusek1wbZmCLSFmAsqFRPjql28gV1t1LQurT8QBeglSfYbkDCiaHiHdW6DcCRGaB0Ia
311P0KmsCO2eBPpkJwW52hsw/grdMUVcx0cxbCPNp0PnX95zikjnlbQOV5foFY7RPKHLV1bXG6CK
gPO8WNYUN235usz1opawNuzISdpxCn29Ls16VAD6mCj/RzFHS7sFqZlZwF49F2EQMV7CdnBCnRqq
GT4po5Gos1jglmCHxffbh+dpZC966vu+SBmJz+QIREJtDddFfaew3MnYWGlCPmp7Om46FTQ9OkHD
sLuMGBWu3YB85ct7c1Jpw5ZbHimbmtLVZRRfMG3C3VL4EiaF0fVHuxZB72rBzV9/i0NCRg5v2eN6
7hYjXNlRDwH4mhKOWb0wd7jqM1ifE3FbKymskxl64lrYAisvBByvq6/jfeOousvn8ETfL7ff2FSq
S70h5dMIq19iz39xFdQiu8d4IvVxSLZbYdVlz9e5Gvb8vV9rfIwVAYVgSXS3qGfSKYX4cTirdFUU
9U9lji49o+OTZNz6byAW0/CGQjz4UcTaVqcdMXzV/V40PvnCQJn5JQHt45O+kTung3du2EA+/6Ja
0mU7lQduDP704KyyB8b28UjPSwUchuSCdA84SNjGMgTi0+Ux+bMIsoZ4x9UXkzgK6iaRUdvPNCrU
zQNUyXinIvQe8+bRsR0c5SVC6CCPrcSPTfaHkviRW3NbgDsCs/RKfXj5oeJ8PmX8NEoOApRojq4i
OMmY05r8aEJvgj/yXR86B4sQWvxiX6BE8EkZcElHvzljubgQtRYGL/18tlAxBBYGs2M1CSwrnNIp
amhQivcHSbRA0yxwjhhtb6x+WA7vOXxIR1d8lX7zSCa8paOam+CvX1jzHP0g5wjmwddmhvjqgbDE
boYH64g6vYDsyk/QG/earzm0NkzNHIqVEdX7Mbytkq6nze4tejfb9ifiWaOQqcf4g6V7LbtXwVuI
Q4L3E0/e+iGhpblWne7BeDudKM3KNt7rr8zSffMFlYTJpdHOgOufWEX6rYgWLQvxMv+SD/jWyZET
LTFQ+OB25TlNH41B46g1/vgPrlaXdUXD7wxXOSH9xgESQbEqn+4mI7tNGgbOQkt3FCM/285jJEth
V7jLy9ZphaV3Xs+3DVd/4P79zyzMpUtb2f3RjWobjG4dEWSq03RX2RoJ1ovaJ0ESSYdHqGzJpFin
ZVy7d22BVxgEhxBFyS9420KfiRB9RWxfXkTNAnNflvc8xlfLjtYI5qrbt1+1tuNQkd3NHZQYZqLI
21r4CDa2XDih4CP7H7T/Npk2CBxUPpgOFAqODjA0cEtasgAf1p2BVCqIJD0ymZnLkuVGNW9K+SrA
21BFz/aJvXE6wWTn04wfnHFYeVz0vrG+QBaRy6/au/9rJMYnYQMvRdXhw5FSL/yD/e3D/jyEeBNQ
qkjnv7YXeZFyIm1caKY9HCic+S1PtPNs1bN3hyuo94t7WTwc4Bv8/qBydltFKWpHsa28mMbXNjKL
fuIqV/ALQNmNsF584Ud47z9XfHYRp1EiIGR8CzIkW54qgseZYdRwZzlAZDfnRPSB9ctxjXtFGEri
+eNEvDsdmMvnp4rVDiT/x5bfWotNVYzh2I+XslZp5CUnkTCRX+ToYpSq6jJdaXG2sNEjrIvRWXgI
VL+A52z457Aqga0Lw0SK2ivjRKAA94w+WzY97EFuhhEQBelCtSe2Ih3j9RiN86GcZS6I0dCuWZgd
FSW9Qr+xQUPbNO+MPqZsOP+r5O8vHz6Nuz7bUCAYQVyF1XT9c+Vh+CZdyLGUQxOps4qBeMNiepfn
0HvapuDFyNR45V4yl6XrrwFd5GhhefSSdm2LktZTycG/OPfhnOn7bnZuTr0UHR0yQJvR6uJlPUp2
hi1Uj9vUjWeK08pxEJOHQ4ob8mXlC3BbZdkVXDL7tYt8uJNqEKE5bMjQ6tMtnDff5+6qj89tUkw2
BRbzkgaeGykpVI4Gw6bvRl/swF1j9eiWqLzQawLp4WZ8/cRK2aRGP9s+SuHMzSDU6jyTsr0h5kZ5
cajL8l21OrcoqdhtiRLD10OS13TS4q7AyEE2i75gGeS3uVxnBmG98nh0VlpefY4pWUURw2S7SuUr
nLCYbx4aY5/YcziTyav3mweqOerjb7GCz/6wUTMi51uVoNJuf0lPCz1KR7xayrQ0hChNRSesl/OC
Biudvliw+moKjhGa4PdN8nMnzdsCbDDt/Ayv4ctbBmSR1JVABMaoprDSKX9QEpzpnw/pOHcCQD49
V1TqThsp8eJPseZr0s7tg96fI1V2HrsTjxb/bu65L5OJGPxuvmV3gyqewkRfLBTCQN95CLCvuv63
MjZG3Z80bDq49zh7pKzrJ25328fDbAKRxc4ALRUhWmuhoB4F8gEmHjK77JNQTJph128b0MTR9V0e
p8/bB2dK6b3aWljF8SuBJTVRHG0IVRI/JlPEZ46O1FMAq2FThP/3SsTLmmfwmDUEM9NuppWT5KXN
WJDXh549rmX3Vk9GKnlKpSIg3QQY6H3aGv4aVJ8ClaGyE1qQPMF9gAalYdOA3O2koBCIDoHQklCH
LwE9opwmn84gRqefm1Elz0VnQyckn9rJ+/NhaeirsnBhehssl8l3LSxzufyOqANxXeylyOMcibD8
WXfA7qs+v2R4wKqL1Sxe4fTEKPnXr2RD6/YtwFG0A9ReLI2STrzEClq0gsQlb+oV0e3Cfvq1vgVm
V2Sev4iJx74ui3ILcYqiJXFdKuydvJW34UcPFpQU8lSLJzWA6Vx3/6Ku8IWfGeBxe45hR/s0J0Ca
H2Ry5W1uEsfK8mNqin79/XKqpNik2Hq2Yguw/4Cr1gD5h5/T8oIR5DDeNEWcMRtTSzDgmSXhXHYl
foWeGxBhy88DRRf27WhppxQDH9SE2mwsjvPaoMSAND3CY2zjBR5hd72nhpjUN/hVcQUl44vTRanj
BXGKvMPSQlz+5rskTbBtmubm9yjX+CJ5xAoqzi/jW4JQZM7zjqBC6S+L7gwmoXU2X++9XmOBsjgF
eKcnFBvr6O7qSwBmovXEuGo1gELVzahvkSoatnZGND0xjheccno9wStxFvM3kmH9tN9Wfwg9ISKz
ZKrm9y+aDdCtI01pqIi2UFUjNoMr0Q5xC64qE8vcJ0Wg6RQlDv4DLTzwg2OifguCCZplMdgJ88kp
ieQ7zJwyl1HZVwgUIALwnzKdgdT06Lq6ymFLU9GlARoucBmAv6DrJ0/X7VanmFQcEfjNit36HlQM
k+7LnVxpoE5/p99na1bv4mMTOy3Hdi1uY3G2LYZgr+OiZzBNOVVarrufsXmRNCAiIJRJHu/Z3ceJ
TQ8HRviz8vZICSeUCvBgddstIZ2GJqMVsJHCsgXiu2/hFtsCd0vFodixv2R1i7X5LqCLRAcyrT4+
4/ehC2QZDk/u2HY4EmuQF5NSFf+lRJsTW6GilUXLPT0ifNd9tmnYnMfHNt1B+hWsjxKkx7cbtabM
OmYC4sNZ1uFvSmhOwvdBHH+RMP5PzSQGcfpGVe8SfYMAJWKsODU4psiJP2kiM4fLLzTK8/gtTJoX
S9qE85zjxtDJA7vUgQQOC3VzMot46omskPUYM9HgME3HlPdV9hXhfmCz15kJ7tZvflG9jZ2v2FK1
xO3fyD+IcNmHKvbuvT3YzXN6HKXk9mQfS+aNjP/aGZ3tc/6+IXmiEYq61D62Soa7enVCCtpCdRCs
wBEi5D0mmagY4zUmQqWLVYI278j+MemXd5sxMTA47NUEuAPwAEguFbttnP7l7YKuIQga5+KJcexR
zRq5hD24zNDqRUuTtY66rzFUyBCnicbXjMnorGgKgVi/EiuPAf/4gasqPfFkDXVQ023W4FluEo6E
o4skZ3TfwVgp0rayfStaeIyAJ1gZqu5Qgfm4uJy4jlXq6y+s//YQ3zh/XaqiIx5skhM6O6twRi2H
gzfkenpOvl056d5Oi7jCte84h0c9DSj21PZrAyfn9f/hGYo2a2Yy/PpWC2LsD6Bu/4BPXD1Y4H3b
BvPnZXW5phc40lFPoRc1sKPxLAiOx0HnjzRe8266pbZPkrrOnKttXY2daYN7M7x9jDjUTNpMfUIZ
b0WRjd0UGUcCMliJ33Ndw6CAjAhPsFwy+zWen8bP0o8Bq+Ufo3l6MsQvbl1pEXebG1jvBWtYlttS
58vgoVD+w6Qbf32/fWlRfeD4fUyHtJRSxmhKRQ1S2qtUo8kAn34kN4j39HWyf5d4viFjodpBEfnT
uOsFwlw4+l8tMhlANLi+Imfvn8bgQF466/XsUUg6NeWtmCWUBn2JJ52VW4VtekJY8Ajxe+r7GEv3
5JVh/7RhRjeNfxCyjX457HbPS72qc42xYIdk7qyrxNnGHrOS6AnyrgJ/tpyjMV32uI8tuhOGF6SH
bjdeMOt/NiLmgmfbEJngzom2P4WWeKDJfJJy/4mOEIj2yOwkGN+vB/DJFMpSfE3pC6jSVIhO0HGs
fS0uQk9lBMe8UAgBDLVRZOY1J9wVG3g3lggnWwmsbSL7t8NJhaSUa3WsmiMrhh2iFRMluVNiSX86
ltoYc51Jgk5WdvbDLmEW/ClFi94cSaGNYFgBXcav++OCk2eziwjolb3Mhl4dzgcLqnOKWahwvu+i
2IXyRFJEyg8uZEw1/EiHwwpU5aKTYMHUVS010K9jnh+Stwe+08l/4dztwrApjRWyviKHAPVP7j8V
Z/8Jy7jQkBckT44ScM+awCICTpTHYbSn8Vp8LiIEBDHr1pna04So5rpW1kk7Iv6DrPLBrwQIueNa
kIflUVDUnnJ6CGflVmFNpVTeP/PJT/VAs8psyTMsYuN0xDo+sUF7FwJr3MOUBFYVg4FHz1aPU7sW
o4uOB+G5FMsZP+zaGVKQ5240Ud7+ME9vbAJTZDEBAcaMJqnN+sJFuE0RL9cCEe1GjEFBJB2DAMFg
WQExAVsmh2a4nm+a75rebIQFB6ITvXswPLAk9fZKMDgdXh5vfvirzEyjsOu9zFCzsDIZhYg1Nb3E
48FoM1OeJXsEC+ZGPJkxP9o+9Mv2ArWjiXkWy3Q5/ciwyIAom1NyrVpTcfVmsWRYi3QEjYq+LGgj
6JYqv9C/O0AdYJ9CrFoFApJKsdu2TBNav+0gdI2lZGM618szgAxP/Q06wDJmKOpqkN9bU/GjjcRh
Lk2s95tCwFjmt87dLNg3MmMTGF+c5cm2J0Q3MnIe0ywMyLrTTUiOoWf7E6haV/O1Q2aQJ89Mrhl+
pcV3LjqgmPdRHngcbBV1LU+8lVlrQWZ6xPb95BuDWcmP/En3yirHQOXpaO8HoVud83E8CN/PLGI1
1kNMd0JvApgp6og1/HM14i8le9XyVCvP1QBNleyPBf+u34haNxwJ4ljikPS8k2J3t8KXghrpo/ra
vkXz67KYVB68T4NnkYwWJhb8+9B1mT7eQoPDA5HAxRgzdJtFUE4g/1whpd+B5auh2nY2OYnVYP+H
5gIFVv4OkyWEMGktZ4Q6KFO8Uv/Fpbg/DrLzabAT1uIWvEaYuMZbUfiFWKNFKLqS17a9oE7/n/Cy
Lqk8ZD6uDXl2mVAXejvka5gFpNUwuUIJIBoHdryOkSbxh5jK01rRDdyjcmDeXcwXV/HT3XowRYOW
SQ3LRK3Hb9JyffqpHEThUDi45InOI9IbMU9cYk69NvhRcInLeLIkmdqNQ0CPWpDXsDv5r+A6sRKR
gwpf0uBuWCEkEDOkf0TQnd4CfHqHBQlYYllvxaCC/2jno/DjHQ/CGJeNcv8a1u5oMHJDrqUmZO8f
bBYFO3KqYYxDevfXMP0Eo14LnAhRrtVs+9MeAF5GksEkudgUzu7U5OgvQnfor9y737hBSQpA8g8O
xe2TIBwTayezxxzy3TPwBPtL/2F1eTfEr8j9Do8ZrbOXF86kytvAESnraHEwrvDI9aNXRbkV1rHZ
ACGO3Mf9DqEcMHq2lmO3bEQeLNZEjZrdebVGLQ/Rg5QCgoyOeDK5nfpYOLSMR3GoOHR0kwMDHHJD
Oc5131bcTyML8lnhZv/6oJPMISSLB+iZMCSgdNSgIaYYn1q5dncxbc2+pBv2Dbp75FnntPAs8oH6
ruo1BDT1EsSG4hLfaVcusd/XQWWzpyJD+c1FHW1iRI2++w/mp7DftOH81+5516Wb2zqrn+02xkDK
S7dr7FPY4029WcLVh1SFasiGvsP7b8/OAbDEBZKkCYVx0PUzF+yCpatXLFAy5ANaslFXTzXUZEmm
3OYAQ+AoufbPL09RBh9imJGJ0ygIxSYBnE0raG786gbVxO352nhTGANxWn9ejMxWNBLawGCUxukf
D09KcLTto6yv2ejO2s7jts5qYNGOgBuYFzxlKJIn7ZD3ahixycL3IOMrWJ3m9qNUfynV0qFM4Ffc
ZgJm8IEO8+8WRiUhMdBEvlywVVhrZ4/NCqRmJKdm5AGKJbxui8hrtCHH2T3nN52iyxj4YteILERr
9Ja1ircZ9Ek7Up7ujteUe0u+mbJjj+MAuCwTiiMJ33E9HYOYiRrhdrLM5KIe1ct4OViPXNAwCx5J
ecZjqucwpH8ARka5mn7n3Ds1zgxhrw3qHs8fq8f9oWCoGkqROv3n/V7Gek4QsXn/D0Mc+VNx4bv2
3ybQTd5i2HCBgX8Km1/r/0h8Oh2eFLG50VkY3Uh60WxovGhrwim2P3I7SuzEuBJuUcEeRmeaqrPo
fRtT1w53o7AblobgkvsYuw5nNjoarjG+aYkUVCaTHrSK0IvSW43YM4M3mXK+WRLKDBDpfQ73ER/Y
+MMM4d4V5eVSaGr7d37MnPXfIRY0VkpwWO0cDFQ/6fUjW256ykIbgZ4da+WaemuI9d7ufmAgowdz
4Ac9AatINaBvO3yMEEp/VDAFQG90o1My1QS+pWrdrhri907hl/1DcyKHjL1mveipT8sViJBu/baM
X9ngpkfIzR3qbwRyn7Wd4Ug9E2hT7pKn25QIc8GZ/BS7rlVr41C99ORHmqbyr8G8MJnR/SZws72V
f6pFwEmu5p+/Wf/nTRqhhNxWLS7dZGKh+jYYNpic/QGd8uRXMHLHeSU++MCN2jgMBEqUXD7CeV3k
x+lGALdoyVPiahUsi73PfSG8/v0mSY+2F6rS2yrdSqLuvYRVF5zRo0q5JrY0lvOb8FS0ZDAK6Jcj
Gyxzn+KP01o0ExGW8IJPYYR51Jg5o5efD1cXdFb21oXd+DeeopYBrxS9i3rkIUBFUUe1j0FUGEsK
Eol9Tuxj9AXvZvrufX3QKoiUpVs3rCRkNkZDQYggp5O/ndtJ/qeImZcH0kRAnYUKHpBZ7gn9rlL/
Upl2v0iKep8RzaVgy/v/mzxAw9/y0SnVXzS4WPh/5/Oiq9CwMWZFR7yMIrWBZngLrAEOsAhsrYOw
zsHOh6ww9R94JC3Q4pT1U2DFYWxLqmcIAA0YDz95xNazgVV2YVQQQkUbIbMEmoSUITUuT9EQyJzO
LBkuEgNt4fjb66l0k0qAvXrlUoAXNRyUMP8pR6q82TRVchRsu2rl56qsfYNDeg5azrDFsgZF+lj8
uXfSMwJytb8HS+AeQW60LKdqgMrYDKA4opbz7hvZcIQYOiRrC9RveaSG5k/fg06px8jhk0DZlQil
pKSmSdeWLA8SuEuDjOh+RHgePva82c219bBv6YRYsR/rjskEfELKvdEjEMJ0LxQAGMPA4jz87hmB
f7qsd0tzB3HpRIu2a1+A/UhVTZeHrl/r0EYCejyKvDP28soxSBo6s1CFyOfhiT3NdMvDGO91Injb
04eZFxuTg5g6vPCk7L1Jp0/YtFrPpstBzpFmulnLpy4Orgsi7tWRgy60kkTqIH2d9gGpoLE1iSmD
9guttlhs0jq9VYpJt0hSXmVMaMjf6idT/vgYQ+Mm8TRQW+8QnI3inZASxc3qOfh9uPWh8PNF1BjI
GhrXVqa3gxEHJkeFCO3uWP+1Zq0lLJk4pE4EUiOXeczozwztZpEoyOcQKnar0IPx/g4rgSck9Z6g
hoFAgCfe3WmzTyp0RgnkgIGN0krW62BAatMAVTJddS3osmRIIwoXNS+UrsRkZYGsWqSHDQzhKOan
UplbebAI2WV3oGP2c+LeeGqB6Tmf9dD+WhuWNXd5aMeSaIyL1ylysFFSC02fk2O7N9a3S79wUk37
Ui8T10FoSBrPOBu41+hLcDkZfZr5jEDOXmgtwPXW/GDs/VY+SZToyQbtFUyy0fHW25h2cxxURAK5
11/Ie7RuVNqSGE/uGkeUGCBCQo+NwG8Bu3eHeSmiqq5N3PE4G/sCHUDfnlVtTgLcee1j1vT0QElI
AnWOY4fFU78XacilVgAsmXM2q1TeWpnVY9qMUIMftIh67sbveOVP6OBSM48EB7nrX0Pr3ziqzyUE
zpPGVb2gFDP9d/Kc/+V96bB+Ga8eHinAS2qPxIpoX+WVgNHNt2EnrqWcKG4eoao4eazAGW0epg2j
NvOgGuVlol1cuRzIBSK/VwfYTwiXWlj2YsJNdnMu1mR8bVsmp/6u8icPZAMwEHJkfVf+fp+RaFRz
i8YG3oa/sg2d/IykZzDFwE1YmAAYZbp/Y6EmNwuA/RBZLSK2+PPvQojnG/bLRy0cdezs0yD4mDFV
iknUOFiLTdEwsoCELRDA6rTisD09GDu1COlNJHGwpO+fLqCbYF27FDPnjmcw03AquSoi6n0FT/DZ
T5XE+mgMFToInt1Bjvo2u7+ToHsp15Q/CZkWaohq1A0CqbfcObD9KAkN+pTx65kB+/PyyFXxQZ91
TfqPoxGn/dHFm07BMlsxLSKSDsgsvc74PM8ycGkGPul15XSd/ElRfjIWpRS3GUraC/eYWdaqqlO4
ZF1iLgJl2YLhLqu1aKvMsqNIveMm/ckc5cj30FA2dxCnZjfXI/+ZZ3qSkipDsyPG5gX4uLzVuwUL
Hph9WEkJ/BH39nHURQFfP8z+c+OT8mRnrzU0m4fH+yY/uWXUmMXlFaMaH0cW232+KbNYDLt6IbPO
7mLpJyXvVQzV+XhDXDl1Ytp5IkqkxManh/RsGsN41eyC8yI+O5oWXzYvkW6CcZtO10fffQ80xi2u
zRk/xeJ3rF+FNwGWEKPetkxaREj3lSiLwPwodXcox2FARbIdlk0l4xUBXvB4iC9CH9S0Lf40LxQ8
B9G3CklToKFV7v3fq20gy8Nqg97c1WVjgh5BpHBlFRGrs3VMIybQg/uL0xXncNy0QbCJkpceWNBc
dlUOogsaXWlCAEBKwiLgIxsqln4bjsQqdo1AVWyx0JH+H6bNjh/ge448GQVbyeX+r4yDgu/stKH0
cO4G8zOy5AxiivoUkyOoojlZsUhl4RftKU8tcT7PCgMLPAeoWzFxZY5q9q6hkvwHkd/gUQpRKUvp
SP3sGEUOhI/bb/muruDx+OMqmSJorjEHDrmfEgcVW5ZwDyIPEp+2KK/9eauSN5V4E0ACedV2pXBo
XDTfQNk7iPyfbrSYZ0EJUDe5IfNFVZsTRWUt8DTnVARoPdUFfT5X2NT8CmtIrQCql5vu7kR3DMWw
IQ4sjNwNA2G8C2ZRfB3B1jgyFEfyFe2GuAFsCXwjVEQE2dfZYhLdg20jZAPb/a8Gu8cFp0qDVWDg
zL083R0ZMtUKUDIAkfwEDp48yqDkPP7utzFr0yNQzwVtQorzPkjTdv0Q/E6gT2UXQWZ/MkQ5PcXk
XD23IWPpYjSdxn6Uuf3SBvdINA9AXOke1zD2SeBzGLZTbUlAiKAOoD7Z40db74j5Ndn7/qYiiM23
wPWH/wKdR2PfvoHv+f+9juiRce1j/esWgW7xz3jlqnqFgjftjp6aF1QlMnFMpnvNBR7oQQMwAEAL
nyZzMBXEi4lvbCH3Tts1JfhZmdavjusWSn/r1ThoILYPNVTMtexbDrNp+AritJV/y83xmHTwTByP
4QNwlmI6mgcu4I34ms9z3JYe/Yb5/YW+/GvB3wyw3WRhYFDwadaPrfybkPuqHG30uuCyTpZopXdY
3qPETqFkzQRpfiKxUYdzo5VbiOEJYgTaUq+MN6qkPICWxkVA0JXhzH7at/uOyggtDjcR6yi8vMlp
l1sBLULsn39JtmHkjcT0btRSQaOsYWVzIo0v9+xnEyQnzNLRDjkrNbuwE+myC6Z+LZ7yG595vSua
XEI5Q9tkAwTbGmG09+DYhViN6tJ9DDHlzXYn83O9ieFQaL1/BK7/U3Ei3+tKxGW7Gn6z2kmCze6n
DIuwcSvnFL9YBxAkGZaBblyEAd9iBFBraDIihg0Cv7x+nY2t/+e5kh8csI8oq8cjkxahaj5gFkUb
NqwG07xDq5WDsKusyjVyBE5LItE5qJ/ZlF8LSteKfF1pO1JfVvHbeTvGEu//F9fwPyAyDxTpzcUt
D5uOP79RTMU922JWFVA1fc4u+Wkqe/69QZDYUhajop0MlIujR6vUXEuJuhGpBPSOq4zegUVpeQdZ
pPidf+sveBIlZm94dQwIH56P7KZ2bbBsVpPjWoLwYJbnzod5nUFUM1akUpJJZi9Tc/1C3uTPWHV2
5yLLZV61WT0EDwOyiVFaGidlKDcksaSTqKMPFmsFKG5Ygyv5TyBBngo6KqYgbLg/sIykmKxG5DL+
N60Ji10uXEL7UW8yC3R0FMumPzVzgznQXMi7P95GoesAN8BgNiAkpR1dgnbK5os33DxP0qkCN6iN
EdEVnYHRRWz/6mHRmI1VbCF6tQiS77nPXkTZE8saadmb76HIMd3tSpBj9K6RHnuEdklnq0zzHagB
smf6ajz/+6cVn/zr0TMUmXTqm+TD6pVsBHCHvPoWKWSNIOOTYWHorWxdoAaCu6FvCOJsdthxCK03
K8p/gdvWkTBkNnRB3ASnpJwP7JuRsjrqBghqO7VFDwATjEjZZB+V32T+pvoslwINhmBOit+wEkwU
h6sQ58Ps5ieqZE0ERHUxTwSNzv7ya1gUxXhJdI1WZWPhyohi+mMRjCn1cC+AdgBv8mWe9s4aV9BM
t+NU5L3Xv0pdvgC9wuuM1MsvxT2azFhRezv3VX+TPkxTiKh0yCJ3r8m0FIHpZzzpM7U1kTiKA2hL
q83SnAb9UDRwSVtNuidrKCj7dxyXeyGknvusB5X1gQvbsI3JRFvyjbizJFHKo6DBFUHtcX2lABQU
xDtouORc4iqjspKIHgjr9QxFxRMZnjMF8o9ACKLpKXpSL3n2hRJUNzR5Hh4PNBI6MPLon+fL6Fob
HPLQ+9CN23ZG7TTNy19HHeaQMo3+7XT5h+KFQ1RfapEts+WAsr+1kw9lyzPbBHNwpfYM4lLmy+98
FVGKYibZ3FOqXQCWA2Fq3j0DxnYvxvehnbDN1riqZa8iM0+wtWyD1ia0VrF7CfRR4K3Yr5jUBjlE
z51rB3vvgoqv6NApEVxT1Ae+oSiV6yxSMIN2aIXbhqDaI7wmMC6sXbboGLWNbpjOFUI/S34cwedA
Pr0oJYYjHIRiG/r+eGwPOY+XPhCOxxPI/PFnfVyS1jjW1MIIZBwYMc+M9deWx5WwfSu2e3e91SdQ
f4qTAb5R5IP0EvSfYhpNquvz/FDD2JzwRQ7ArvAxqBtX66KZPSo9FTB9+S6VD+qqQ5z+MwaTc2yv
mQcc7Y6Jn/PvoKIrttVHZ+kF+tqxswxz0rqJSoXFVQ9CQ6jxQ2OBAqA/O1ICOpoL2z8PTVpirKrC
mvGCMAMwz8ea3HsMRZwuVSIcVVC4cJ1lv58NEtLP/ObWLO0y+PewTWcJSd/9yUyKM4oa7CLynrOD
OU7zUJhY4RY/0+GMcLMBwhw8hdIXyNaSkhobzZqzwAlnmq6FGemvQzbmtSG7y6FwVnuuLzcbodwj
zvzcum9KUPb7I6ATtuLS3+gjQ78VDgpbI44V0fLoMKavyT0aLPpeddsUUlT9535W6H6e38GBGuXW
TxHddxWrf9SXSAScjYGGheQl1QjJ6xP+SMlEIjGFzZ8RGm8KqXtgoxIZ03sNUL4hDt2LVWkDExvh
FM4SuSlqfKGrbrdntb0l2Dj7Of/LjZJ5L8r2TP3EUoVrW/in12NHNShPbAt7y9AYMxbWomC6J+AL
OO/YbP38ShsXqWmCizpYjcxnA3DbOj+TepP1K4o4fUomdBXllKKgyJyRpKjskamjuw642URJhSwN
hnOIXkn0PnPrA356o3sqi4RnS+ypcjleQzRsl8jT+K1cGgZbiFTLXhIdQffhlbq9rdCX7jL5ANAA
LgLhMQ+ftd5+gVzGcds1zINtBpBADvwQlfTTpzw2O9titG1Qpt4GZt663AIxZgEJ7HDZgNfzk4Iq
f5Za05RzlH0G15bl8RMjYl7HeilptD3gdctUAuhdIRiBDzNqer9PQ5Ous5kYDZDhLRvYpTw5CiIm
Dpj/umtHwOQACdAGVqT8VoIC9Fb0q+ogq2YPbWEwdMXH+/KL4s6/z5nF535h1/Vm5k4qM7S74x4Y
YMM+mxMw8zhAjgCPuXu3AfgBc65qW+viPcnOTsoEFO25PXgKbOUbv47GPzyeQmDPN0tSon+X+m13
iehakwdLRXl8cjJdlC5/yL/YVPfC7Vs7ZQUrcEGf6DpzLKdj1439n4luSnUOmoUf9tZEWsef7AbX
fqzgO2p0LADbq+Dy5EXGFb+yHUMkbwY3d9qw0Z+kYuYhjXp6zt7cXzsR7RcZhugFvrCvbskZ8jAP
sYGjHhzRADbxzDBABwGmggLZc+JMFkaKH86VBu1It684rjWESbnGeIdN7NPgyL+E1G72glsHHlLz
+09z2Ws2nOiQJkRUBNXjTs7EpK1i5bhGjjAqffjgtuHtrv3gF5xJM4qoUcjYskIGOVFXY7A/X++2
IRDn4YtWILDkVwUt5qgFKliggamqNaWXVyTV5ANrnyiJrPk5ABdQhiGpWOYb+2NVEztjvZVuQ4Ff
D0Bm6Rly89n1b58sY9ovNyxuiQay66AtShAzXZaPJaXARpbnd6TENZ9vj69G2qEMymvDPIsm7l5C
MRTpBXM1DgurJRZ01cMji4NqMcsSR99ZV8wbOtG05OZPnrF/MikQVJPOnmrK2w9gKqBJhkC66kuc
BB7T+sT0bIZqi3mXS/vaADgbGZNv47lzvEHoOahYNEpYfQIqpKJFGk4ANzDYH5OR2dewd5W1sTu7
HS5Z+y/2HQm4UboK9Kba8rFgFuV3Pg1IOjdvXhB04jDPCOj/NQeG99Ae+t7ft1ykzO6PgwFB/GcB
5leOx12PQwRe2OLMTmJH8y5A7n6uCtOv+IAU/Xv2+NvNhX33utghkLCSzsEv8Y9ZnNVuRbLo+Nx7
HJWaM6es67gwwVj4e5a/twFxdWy3CraBwG67h4Z6SAtXHYHgH7e6pOZCAdx04v23zc6h85f/Zu3x
AxnPTa3gzsq7oX/wcXv94PYql7MffPGXo5ZxIRXmVVKNN8hzbbltIK9ein+SlxtpnBjZ5PGRs9dz
Hk4fFBMtKYSza511kp1OqTm7+rbEbDXi4L9afEl5MrQxKg/4thYgs2LzFanb8vPvcarLalDwH8P0
/ZE6s1hw4SvrSqD9DEXqGRUl02/vCtYBhh/12KjbfBBQJDcGNoRq4AgOYNItU4dOnERH42TKV0yF
IlXSd/MUN2NnNiZ21omMZmcmP+3Wu1pKOgvcC5vkm12cI7hKrOiEF5LoMeEB7I/AdsI4u2OKqoy3
BkIKSb3mMCV6xdSkhKqd/n6BFeFZC9X803bNGUdTxWp4OwdG1Qg/aJGHNfLByYR3D543etoBPXme
V2MqWt+KPrkZjRhrz3bLWNGxJr/D7rHJ+qe66B3n951oTVBv43vWVziVW49GU2eDYc3Zuwv1F8Xu
/gEvokLgfjM9pQJ9Po1niwacfE6dFRxgITpvm+9DLaKAF3v+HHeuZo4OF66cTBh6iYB4g8DRsB3K
8rYsndDKdWaRo/wwfRfi2V6SwRJnnCymDmAfAbURRf5KQO/PV8BbuIzbsDVSuK22PMJ7E+94JFxL
uOY8uP23L4Gt1ENUckXqOweYvSqeChFe26EAw7Pp1mIiqiCqZBwVr3IQX2oXibIWcQGgWrSEKVHE
6q2N0qGBhW2FcyYqKlXiu2K4a6ke6HYoumJtiV3e6TFAzhm7SxIkBaJUT9/xnqGI240zQqiLxVcC
MLt4KPzatuKFetenORRcynqD3ik1nyAZI2tukxe10WW6Zi3VhQ/l4T+8RYF8TcnYSsbLsvQZNtQd
YKqTbSwdWeohHIcKg5ra2P+ANg98jnzbc2oYJe3gu/OEICIhRra4ZxRJUuVQlmNQ4Y3KbIkiMU0n
1b6MGilOhtK9GhhYJwkqIxNV9KlKuTS7EU60TPVfXa4L+OTHE4YRnEkGPZe6jVnYFuSrSjtBQrMZ
8mtA4w2Id61V95eDhRQEtlxOM4z4KbvtjMyiuHnoh+sFlTXW7gV3kUEBhpHfPlX43+9Tylxsb037
CQXs2ukX9nQnMzAWS37uNHySdvPxOdsMAJbafnfHv+Ka9JFkiyGzRw8T86i4FSjoZsR75ayfF3Qj
bTfpSIOyJGrx6thNZDxxkph0xu7CGVWOVREIEAjpuqQtgGdwMAPoVbze95yd1WOPB1m5CylpwkG+
QPWPQ+PPq6/NOmbXCGrqWBJ0O1XvuF66LuVZvEO44/hNCeoc3Xvrg2zWC1Kysf4J78bgwQ8Zi4e2
cO2+pXLNxwg0gIs7gWoveuK8hRaMzayjeCrvnyUm0k5hoI0R0updlzcQu6EihlT9N8+xLsG1afHX
gBd6g/13xzliKTLzTIiOSPhObVn+9VpfK5PwKgPJf5XRRdFSbQpJGN4Iam2E0hNF47af90qBiGC4
iIPJ8s2iLa99nnQNvOtwwlD6Hz6tCS6xCXhrtm5t2VGKK3SAMcbJ+03k4jX7tncx+9ZVhMJNjKyE
t1WJ31qCGOdwpRQLTaVOyVPC4evzX0fvkPPZT9cHaTGnt2q/knk9R1E9LOfoB42wWn/8DC09Js3d
eAIAmHgUcS2ILvGxBijiddJoDfQjKWNgqoPknE01gHz4T54/BWk6t3y4dgxIMyP+t8Iniyh//v24
G8SS+1S+sNj/krRf32vyMdz4xY5bpruWj9v6d4xbrkNm/CqPCAXVHBq0O0+7C43h+eHCPJ5zvCiT
hIH40QS0iDfoYITIGH6ap9/qNG1zgpZgjdrci+QcDaS879oySVG0eGhRxb8CILQWEox9Gh8pLE2i
ul6f6hRZ5Z/8q/XraHFGYwupfJAPYmCLxbiMVhwgV/F/p7nWxYinvzob0DXmnJEWccjx+Q3zwgYt
PdSX6LMN9u+PiXoW23OtAS6MrvHm462rM8ylW+ZoOjdYXrUkG4IRr2pVUoGdCe+dDiTRHNI+9z+U
k+SrSgW6Kh44aP2ImNl91RUVhaYT+MpjYMrGUv/ifDmAGrQWTREb5+oFLJJjePF0weqXWqQO1CDM
teKwkQCTOnUGrNsMW07JkEvZ2NFSbJDOpzjlmyHc9Zw1hkgHxM3DWyZiIY73IipOYJJjGEAaFfe1
9zuLT4ZGcwQN23N87yQ1MwhlMPIzQ4xOBi6tD4HHqnpVWZYFyjkrygvSgp6XesBa08XOzuQxGzxN
92nTSRggB0oFOFhLLjpoOGWmUhELj8MNxcT56nsGdwGIzj+fs7l7iYVx6sruzbzCeB5TZualPosm
b5EmXPQx1ddXtxOcI4aWJBwkxJKTZw3ztmFNKHe7sEmGUI9xqY+3Kzn/DNGO7MZ5M+Ysjr2ULSOq
xAQ3Fc9v3EcpKQ1w8t/EpboqrvmmhBxaEmyiXZaWoQZtMTytKeK46inOEUEsXJNk4hqVYN8j9foV
ecr6lOs+qyaSYJ7bbIkLsEauKAsjIfy8ie7y87ZVr0ipDXqtY9u1kLNN9wd8PHDBBZwJAF8swUPL
sBZ66zNA4/H+891Wmskuw7kvEDfxpRhwud1PYmgoQQRhlCzqPLt7SwxwYZGZz4Ojvu8+rHdNjh96
CcWJe8EEs+USFPWBfFh3lh8hK5YCgDYGUVyBECrwy8/K2RGXFiZ5cHtnLtdaya4j2FEYn3qQ4Ytn
k1aBzhDFSIM2X4cq7vw3JWCk+ecElMgQkJbepTnAhqafP9P7H/9Im1lY59VRqfq6rdsuTkxBu9CV
aQc1WAkRQUJQBHKLYGxbWd1feqeeYKQqfq5L9qF2VDuVHykXRWYxu4iUfILBrdku2reGyc4JNw83
M3DHjIlXvE5ODqFpJhTyFbWEgv+f9WQWCFKypeRzQgtOV06KgzUQqu932WhgatWdIAsFodZET0E8
HmAtUTCGC/EVvznKnXMFli8BrC5Rwgcud7xhqiwKXLsjCWidFG9TmCX5gDzhTzLcnFkAT2TGRAcr
Yh+L3Mays6eZLIJcC/3QTbJL9LguwldmuZR51b/vT3vrTBL6Cdvy3nZGCUZ40Y2RHMYZBHsUOyuF
2mteRQAZB09iBMmFxe9A6K/YdWBoETql9jOAPE4tICdTpBV0RRCDU17uRJxtduGmIzlECS5KP9Kw
gWcdOnzrjrv5Snr8Rtaoe/9Drc6I5KUs/crb87S2Hr3U0lmw9qtzn0ZfKsBnuAGwsfgjhhfMwZ/p
XgRmnjWTTezECmTbVzjtnZixdsDjOopBUUtUH+doFxANPwvpBbrh7gEX4qukj2BldVklW/iw8h1M
og0T5G06xVgKkImHYcHEvoC6ndHCsmyeeL0sJLZFIlmDPugF/S1m1qPaZhVwY8sqBjJN87mdP9mi
F6G321Xo8zTVk0fWNp/N8IFV0ug8321gQr7Qzn6LBQo2iqNYgjdEyMs0IDtZPPx9jsqs1UhsVt7u
B1n985ahOTx/CFP42fR3+fPpPHTM5r8bubs5egvLOHe/Naq0JsqVVnb6JjyYwXZkdfXJiW934EIC
i3ZYty371BQ8TqI9WpUIIL7/clJXr4cVqd05j6fxVa75WQDjMurHfnVAoi/dXikwvZErtPatddLY
njDrgj9aiy+9Zkqew94aKSGNPjb1K00XNgYZQsH4a3GolnEjOdI7XJVWoCGpyGWj3wWlDbQyPDzS
Kf50FlCgyPnKB+pnXO4rOPwaCk17XP6qP0radVKsQdHD3H3flI8LhG6R7bm0eJqNxHeqmG+8jrj1
qJhspoPLWt9nNSxlsYFmCr4JDW9Eh/9ZyAVXkCjPapR/Tb4kTHwAC8EWbntPjeyzpwcTL+abMgMN
xtrpWU3XDJ17qBf1H38eJlmWt8VxpWcUeg1KcoyWOBflGOgnamjBNiKg67C/l6AnZ3OuuevlVCXQ
aebiCx6qjh8P7ToII2XCPJ2O5/cQmN026X38cvowGToKuW0ZECMYiiI9OGiovbmkgYyJWcM4ogpH
Z1vta1FpYnktAMVkARaKF5mQ/XlY97unch97U0KifVNKqQ6+YxhsB87dmOIaUSy6b6G0RPBy61Sk
7+7Xwwmcjpa0F18xX17sa8HQggrfkvGYnLdNdE9qXwUyXB/OzB6obKovebL813cMG0gtPpSmgIDO
8hPBLIH0WlVn/8JuaSwNGQZYeF6YhNBYnBCl4uppueBTgu2IwlckCiFPzWVqDeyp+b9PY38K12+F
Ey+ysRiIgmk4XVIaFDSbkUByIRod075G0Mj+WZkvwZbMk1wnNsknXKE2iGwyDPifyiK7aJFMzD4X
jyMpdxxPaOWLceMxQaUjG0UANyueu7GQHxv/sy2XY1ii0XDbe0U9qtFC3PjmfW+iN4/GGcGpZ8On
dx3W+IGkDiij2/EonYxKFkvFJECcsfpEXKDaZQWdvyz3sd8uHRjiL3W/l0S64ms6dcic2yZ9P9e/
N3X48VAB8fBxNYwx7s8VFepY6+RsbGTbU3zlAfSOTjGya6hX1SGoWfYpm05BNkpS3I+v/REJdvPZ
lBrCtXUg9gd6l9XWS++/sSURq138xbRf9+20gokIrQol4fB69ICFOiaCfdyAiMiZAdolNpIE2zf5
WTlgdSKC94NDcsrWTkb+odMea+EhtQAgm9ztUbJMmkM5urwVSfG9ljxPhXTaAwbHk3ExDA6cqZg9
wtmfnZMZHZ/q7jY/chSSSHIm/5Sby9S2IofC01FX5TuKCa+xsDD5pWjDJYc/v/vnO+vPu5U4iCfp
p8zVqO6cAal0gO1CcUMJ83LYd2uA2Isg7nIZsHrxdZME0CKfsIQtq+DG2jsX2IsatmCwcnlqo8J0
uoRJYj6KXI1DkAw0H3hxTPyb+A47TkA+zEAnkiHXADuq52xwwemUSd4d48j9RZIIzQHYD+5K+3vI
BP4aNtEBmpHIhTKi7ekm82U3m7+BOAt4ZdXAzwGDslonButh8mjqkg6IM23tCpFifafjAevr2qS0
bsYUKDrdhumOGgeiLiI+gDcoLMz3wLjAEhXYz9TOTAqLuOjKHRkT0LPb3Ow2VJ7DaaoRU3lF/OJL
FeiGcid2zRvzGjYp54DatxIT/8vNWffX2cS7U5VKlr2qTcG+tff/H/E6GeZ8Z1T2yzgrR9wAaNFQ
lbmK9Bx+VFqP76ZraotVJTQ9MYuCDTQ2DqYXSC3GRIrVnHVEoBP/xIvr7Bf30lOgIYWKFd8UXDS1
4sg2XQTYFt204Qx5L1AxhJnX95GyZlztqlHFtuDSpE2R+0s73wmprCSdbeRsB7G3mch0r0RtFUSb
EXNhTNaqAn31hV96Ha3xjpx/4R5/3ucP7GyuDVPZoz9gHSQuxCKcX8kgk0E9av3e2vsAphYKsihH
Hc8lRoOuRKmZ+csm4Yb3XvgV8kXnYBWhB1a6WU/N/C4zgfF8HBYhi6KFv6T34/Vz8MmWD40oerKA
RCGU9omEi6olLoB3+EXhcjRGEkk1iuFgl/a5muSbn7yCT1K8dyNykNb5c2DkKa8M0rMjnYsYd7oh
fteemI0XW+bsdajtvn61riGqvqH9zPdjdUC+Uv2OEgp+Uciqm4OP81RVbf/uSF2YNc4xXJ2MNo9p
QXRrRI6VMjL9fkRYvsgjLh7SR/JswoD9dlTWqu8SGBBCkoJW7zdTmoIFIahlDKAn63AT6iIfqNgs
TwI61RaA024zdKASUYlIS2OR14xYYhh43X/XxTbQXIdx12nsS1xy4RodtiVfV68UxH/YZdLlkLvv
xhB2sFZpFOrr767P6+VCm4cuUiY1AH1PCRsAuyQslxwm3VlelxelB0E9572w2jmsPOqmX1oao1Ca
cg1NhoYD8pnO3dV51RShpDfBshi/uqRapRvadHdI1sXOSoCePq762QDnrV9RY+pXFILTQkdBVaJO
kn0pME0cebEcM+2yYNak9p1BvQ6BVpJAJqZlpS6Mn6x1C6rShldJQwltAokFRJwdXMH4bON0t4ts
P7r60wQ8wMdtuCnNfbBidv0iFs3jBb2us7a8+yqlXzUP+ryVaQ4Qw7l39ydt2l7cuBzVlwhJrv54
RfwhS6RkSM/QOWsf+1X2GELuSy5s2PFrSnZrfzJun2biQFF31sa1h50/qKZHYLShBpcYiYvt3G8q
MT9ALhuE6p9zMyA5G1PX4n0O1a2z0Iy+l2v7vGt7VxkMF6iH2nqEBCuvAfd8NVQAs1R1XlRRBSad
fM2rkCXhE1gwrV99zkFJq1YETqx+MjTEnQ+G17Rl3EEGNyy85s8BBQOk+Vjydtm//RjlzPlIDPFr
tfOOtDEe+7o41ITKaoADn17V0MCMqYRPYawjeDbGnhVjGpck1aemFEXr+B5nixpbB0x2X8GnYdtv
Rwjay32wG07dhA13Eug1k65kegGo52pfsStP9p/PG49M/8tt86D3iEqKw0qKb6j1NnRSxgsLH8vY
4T6POiMshwGxwIqRDdsacNPa2/tMnED1sEpgl9oMDtdlz0zK6q37RbBy2aUm2EUzjYNDDE8rjIxP
C1tYcI43G8SdcyM0yD/ODA0NGyqdknwIL2NQYsunxSXqZXCVyIfWgvE8YQDgYZPlPiMpZy6aiXls
fthMepUQcGGfV+xyctOU+cwatAKiAgR0adS1wTdoEjLdm/rRU7ZDF83myllyCv39DkIHZgfJ5RnE
XgOPhpnNIsSnVKAnjMWRGKYzL6BKSuHSqIeCrnb9CadTjf8EZ4kGMxKqENTa3mRmIkGl8jQ3lvzY
JXJl5YU98hL5x5uDQMLk0YIoWeAQINDbQCIK9cPwfd8++Qtz8vYTO2cosEMxT+4T0+du8dvbkJ9T
UoAFOslmX0uoJYPddPDc1eJx6O6PrjtbrVbTPGzSARx7ljILvSMJRSohzuOwW5tLpmKbM9flQxUO
MHuh+EM5ERR9NSw1hkNsBYT8wGa+DcZUAk5oZvn6mcEN7WgMQvLimbVTOKxJT9ZTq9LZ3NPYaMFv
fkTE3nwhL5KEtONv6vPdRGwRVkMyxqlekIj9nE8a/w/6/BX9uy9UHJ0m2vMTgIMOuE32fokf/AuR
9Qpy1p1xovPNBQzx7ggJqr2bUPyWByqq/QvfBV/vfWSUMSdd7gl3Eyljw6LhIoEE3LOD8Z2IMYCs
LKDUpaT9Yczkl2E5qr7PS2hE4EFNReTxndBPbDtilib95PqydcH2BO+GR3mO/YYYKEbiFb/ePpfG
ierb7nApcj1eresukQga0Br7WaKl78fmLSmL9jwlEf3EFeWD5ukulAtNN4RNQR1vdhTj+2OoTred
wVECVaC6SAMSjjpaNIwflvUHSVjqRldSAZV+HRh42GV4oYekvXKvStfeXvRKlYjDSgy6s8JG0q/l
UtV5MRIchNNIcHC/fg5qfsQCmzTohWWHhrQClyrLiMvABlVw/xD+uyv7FcpPAlAGf5cRckIMsGi6
JLDRSYWNGyy589IOMheQzY9U+XnPPXXSf5XSopCwLNr5XUnPwerCwNqb3aIffHiwbP/9jHgqBtjk
QINan27FT7epdf1ZW1TOqx8p3S0DXEZyXdksdkk323Nnk2k1AyDFjISUcjkN9eCqOwv5GphMNNvn
zYAfnniSCFzTH90mxRRH6SYol1/SbiA+UBLIvGichof1GTYdsN58dc8mo0aEI16/jSwsFBoG2+0t
r8cuoAXS6yu0d27Q3BHxqTXl9YBWU2WPgdViLkJchlFtAo1IjRuN9Nerq+0RjMHIEEthMsSEWVkp
vQov7J5NcRC6bPpTgU8TfaYcNH+WDl825ariYdoyTzFQjJi79jT9Vt+EKSM7sjERWC4ODjYDzVH0
atHq5qOLlRHODx8SKZovDVSW5Lh8xRzP3JW2zhSgyivv2QHf0WBULxzbEYdPqMY32aC1WSAYreCI
Z9SE/ZBG4v+pgf9NATM/DCVyEBoXEwEpSftiJz8gzp8l90KQmrSd5I9Drez19LA6o9Z0B2nVrDw6
WrinFODFeBx/AFUe/hgCRg4UcQoh1+1xTr8US5ji+PRXSwuWKHk4tJjGyncDogQiKhezX/ivXYNe
EJtIZdBRqJ3tsnVLaE3RPGbwb1F4tKMQU6gKT7TtxAhOPadI2gdFzCDExO0SukJkqIPIgLpFGXTh
Zc83oKGkCQlD9MK7bpOpTRRmbujluzRpCAI/9ZGo3R4i2MeoiFQ0Zv54D3QrIXvJ8GYANi7JYO+/
+rhS2O3fs8geya+5+Rog/qWuPWqeWt9PWUTu+v+5yHYM7bx/fHDLlUapJ82VWH34c1iv7EGg5cnd
tWHDiwNOuVLE9Ll82T9mSU+DWgkkqnqgxZpTAyr1/ZPftEuvSHupZcAT3JwvbyvCMnX1EP3sgBwm
GgV31j6qSnJB+7gtGGLhXr4+Unqjcc6zf2YA2ON9f+/INUlNtTdESzQ5/ZbCNr3nqouo4947G4aU
qgrVjLRXdBhIjlC+hnYJEJOwDVM1T7LbrjBBwvJ2eneKFkWnWkaym0VjOIaEnmk5Q+EsYZJn1dMb
RSxelJXKp3YHKBfsQJ2i5yHC428NppjC4trJPSnydbw1ybamd3X9H2L2n5rgAoCHy7IcgOswj4Mx
ghj3Mk/ZPSj8u+SstOSXlXtEfotnh9ahTuGu8bhnIx8ovH2vzdQNFS4zBri26Ze0nW8ZV1mjluo2
NbrG+O+brrdmAiLFQj94cF+lSnbzTfDn92qgw+Mk/rFsIqRFxNRxIYkcahZs6BSeUktd1dOYh8Sj
CqcyzEYjERhmSi4wmlkOLS77/heA7w9i/D+XTVT9LdxrEjd+AgKgqigjR1og9+fEUL1kh310i9f6
P4Mlr2nel8pe//E0/919i+O31dtYOmSM2pGlpPEciDoGySs+YJ58vj40Rm6EvB9UAWd3Bebq8/it
ZIv/BINwnu9MuTbEueijraUC/Rwh7oxM9AK3VkL2hfP2+Bl+uSJ7jboVHxvcxfXPiMqrF2edTuYB
BuNYroxbitF3XTaz6QBt/2SV/8TeLzuH91o2gaBF27ftlfhz+RDY3qGnlPUmVBxUkHbCAQdKmiUh
6BPyO431+5UlR4T2YPHPq+UK2yDrjBuiC6UloWETVGX7rWD7WGOSOW8uH6C6LMM75WLv5kxLDc41
NVE8UZUsIOzgjg08kCAY2N5zZF360//nER5wjyrT6abzWVSgbSTwPNpOxoXRptoIDq87mbxyHR4h
1SH8APW0C4fKaLG7geDq+IiVDu5/hrKgoR8+R9prH7DKcMx0jcvy7tEO0B3fupyR7foJr+qzrPcR
mo9q8//lwMzJtuA3jp/jK/yb3DVabcUSBWnWqAByPfn3fSNpP27xQLafN4Z7ZLtAbNJbHBCc1rco
yzO7BcAAdYRANPiTym1+PwdrRpjFDWDDEojvbyuwjd/SkkfeFdUrS0dmPfcszNDYQ8ZyJ6sXDlx1
aOvgtaKGFgbIBAuEJbc5MfVLZhVOzzn4V02D7UqZQf2xEWIM0DQkBPkyaoDPGjdBFzhOcoZx4vu7
bQdVd/I05aEfAWccnALdNVAeC2SBInHvWYuijmYWcmAU2YF3V/QGMLlAo10B/Frv2IH89MLkJFMR
tT66FRrjVk3Trw0hVe+sQfEp88FGIwc3nxE+UjMmf596+81di5p3rmRJW7hv/YHhc+tm47aO2G/E
W3X2ZuQCz5m28Du1sNu+qN47/j5aU1MA2cpoybA7f3tF3cWRZGuV6XYQxc2ne0pi7XGuhvHnRMlV
IbkXgoF11bCNvlCqSEGKsCtnDIG0+WB+uS85bmNC+cgCq11bjEAzIssfnWHUfbOj8hK7RSrfUMXD
ybqqgZrZznxZcVb2tPIgN9WZdfk6I7XxWLdARbyuke8IJMMgPP9QwithNnig9V1+1UOgIgCh8Jme
ZKCTQeF2QGX5U6H+Cb9Fl+iEhjaRhGXWCUWwQyKirkfe+tOiKqxpdURCb9KcNuS8uLaIQ2nHs41N
tcrb3EiUiO25c67TjePqBEmgVZ9GkXBID4flRcItw0vFVMvLH6f93HeJNUpxX67F/gsH3vjQAeYq
gndhgp7W5qEElxA8c0MpgaY7B3GU47z3Wl72yiyq5tMTTB1LeO2QcUDRcG/c+qmlz/AgSAyENadZ
hcAG8K1WPLJzJng7+62BAleBO1Xr6A52n+l1oQ5pvjpqisgSnG47Fgf9BsyXO8uPLeHX6yvk0rA0
tYyaz+EF2VTjZB6BtALkZF4iUZde5TqgPU2I9r3pwjUMXKPm+8JbDCqDt/rLhuNQdVPb5Zql4+UB
U804FMcA1KbJoDdAFK97UUqkZ6fJj06QlEE6kq2uF40/MS3L3gDmxIRGR8XowZpp7JRtJXCk4mkc
DMe58X/1gezZWEzJh92piZ1Dh2WcdkoE/Y3bpSD0OLZZsTOzTNWorZfPtE7vE2KrWZCxPfbZZ9EL
yGWefMmu0FN2TITrXE6T0j32TQd63WekEOPt9r1/99MD2uVsrZOuzkiIp/XWz6dB67muob4TXCNp
Rd7ZI/wbOsxq+G1P15FsW8dIF7cFXz7TKZ3Iuv00rcyACBESOojxPojrQel+i3Yk7FHrp+ysS9VT
NoC2Frjxs+zmdJTU5eiYQEziSPi8ruLyBwGWT78ULBfT1pAXGEVusU0fg2HS/FMCs1Jq6vSuXPrj
NirwLogPOcpjl1nvsHD4uQ+vTqCjzcnnIACVTauXM+lf1S1+hfBRu1oj6bcc3DABAmLfP5slWa7d
2LpEc+2LQNAjQMh6p/YFE76mkaGz43iPhemn1Drd7x+AnwbBQePTydhG1TSWSqmDUuXC5b9xc97a
v1mEb3dgF/kq6CWISPTcVwiRsOeKp5P8E7y+sASYK2fFyETlIzrdnZ9ApHlrs89SYb+MusmDKyju
TDFHVa8ZfsjhzThXbVksa2s3xRZkIxh922LYIKtMIySWO08exYa46VZAlvA1GVhP8v49VIPJpd6w
3aDK7pnjpfo32LlBqXrDBePadE2C3WnsmUqy0s6fztbK2+zgG2PcyJ5nPtTUkW4hhMH2NSPEO9cY
/HXdwcYhAJBjPITD5nBmQPrq3VbNLVxkOp5MLKVewvME8fyIX57eY0xARsKJASe2ie532qxOdD4b
PzKF9rlHFtQtGe3IirNs0OstWvqe1KvZPf3A+7mUlQUr1R4ku+tvqGMgb8YAMvM1B5mZJXcW0mD9
QwhxPO1fq8FzYIFInmxH8mR5nIN16E2esF8QOh9h4g1bfzRybcPz9B0EWOGyBBEoAlxVBliwhd36
6/b4shpNK2GivzPb6XHdyI6bvZPi7xxXXxHMxay9YHxS2Zml0vYsdDeD7K6QOBghuHLvkPHJM0Ja
XaxfY6i8f2HihZoCImsBknGkM605xZUGcBIgy0SE4EMm24PC/o7YUUL3Mas5+qrrbhLGLW6eoRKO
te9KrSWKcvaDV1aHJTCdXW2QMDanvVpGyvDHStYwZkNDXXyOg2xO2C9lg82MTl1neVN8WPdDRvSA
wdRnrKNsB0pL0/zH3JVTYfrc/xnOUsRY7vd4w3+yFNBBUn+hXkjIPdGzmznQidYLCH6yRq2MBbj9
aA1maG5/8GKMN8+LnM70XapX02NskjhdS9xnkrXRR9b8fk1EezlZFDzzRAvoMoX5opPzihavZgAf
0QZa5qle2XnSr0L/XqrLcKri+xCgCtG75pkYlfTB9UOTwRCn4h6/Dz9uqXIasrM4EkA6i9nrt8Vi
GuruSaQeU05ZRL0MNW/LjkLApnmm1t3+/IehL3hNn4XqwB1HHYV5u+cKfe2kFdfDGDaBSmesza5V
+1lYUgmkbQT/Vm0Mos6JY5UCZSpRcu1jQdhW+lmKi3aROS28un+qba+uhZQZnMygN63Y1JRNTCin
WdLN63cK0KvLEfZ4055LaUJWLfpX+p4fqTt0kEBVBSLt/+OBMTp/MCsYyDx2z6BF2mHDcX2rxlLC
V+YYVZlCVMlqPgMg4c7VQPh0U1QGOU+U8xoAJHtcLxvitFWO5pssvEC1wpXh6byLMr+aRVFv1v5D
5M1VQywOXwyCAsfDRCmxr5UVb22d2IWb0A2h3mY7lueCPk9lKWNYl3zm0tvbsTJqfdJMgnfQN9Pl
fYy1CYaFIP27bygIroQ44dqXReDQ1sYmX2/Q8jEyjjUH03q6OiDbIjIsGFn8HS3hNb1428i1NWaB
QoGT705yLk5JMDofSfjpkrEmJk6qCHtBsstOix6tXA+IUD5HmVY2vV7DwPpb5f38LrFShHo627lR
+9iccbNQlTi6BsVAeV7UkL6yzxgCUyNgxg93nbTlPSNzNCuorxDj7G94Ss7I6pXaZU8rntTqTMts
sf7SEsTsWBa01Tk6I0OzqWdH228wNQ7MKop2HkhcjSrniRBhwlr39Drf4Woy6rN9IWPLalsWe+NY
4OXmB6n0yTs5tZfic7/Ys0Lj3I0eBWycocqe2HFQtjzfZ+OhsQ7D/cOmJdDC7Q5uB1lAuqzN8GU7
C4Hz4kATPepmdLf6rXLRvVtiLXYeEs3EjBhzQGdhbxTo8ced1OeegBhQ4EK+f8zAMggMAx4cSBdT
uzoKiLLPWRVWGDEjviefxwIezI1INmRKNCjqbOm/Bvpo1nix7tlh99iDIPWxEGtjNHHneBP/Gbd7
o2HgeCGYl/06R8QG2xCAfOfq/ItoW5ArkhuG43VuQ1SDtgjW0mEKgY4w/EAxszMUNmPJbj9qgF/J
/Zon4r5OboxuC3Alr03rEtUWC3+X0OjigMU8Xcx6e+6ssronfsdb7lt00JZrUqfElYB2G4/Uvkpy
8YhCYGKtg2gluG6KCNqaymFubmnW2NwqkNFEYkssWs0GBjCwM3ISJYHTit2nYfw9NZQJADnhCPUz
vH0nwsDQdrak4q1iE01hQdV9xORVsdadQWywBe51wgLgXrlhtIREuTmkvm7GqrQt5V5samMQWzUJ
GA/GrngPqM6nzAE3XezFScEgJztJDXKDpGk8pZSZKUnV7VtGkbKJjjtaBdNypqwvN04l6ndZZ4HT
4EaJDImTLDrbCOgxXsn0gcw4ItMcDhNoR81gBR7N/odnsOvA71AFVlBRBy2QrG4yySKvhQj15DYt
qAPNFG26k3Xmlvtg6dpw6toyIalm0Fy95bh8+lCh4dtXdIzKLe1ERVwZhpOunBd/WgwR8yGYVlp5
3ckfzA5w4nDuHsTezFvnAP/krER/YYokQmrA9jWfweM15nAiT114ws89gwtPud/WIsx0GW0Et+6T
iAiulSeTFzS2JMJLkiYF05qhUr/1QQnsiBcIy7bxF1zpXB2VejKSg1OaAjm2CIYZp844n/NxtG1p
fzNnVJslZeiB5b7f4VtMYfOCaymLHY2UViRm2bM6sUqltVYJYXDv7GpxTspsJLatUIjj9hom6pX0
J1RCw4W1vw75KIcI3fxLlqIRNr/TGrM+d4gAzHNnK/gjciCRPcqamnG9Ll/FenflpES8z8C3zkrn
Xgp6FBYt3geyuPVtE9tGPQ3u9XNBdwDmjnemgolDVHWcAWVGpZuCoqYAb9d1scWFV+56ggLTgnSC
BuFHmp+pUgq4GpAHJWZruhB+c5LxtYeTeTv9ZYwj6+brGfdzAj/k8FxTOLO7IsYzxFyHusoNTgCk
kRc1TsQKecLeGcsfn9w41ftC7v5uDnPMMw8xF6ff0ii5d9nTpxlcj5gzQix7njA495ieBj4nlke/
p0X7lMP5OrwX79EqCpnAY/NTM9HqAW/e0BIZZgi5aXLuzC3kfNWs9aMYMKMTLrxzRYbbzNJFppw6
NIk91MZwHHIag8HMpreqRwAsZ4zb0VKATF2MdCuw7T7sAE1p30+3RhQgOafG2ZV87FKcN9BL4l4E
1ef20edIyGb7lz38+lTR/PbBI7sfSIW9gH+E/bjI/V0zqenl48DvtNpJ4NCZ5GgB1zl25Uyp0VGO
SgMvUsvZ57/ipuqQLjAUJ0IoUZfarUrMR2USCKX7BcXUyj7KfIFJM+DMILfYv+zqD+ypng0lqUoy
Bz699GKRuKPltulmtz/01Uf3v4PiuH86RYWzDQZghh+JotrCg4IGM5asxOPNQRlFHkx31ItY4IMg
CqVOmHAoxjk+LJXF245PYsEk2TSh6X+G7FuwU74aN28nFx1vWUMWIigQX1YhL7nJtPJhPu82ZjGm
sjiNuQ+/FdBf4s0M4jmdx8Ro5Yin9N+iQf5CpM/0jVlqmM7tWOMpseer725Qzmv5ngnDjb0ntu9l
9Zw66XNJ1iIowgLy+q3YE/mOfSSKZ6UzsUbMSEfA3Qj4DAD9YUzUM6BwQhyF6FhS7tElel+myNMo
Put2GzQ6Vjg2RdQdrf+yYG/59tnr0O3CiMR8YQ5PdtjZu8yhk+d7CJDXUqNv+3fXRHrdDekrwjFI
1Wp5x7CLDxO7uUcuR+Krt01iHsOgVIms9ITBIbvQy8owD1A4bbCE0a5Mol1w9VTp+YaOSXVFsENs
8jetNe11sHl3vpH+RtfkB4c+JzSuUWgMas5dk3jL9WcbWToI/zJQ9hKh8e60I6oARzfO7+NR9aEG
4v7avLSvxx0UhZDhXkHH+5pYmXscG6x8Jcp9nvQYXFPITA3uSb8La3Iyh7LzBK8FFULbuTDh/pTe
Xze7NNjIYbTtZvj/22B+q2d3zm7JYpcVrjaYXxWcMFre905gLTnaTgCsPHOLSdXnXrRb8Ij/Tqnm
9sszvKNY4sVOeRkgYfkFG9OnFIl9kYtdufQ3hCKVJxp1BZrFeUzMwqQD//9CyfA05X+dET2IwMvk
uBskValnkIp3ChXNdJXDNuJ7FKEHxkJBINXoE7EvOH26ug6zyzInon2eTtsx34FrM+A5SP24NLmz
CVu3FnHbzH84E+tfRc3Mevz53cw02WXgySpqIHZA+yEAfWyLCS7MIz0zMyVoPssw+Y6gp2pab+BM
7WV4yd2PcggneTAWKrZO4YDD3OOpWrxwFOf0WZAiW9c2266S+vxOm4JxcQqY9BcUEm2BLK2RP1zt
qa5lRiGTDhjHui6EcpQZ6o+20n1futhWdeevgacUWuIQxsPPKlARwxO1oazLZDjYg6eHjK9gjJtH
Ueyvz8N+ztU6CCcdv4RdbH9bR6ldKVpX6DPHvGFd/hkOnQNfqHI8euekSaTuy+sZyjMzfzPENrUd
blUfZWO2HVu4VkIZOZfl6U9i0aNm7dqbA6w7EKEE27AVpkKd6LkixUBenx6kMNDk4t1R2YAVQTpF
fggt5mniMiH1w1l37pzWdgXORJU39qHyczjxZQxlnLXGimXrRa0YutvKbPv9sz8BmwgFTIaLFt05
cY/x3Z5d9A2rDue3xVkl+5m9ZKiR2aI1J372wK+Lf/soXV1G7sIW/TT2DBdk8GSWBqoYR3kJMyOE
rh3G5gqN5itFVSiaYPxkogTb+eWi+X4Sh8sgv+ZFH1aTdz0LKWPNtbyrUAmixflhhO0364yhRA/l
6JHwZfMXuD3AyKLe5jk535S+NYadiOucjGxdVCCKLymzYqG6W6VaJLZifIDEHurQ8NC9JTn5BZO1
ELScWt1gmEhy8i0OT8CH7JjP5sATUMK00V+VCVhQTRK70/yTt1Mkp9Ozz33YnLWFi7bRmGyzcmd9
xPtJOutCvs4MPKJgLYbz0dohILPyDlM3/Vo/nZWTL0pePiJMImIE3hs6XHM8gNITuFTzPLYalt4E
yZpeLwAlHO7zk/P4yfhaiy+OWLcFGvImjSo1ToqkQVRy0BKbVIL2RCgWlgrR0/8jmnFEL5P1nscX
scTYzO6FzcGXcEhQ67dXj1MN9IZSAt4CCNMJaIG1qkD4yks+z2cv3fFA61zwc0V5cCMEEs+v1R5Z
hD/eB9SKQPckpppc6Nr31QKwu61+gogWAWACZLQ/cGhGlB3Ul7dLsmnbQfbGRZwdFgcSIcuXziS0
SUvkRxjnVzJfesyfkgJI5sCwNUpnAKv9LocDagN7OOjH3ZL4rnKvE9dfUO5uI6qPwNJc5KK1G1xd
g65VrUWNgP68YsmyuZ+1YIaloVOVLyDNlnD0T71VMSv66xTcUfrtzawAEDBrDHFY5Pumfw74t9zf
u+H4jPlKYZiiRH4JUuZFdA9M2aAGBHO3AT1dcj7wj6hMhYmtkZ7LfpbbXpQixPFAHCf4Md8f5YgS
ZhhzkLYH8u7ViPAJ9nmpTHGaWdS2mFO+2Dr1NvGeEaijk6ojLA74y+8I7N40JilkwiYxefyk67Uv
4GTeohknBORcxchNYVRQJ1ImXhn56gO+s6Qx2Dp2ESNH+MZUlO8/PJBkGBahIUfYy/VEzP5pXAhB
GSM6VMI1IsCZ0dhmRUaMfTopmUagca8y9EY3/5EI1H3S3cyg25lxpMvYbuC2p0Tmd4JdM5SC2idY
m3khnw0JVmsiPaXWVnVfwS2NY1oVYQjlit4LPnWj5WhJ2htV4sV0/wmNfP8LfjmcWAwqzBZmghPa
Uj6z+9jYQmzWFDeuMylxqIznMMyOBIakvFGfSUczLf/RTC0GFuy35QiBhI10AK6M2OWQSHaSZdj+
dVn6sUqGd7h90kFS0Ir3IuERgYTOhmK6kc3TVuM37XUVMtPdZdmg6ZlaU7szLCGkq55cX+zvJosv
voLTIyxWMLyla2hJsAJn0WIXDvz/L155qYRmvauAW/smQwGQgpCXgy4tiOARpDN8oukLwJCnJ0tw
Vl//6nbiYPHpPBYhHiEUKOydDzSiqCnf9j4pkZXDcmr/av6u/2yjVCWLtDmLogzjTh/A9VuF4d24
2nb5WgJfs6h13VkOy4HxrQZwy78iXXB4yeImWCMKHgYc73M5dub3UQ2/9BA0ShGmx9StwlyYfOwc
wJRO6OgD8awpBZo8g8kXjWSs75vZoZ5rkZzJqUL86XI2hhOGqCXBZ4xGWzE0gUv2wDPRzRNDWS5U
+xviSb5aIivcXY3Z2+9Uzo73Hb4aNsezpjTJlkF6AjqlqZTKr0mHZMsl1ktb12ex2v24jdvvBW2x
l/2pvNLjhPrDfsrgst4IQImkcLNqPmAHk/zFTBIL1wKIJKAd9Gur/ginT3PARjUOnHBwZRirKbzg
QHKxhpwxOXBZ40zSRBCZTOuRdLeKlK4b5SIaX+TE3cO+Hyc9sO7mqR5yeE/cwLxp8LVYI7YdEQNv
PYf/8rkapAj1NlGFz6F2Dlnx0TCjmvA2d1SpgADxrughnWZUdQjJf/YwrvYukNk1f+NJB2jj/4sr
v4O2770ZQI07UVW8XYP4DwtHeFneyQ8NXnj4bHuTtjYRsaXSjyhF4EFLlbJJ95/Q/D1Fe/5octiF
54wSk6fK/mjT8RXnpzn5+yV3u6xabXmm0WgWUVSzOR0JnKGqJ8yZ6kDRfErgYLqGYp6C9YcRquqH
Jd+LGPN3SMhGa/S0Mk4bzvyAxyBjuGYpGam2RI6HAzqLZqqm9zklmEG9uYuSbr0isqAPLJKjM8gC
c7VsOwP7LAbp3sCt+xvQBAHgdVEPHmE/URugQACoScj/Pj2qm5IV0wmT6rEvGi61ZzjHMMYfZIfH
jW5X2Or0oVbZsnLgFheBVuQQsq7LKIP8ah7VmxDpO1xgk5lXBIsE35T5JH9qhCU2X8ZlaEPdoSs/
EClk2dNSKHAr1DAi59llV8Yw12pvMEcZy946hyN7omfBcOZwt3Hnle9p4/X7pxdTZDPrXZPYeTA+
X6xQgYdMblB7FGP/kWn9jAEeCQV9ZqnZBbdDb5p1cvFsQNGannAor9nlvNieljI9XIAJZnsM6rOd
wSNwnReqLo3nLiLRiUg2BCr3HDusbZK+s7g0oCVzh391kjR76+RnlD2rTSM5KpPnArulxZ48pDRu
+VHXjN2eRU9FsWomxvIL9GN8qeVXGW97K/JcjywkCE+JZLBqYATnegv++zfMbemSbbbhB4C3Qp3i
VbER7ilHavtjlyRlx6ey8ZtAk8ZrRySqUHwqXB2dxUmEQIJ/10Jwanpfr81Qe5cs/vQ+fhW+AIBW
uS3u8/fAR8SLp+ugT3Y5JfcdVb2pHYCc35LVP3woHTzdpltQWEG/IF502yFOMIUEFD78aA8nVk0C
/hI1YFiEuzgTiemNFxDg6m2xmruENC/CNPXpxuQrKg002WC0YwvGFToh4GC+8t0zS5hei2amVWt+
w1Gqn9G4lCcEsGCbLmr8Nbof/b/8e6lC7Ed2UKh0xoMvRk7qYSZ+xJtxP70FTDcJ8gQxSobQY36W
25HofDbHBfszhv8C7FG5DLBWHQF92HA1YykkkqWad7j5X0arMw6/7NqkItIGjT8bXarBz0ruDAUJ
VnFzoScLmDQjdIQ27j++LoRqOUCuolzz9BWuySJi3rxhXCtEtaXzD4w45ADHosK+09qAEasMNLpK
byRIxy+4YMVCbcn1ACR2KgZSi3Loz/UA02I3ZPy+j4c9PFj0DnrHNiDU7ndggvZcdRyGgWHOeL04
o61YAgjQOcd2cVEIbXkybkrfeRj1Kf5mtci9osnMCEec+BViub9fdNNQMKrM8BEmjHInl+O2b0ZI
v9wJi9vhl/KR54VreG+UxyQ97dzCnZzT1Mzmu6CEqL/opsgkei4IkcE9xHJpuzHyvBujHk0qJrwU
aCBAkuqpfT09f2SGwdSh8ZWTFGgpj/TahOFs3Ce7XZ1PgKj0E2JiN0/PHN6a4bGf98Cm8JLndRn/
c2tYOI/Ll623bzLhvsgXYubocszpK/lh4vzA/N7kT3P/97VWuo1SzpiS0gdZ1hPWIazFxR9F+vmM
atzuiZi5G1VqtWIjAZNcWCkZblImLz1vcko5J0HhOpNQdBPn2H0b7PtWJp6IrmAKdVlwSoez5Etb
sl25hgpRkjgANJ7aLCk8D96gu4luqS/xJd9gHamQkl5Tljt0MJTrtBFJaUv4f2dOOBXV0T6Ki36K
UOo57jyUg0mIGB7SXXON0NoPStmj0cabheOMfu7IskEh6chKP+0wRYqJvXu3NIXkD/HmLb5VTKGW
F1zoHsBBbF6CmgNVa4HU+PVhRw3hWx7t/BRsfVFrOFMJqoFcHEMOo++F1JcZJgMhLJ0lIHDB4/2A
eFlc1Qq5IF6DiTiY402FewXESdRamBnjt+mYGb1uU5lkgw78watcHG7eiJcw5uL937JfkzkfkEOr
MTqjpetBoXJtX3kWQPHLzUc9JRpxY02ryCgZez06s5q4+Iz2zxPdPk/WaqH9yIf4RIEv/gsxPkhK
g+bXkAXESN6kBnBAdyeRQmvrwhYnoyuJgrvRZEMIdkEHJwkDvWmH2etCGLAaSdQVtY3u7OXmTUDX
KJvePw+SwH+V4hJd8K7NYJ25Y4VS5e495MNn3I9RgP58xY4Sak9oVYkshyk2DhQSHpAUS7BiAypM
UwdQDn0yyXP25P9TJ/YC/alKwEGLRVjndN0HuBaytp5fOOFx/uHmoL+I6Slcxdag8rlKrf1HRZb6
lKjPinWcVOGZg1r/PqnrakgXODoW28nCHcaZzb/bM6gn7vywP60tAIDs3vy2pO7yP6HcEMy6Uu3A
nT1wo0dWA7ykiZt0alPSxWjEcZ3VmIBc4YU3kJNz5k1xEyie9ZXViaWKhLM1uivgfSwQc5P2FthQ
68coG+ofQSipqcddQ4fZYIWbGknI2M+U/Hwe6HBL/7KvGjwWyUh3EWtiuHfouhrU3ftk/gSxZBuv
r/k8nvEiL5dY9ToBeTokk0xsKpv17wDPRjQg7YZagXOEy+Khp1oOICwyCIXV8SPAm4GFoFNpvkmD
hjsW2wQTkkqEwvABLnrvUAo+LxboHCD6E3/BL5hmSWIcdGR3SiROmHGofBIaNDNIGlrRa14KakhA
wj1e1ElnC6+1gFfbN/3Q58AJ4lGUnadHTIL48zC/CXlwHoTIvSIDOcFULbQARjLkL7YVeqBkHcjF
IVWfemWxxXKu2ERgPtMiXiIGLUx6EbOZkAFe4JmGrig2zxLZZ9ptXXMUgOfzAc5o1fv8Tkrr9OIo
A++ximXgj6AV154a57R6roZ4xRAHCiR+9Gkcdda/wjrzQJIj3F9fOtL+1Er1QVuEq7rvRlYJIXH1
Wwzf6H3ASWq/MDuIUZWVAN702dEePTDJpIN8eeLkldHN08pqyzDpaqsn+GMpN/+KGgZbqpgkArCJ
dYTdLLNjPrAgM8kTwakO0dp6C5e2PwhCvR801P5A0bQNf72JHwFXndtvBN+nWoQLTdBFetpFhojk
l1ynBzA7alTuymwfFtUczvc80wNObmotmk9zC4MGSrYi1NlM94Urj0UlEfbc7lXRbJvrYYUm4k3i
dzChoLhzTQ+HGOdOMwHvYEhG/7prbGcBKAIo7A0Nwv43eb3Tg3IvJbSPjDkFR328qIFDWWN1UxrW
XSN9cbLAonLux+SjsgTh2gPKTW/7sDX734180yuYXknbcfnY4RKepYkdIN/mN9CivvifsPR599G3
ynkuPZNxxpSrX0t1DxHhN0MhEW3WOpsGWb9baoLWOxRF0pvcYglpw8wV6m9/ST/qPegT5K9JgAAR
nvyhWolZI1W8qLW5NAIKLs0CS+zYs+wuaNv9XqqNJNVBNprV89ZE+8NDGgbKBTap8eFRBei8nE4L
kc0kqOzVwoBDYuFGYG58SQV+5d1gX1OwNsrM9IX5e6OTFAzoakUPZ2ix4H77K20B1UN8ED6BEHE8
y1GJ/lMNspyc1AD08j4fLaWAOaDMZDNUk/fkx7st9EHTfp6K2tGrPhEYX5toU6CgTisWVgAZp7u9
Q3XHAnkDJNg5rjAuOhjeMPPpoKVHLtrORMQONd3gbKkxvjFb6UCfXTuSLybEBkqyuOefqwr/n5RQ
32HaxcCeh41VCLPnw2jzJ9UdZnpKuQqdmsvcfPeCNmlbFoEGHa1kzXw63atYIYwMjUKGH3ERaNHf
vrjCkK3dG3aC++TTN+YFoGYU9gjJMWLJ9FbB4sP893p4zxUsE7aBJ8+eQHpG9u34kU4mvSjBKYCc
q2otLxAluN9aG+bgXSUlvsSUZrLYbcKnaT+8f1EmD2PbCNOiFVOcfvieCeUlnoJjhOSxNc4PPjFA
cqDGYKUyiTRReG9pvCiRCONsG5SUQYnl3sBVhn3MXCnYL6fN/89KT1xCQcwOvrHPcsDAv6c7iDtX
IOMiAZm2Wk4G+MBVM+d1r8iSa97Btjf8zG9EhxWWWJC3r8BGH1IVQFWQE5AwLuR8DjIMWR64hUzt
OEhRn5FKangXdtQUnVSKDuUIKl9e35dydf6zfEgNTC5brIRoR8jdk6WeHkntMCHuqFBvNXG1Wsl5
gnV6wxusNWJtvK/YxGcMXUpJDcmajVvG8bDkjiKtkZe2f56bremGsosNnpHWvLIV4zAGZEFkiXT4
4a94iF6ndIUQXssP4ayGeKgTk1ttlmvbEGP5TDnOjGlo20EGQ3Ngagp1A2fVIJllBjBCMMkBXr9A
0FtcrrX+a0WOa8wThOrHwH5o1MikVxLNfWN596G29rmDDGCHrfzTHI1Yhkpp847WfkLpL4AdOc16
4pFR6W5SzaKvJFrdoOKwFSXAVsRzTa3S6DJfukdt85KGzd7NMDxgGS1qwrnNBsQSJ1a0uE2EwHZx
pF57Fe3fJ+yvVERYV/uTF/UjOqns9kj38RqFT3wN/LIG0G1Aw80ErchE/yr0H2Bphi6QdTv8ld+C
Azauv6w4gljky4Cf04RXdEg73oeeGvpnfM8j4k1gD4H18/NAEfM1B+5gJv8maibRoV/OlKHCUi7g
3aIrQi6Ej/l6VnLUGdySQ8bQoJR8osKhki0uF8lwEoj4S0GUza1PHNN7SR9D9fG3xJ0KzUod70dB
lQ66zj4h+CYcoFhPHbVdYevMWF3zzS27TabnCI+XmVUhzDeI283Hyi7eV8/vIVAhMwh3PQnipHuz
/xHVmMH5aDErQgs3PqlaF4pCH2TCnIP42NKcqQDfUOi4JjgqkGvGtdULdXJRsMbpKetkGUpItkPp
tRWdW7MsCbSflLKHibSKeov4uJyTKeKzYMfjY6VckbffOyBYqQbR4nUJipIodwWqxBmPOY3JH7Z9
Bm4B29HCMDJIlBsQ6DABq4+cyw32VHBaltRLOCHBZWkoFmLKcJTdi8i0IRwO+iHvabGojtk3LWBs
1+SzeRIGUExU7NUUZuLFeoSrca9T4lh6tdLL6h2ixexhZlKuMtUekoBeAuj7P0QfPkpdMyMqbT+t
T8+isIYrRloCqmPSBFdLJBHHoYam85ZiqVk5n6JIZL4Z2n4Vvgat3eUjkxnsOwIdGbd7Y0jZArTB
UaChtVFRzXXhhWerO+m3Oq7yi8762QIwGyhbw6QoDWNYWvchLeXHRJAZauuPISqz/398bcSPOBwa
f5vJQlAz7d3JqOG6X5oFZueYcRh0hG6lufVwIes4iDM8MgElU2HzPv3DiILWjZMmgnt+trNtBdaD
QE710BBtnjLy5NBXFbHGHwYw78wMpvoYZvUVY/HVTw6WVtQ19waIiL8BV4wbwVA0lRFcNejSvJGP
6Uvt7BAFFD2XFF6wNUzzrUtfYek3vfFfC9mDlrmkPdiJJL5ypieLArDP6BuOfg5XI9YDp9FCp6Tw
wmHD2hZfxEKsOodpbEDjZR50EAmVhkf9eMxIiUXmwrjWySA/EDvUo6mbqjmeXK/DicWRXB3nQ8rV
suQia1eOtM79hz3P2vLfwNkg108YXLxwbHNvamrP9UZt8mX21m9nGE//wcDTFHgGuo3mBKWZ6mSe
ZdEVKsQ/Fkj2GucL3O0G8wh579vt5tWtJhW2ChY+kUo7d+JQqi9QdPDxG/JkjF0CtuJb5BlNvbrL
qieoNI2gfhOAa444EHd/D2CS2a0mNTqv9bkZeIk7hvA0ijgetiXsEyEJ7aYr+6WnhwtbAKwnu+yS
wd3bUVTXK55xoAKja0pE9L3jlhfbfMfpdZZ/d9y3tTQfPzHGkH/qPUxt+jWZfJoHASZGKLH8Ot6d
8imv8M/ns+7hfWWBizgKVxphvw8AlS2q0Z9XnPTQLfVoMpRQoCF9zuXay8gvkrZsBBADvrL5mUZi
cfBOC/UIxlGbz8OGqCTUCFbsvYXVZHzQWdh7hGhyr40PmXiciSdIxh1+X9HwiVUKES1DWxqnvzcn
iZ7n46bZoSwHo3XmzBKfCeoxQ9/LjhWQfVCMqADM9AbTs+YxcCozTLnlq0o6gkwpn9gQvvQ3zDAa
CsecQUFKMAsX2R7Cfl6dZMPrvrf80vRu6yL3CNpLT7MFTG23v5OsGRsP5E1yQuYr0RxcKcYvAe1R
/B0Epi2mX/JFQyV9m+3/rwCMfJT+TX1COY/HMyew651pDTwNgL5SjDesm8KaUnS9mL/J/RAB/cCg
GOHlZ9qTxYTWyE4Yv0Sq2u6ilRIaQD83/Ii/+6aFkOJRMnBiGchAFiEWosEIMVRbcfT1MmTn6Rja
SIB3PLlEEyP8PuVc8KpSEp1IWahuOjiwMWC1KctI4R2Rpw318g15C02NR/AnFSii9crEUNHPIDnb
8pHKn6XrcnUsB2SPuflK/b8fls0ejJ85glRB66UyXB+gGEBhUawlrkO99Raosnz2oUeMMR+spjaC
9gmTBbhcs5osUeWNSIeG/pZ1DV254pxp5yTiD0a58wXSzplZwdVFgMCYJV6jw5TZqcQQG7aq5CEa
g4pcsroI16qurVpGq/NrnLmwv5TNs6Ayy908NJxLB1kyw53ru4YMtds5uTQpUaQwufHRvAU/RCW7
Ad/cz9+xHzA3BozyfP0WbAJYok7BAubxcgbQow8s1GVEGAwlltEiOSlX8ucxXGDsku8AqdhuTuRw
ukFmchmLkTG/u3JShz6tc+Ot6rt2q6WK0zV+qQY1t249+wCxVVxslDrGej+sw6v6HAndyQtKQ7A1
3iUCbmxULXExfrgcRX8cftEuTqMzRA96uxKz4c18CE9g5q85mk4FnOUzkUG9QMxaFmzZgeH8BEv9
aCQxJXOgjihmzBOJs5DJILQFXf1JTdWO8i6kjuhbCx6HtnFNl0Xc4l48RUW3DhrVz7QLt6mqtySL
d9DkhfyhXTGPufFom9TaWn3v28z7ah6XStJreU2RbuN3oma2MDM6+iPCNfLGAdj2wBQ3scfvZuBk
09p+p2sLOKRuv2dAgYbuKE/Q2iKwHPDoSa3qBj8ZotawSIQUIJzAXwgSjR5mLuqI3u0G26IeX5l4
w/74Sw6yGwokPPebSjjVwuqH3veueWaHAetcrAHvE24uT00S6Q5P95beyaxiJ+4PJphqXcsBUkRr
2V4PsSjXhaSQrRR9eQNDbnl1zG7kG3gpkjvqorBbJhdGNh9COIHzIgcn/PRFl44kUOooSUSv/Cm7
Sa0/fvHsz8scm97VOc6J8XH11OC53Fh59MArmfUvQJBuaRBF8twlJtCjhHNuD9OIHvMgHMuzKEIk
7FZqtmI1eY54DEUjezmsifftUCcAyj77a23r7V/JaODIDl2rtwd+CkxPqseIX+jFDZD8nKfe3JcS
dG+O0gyuMm9M+jyRZmgpbLyHAir1yqgNbGu2raKHSmvppRdE3APhXrVTr099qMw1t3rasUYmKHqv
VBg6VvHrnIHCk09QEbkG8bBLsIO1plG+HuruyjZkYd93MMdEcEbkMwKAEXQ1xMle3K40ucS6RaDW
q5GHWT6+QKMuHmPZH3S7QqVgsxmtwflHOQmHwhVor0XKnEt0WrFNisqYkI7R1Buq6vH5vXd9vE4q
O8ukU0jboJ7jnUTyoTCSTsxN6v2a1MYqTeooS0MogoRsAcEgImjVgdeOvHt7j18HZya6ruuQ00i1
zmMLPoRCXo3FhC32xLL9dsCNGEts4KG40z6Fk702ho8vI7kCa/ZL3wB3ivJ43OxmQxqsMIVJurSQ
jWVp/2uSkC8Q8VFG5oN6TCSlMB7jXYbgeAyw54YNZlSw4zdoYitP7o6dR4GxVR9iyZne6y1L9blV
LaJN6HYg8x+o3H4WvHGzugiTyMWd3xikkaQXUL7Hl9HsleoOUePZ54k/vphrxPhRbGNSFpnZVpes
o4A9SC8yzChatprlJnW+XP+Im3+H7DxSCFQ1R/2i8M9Kfqi6DFUhVAB7NNyRT1AokmIU/AfpGD4J
+EqKtLmjsU6W41hNVDilw4aplAZhPxgEGCqO6mgnE1EQ538CYpnUkLkQsDOeqf2f9eUKiVXrfEr+
tQxZHU5dsJkT4TVuZ8Ul+oswFAcGGgciBMcRFvqVkh9jI7rnaSDUKgWqT9RR1b1t5eKeeAIs1vyr
1vE00kNGszVhPoApXcmRQROcUad5wqBy+oP3+eDDy4ms4J2eBhRjxvdX1OtajKeIMUD4JpqiilzA
66alGY+/1CUUJ3qpyAuPnq7ff9vLDkWEDYRvbmXENhfwUAaIYclXbsy9JLgTzjXhD8opZtYhICUP
vzQ7npM/72apiFmJHN2gOCPwdOU0VmElzZ1ndSOTt+z0k5zwGBa8NCvyNH1H+fvP0QWh9p/1U0fA
9TLSsAt2tQhBMpvZfc+a+AVwU5fQzZ29kpC74Xm1U5mmHbux8qJ/2mcKZYEYbr0bqsqBO4INk712
rvTUEw4WvdoxuvEejPmCGXh0eAX9kyDBN6vctCKy5f4KULwryt4nw+pJCu+SyckEIaoAzEfHp+mf
t7yYuJOeJm+Vg+GbiTAh5W5CCLxXB9z1lvmsC4YMQoehgQUoXtknefz2i1Yn4m3n2mNCx25pT0N+
fkDsobpbun7mC9ufaMt7D4VYB0Ffv3h7z8zvj44xZk6kOhwZ4tzbebqo+9vKTUH0xUbitbu9Z9nQ
7MSnfSl6c/mSO8m5xEztZur/BIBaMhFjterPpwfKh18jirBpPNjq1ZPnHoi5RtuQOjKDsrTPdACM
BjXMXCl/WBsv2i6lBrm1TaxEz2EjildkkSayWnLleOdYVsUodMF8myxn4oIbxquTVwoYZRTfKIZR
J10/vB1EjmJBYAj7yja1PEM1TbfdcHWy47NFYdYYyzaYnTcNfFGjCKgTSJ8OWw35eDsmn3eSNYwT
bSATKswIrxZ9X6RL7mCmN5AA6RdTNuvydfHY1GktcuydqJ/bCKAwdGQUk8UTu2vHHiY4aw1krspi
OQua4R/0DbhkcR3hynbMd702sue0sMYIp4tfOGw+t/b3wMfxGs6Mff99SEoEvgayj8LbzvdDBm7e
xIR2xIPvD3t3KJ5mlUe1SGAm6tndoj08k4kv8e3/sVoBLKj5WTN3GfrCsrt0qsCSyv5TfdOG1Fl1
T3CvAaKwmXQpg4MUuh+NAyjnMxmrsqmcAeDD6/fk2fqPqg00eEn9Hn89AiFO+jfA4TaeH55e4Hh/
M/CHaWBEKk7XbcpLc9wpPfLf9Pt17euOFyLlraXaFP2x3QWwDavArd3l/CrxgCkNvutDtB7x16Vk
i5nmiC9M6sUaRbQeWTCihnT3gNDmkDUSZS1/0f25NfOOJ3b6gL6wlZsBRYyYo8Ya3yOYrSDs6kfu
qQrxmDpI+GcSLnXhocuvBFW0QpXmcAj+j5o2rxKFbDnYRf2/PZfnp4AdSA8IY5Wbpi+vN/uI9SVp
kB/hVC8xX3tStpV3B9l3pFzVSPwRkkEPLKybnsPdh16IpwNr0hqDFH/j0I5NJmxjxY11sfQJVeGy
PXyXBWPkUmeU94FS5UNEx+u+wc2bAyZDRliDOdjLp3iZzTc0/h9WQziBpT5p/zmliQJQ7vzhC2L6
2af2u0ohitvBfDdSvqmcNkOc/KuY51trLsl81tWNSXn/WCOH1JdnzUNFDjNfGjq5fL1xLPF7Vg4i
gyS3Kd3xy5Y8/4ldTSK4fuNm5IBfMOdxPm4aN5bZY0dYU8pDIg0H5y0JyS8yUl7ALfp2O4KaabYo
qziI6N4Y4LtrwpSV3fL5LnjQWVGCJdyQlbwWY4+QLp1zisEBnpFKE4odYcLyBAfOWki9f7Y0nxXZ
VcIdMXYklSKufM4t8n4zI3wm655S1RFHiKqKxMmPPQzGJpyDm13144P68adYMw3vSHdxjzh4JDEh
AWLvLYXLSY/+E9MRmJCd9fDm+nIsSPQ9u+ihCeqJoNQ23dSx/RIyglm9vXH9V+Msn2U6iI01q+ll
ibpno+X2XbxfSIVhSPlJnYqmoR/5EEqj9qC45juxoeewQ6iaiy2tzaNtMUYr9gW7T8Odol0lX/DU
dodDFCwehDKz6Zv2n9xzVWokyoScUKarWobDN2DTw5Y6G1ZxCSWBT5IjKRasLPJ08eMg7zCNzJRG
EPuruzfn6aZeAda+fvsNHl1NuAtkD9w7bCz/EMwIDhqydVxv6RZajCm5tK1psCCPL6GbGhlmmRUL
M1Yzj5wMmqQ4h0Kkpr14tg2HmGFlAPtrYteJPv1/Tt5gxlZ52zoIuYjkTx0I9vKFya8FFGHy3RsK
k/Ptv28TeQ+rLw5duWBd5NtPi8bE5w2QTcCfOh/RwqFW46x+OvdP26hmlz+V0QQ1xH0IBH35Y/jU
5OHq8F3Smmy6Q8OsCgCK/Lu26PIvij/dKKsPr4qIAQXOBkDICSjEEPBEwKX4QQSRCWNKDKoaVwbv
sd8XDJc0fHfRMTtnQAA1DMEUCIOkTqe2c6pmFVrTIcvsj2JLvCclGbkLRPm2xe4532ggdjHh4CJ7
a9MbdpzejmAyrh7SaxIR3fuEDCqnpqR06aunafZepcSm2iaQJ15zmQaRRJ6xZwMIIrHOZ39eOm1i
i2ti3o0Jo+WRYCx82hSFoRw8dF01hwYoiO1KarotmV1eFyrbxXvJpZdnFdCYgNuRcOyBQUvdd9Iz
zAxJ/usGITYwnjZEhR2XwBG82h8m2xsszJlPR9zrymgbYK3WUrS2GRAHsGbXPB8sbdLv9lTsfsiH
ySAZcDau+NjylTTuXL0vX66EoOxLPmzOF7uftfwdH97zH/NE3uoJWK6g6WBYzAHNJbYU7RPbjShA
nhOLLKm28SQETq62UO9kq9Z/hcbV6BCrfCw258Di35vujLTRlqfgNlyEwXk6++kzxvHdzb1Ksv8V
B+rasNUmSVXXQYxByk6lfqsIccPQ6LY1ATxVlFFtsHEVLN7IStrCEAjKw3gkuf5KRra6kXOAOkoG
nD83u5u3kPWK7Wl243ZAlfCvoaJ+Fc2PMiLyiUbifvVMtW71xmzzRii9qPvDFx+GlsWQjgj57Md5
5F44VEpAA6u77Q8S7MIsGfMxPZsslzWl+jViV9hFSY/nPW43I7CPz/c8B8OzOgCtk0gg59t0Xhek
4ECplSuKMsVNt3BhyhwbiUMX8ZUabLKFVgjiDoUq8Q+OsYvUyTnuPsm6tGIiWRmocUq5FUhUthsv
xtJaE5aS11vYPy2DbstuNAlzzWsdDO2Jm/zrEDviHAyTU9z4Fq8JPRpM9OU7qAayXlSuWkL5naix
N+1YNB/Gh1dx/fo/xBDgfQBu3dECg3zozAEh14AfCG5VARBoZQILlSxDPFJ1CHzdJSI+4Z7SM5bq
DAwQ1Rdt8gaP0KI2SJp/mYefrNLcEeSPuEbPpbjdIHBHaD/JKMsCaAoRWa6zB2SbVhYtrdlkyrD8
H1ezP0g9IAGprwPumjwNm5M8PBr/YMZ2TGvHWX72savJoAPcX2uaEWN1I9/9LGh9emdHUh+sPv7G
r6mNRnRjeAm7HFABn2CEgxmTszAXuVwltCmovpBZaoF/CMQlxnR6uBfMLrTxDRnr3zEopWpaqjAQ
XYUW5Hmt2y2o1d3G3fN6tn7YRlVJ+NNxPchPOx0p0mvBxXUa6I25jXTRL9pB0SIrXU3XzblQBkv8
m5ccDapcoM1knzgHN8SCpqEOMS65SbrvwWBnTjlMSBeERDZfb0cSDwrPOoQW1XDbMaS5A00iBf/K
HPDuarDg34QjVq16pxgCIVTWNjYDgxT33kXhLj1KTIlzT9sqNaRTBA+6HfHp1ELgBS4mInC3gAQo
gpDkaqdi+vGmWkNLCmx/2/7r8xDuSRBsR93qgfpuf94GhW8e5Eqs1rF+516H/pWHbdINvBgnJ7Aw
igtU85KoJkspXuZkPz3xRF05t4oge18x+mAByE2YO14ozO+CTiS/PPfQPUXmsbMtfQwF1D9J0cht
vAqZSRGf+gnMf2G0u++du3P88SNAiAIyA2OuUq7pJTBlTeM+YVkw4lKTm8wrJFhBpDms0/rVZISD
80QOyUdkbd7aVPNVzSJCOT8TSndgwJTpn0uc814YeMelQojXxgKCvv0bWsEZlrzCPPNeoqe1ifRO
XujDqqjPhm4zSXsw5Pm6pzaF3bcvlj813B26CX1QfoviPRlFSpd4F5AMKNGt8xl/FRrQnxrGz0U1
IMET5fFvdB+nGWjgGiOUf92Q8UhhSuUyKyoMPh+pILVRJ2JrVZKfngDGzcaeqm19WwIo2kIKD+z8
OOJKxvS3XWkVBC6OHz3q9fxfymvxqUwTnP+qkOs44VLXaG6LLSaXxOKtdBF1PPWM4h0Ow4vjqpcB
k4dzBVjs814AN1YBmfH58L2MRCZnpJfX0q9PfZaaqgHC8W0kyU6VLquetCbPtweb37nW8dJfdVNA
hNqwy8zgAOZqc6oJhOQybvDVhx+pTFeAD+fAqcYsXNBQaHDfObdFROtGeA6wI52i9eyVesYciP0D
8QjdOyMWVNhU0ABfCrHmku9t8hm7ACo2vKJWQltjhvA4b2tawsaa0pavyePy0Wi/zVmzPcwfSWeu
+TkLZab28U+bLDR2TuzlyQHB1NLvwjBQBRXCM34byiLnFBQv66yO3j47LrNxP1zikjx3JB8kWkbv
JmmC/dVmET1/JUREdNcuKMSiBxgOMPr8Galggl1m/zZea7v6rU0sukpto4pJEUGgCUmx5PxpxNF8
Z0A3Tk0GZ0IXVoW68Gdm/1H+PLzmwSdB70bg9U5lTldtL+/vE+rP/t8+bFH4sS2H101kM8ghXkoJ
7BCE/c7kN5dGqD/i/dP9yB7OaZmBuzYcBsp8UoReL59SSm+DE1fUxlzRr9BuZpPIfVCZibfJvoXQ
oCeUccV+NE4BjFEGPFVfQpCURK5OHMJ3IpDZEyGrACHbdh/v6DNH3jEaFhu1Q7qFGky0FgLomAZK
KZRrvzxp8m23xjInANbBpZmkiAv8fYhsfH/9IVNpy26zrvK6PnYJ9Eaucy9ZRUqH9kQzOKhWMbhm
tUcX+jbbGCOxBZifimzoqSRJRBCLNVVVA7QENcF6PR5jhqt/4Z4Yv9+e+47UmAtEPn8cudVew850
e34QSvs1pMndohri29gFbq0iofmPx/m9tHI59YUdTz/GfI73mCNQWlUkm6W7atmftwUkbNj30DVN
JWsho2lpXjINcV/ojNoNypW0g9jtQEAFC0eh/eqOLE9GZoIbCIRmzCC9mA9UAF4+E1PZt0r7Stzq
NnW47jrR70iKYs0dLgcBqHY4kxr9kg7v3F8qPwC09XMQyBm9y2Dd9T1M82oM6sxzi4n7ZqzEh/35
yCrd4M/lSkR7VK87D5aDFK3zADdRkUBqQcSTXstihIRdoYq3o0weIOEnT39u46Is9kwRGL/ekHB3
Uy3cAT3Jqgk4JRBm796fmkaIK1xR8K2dAalc9tK9tqi24kpCmSsgsfcNBCxxeyutR2W235p19O3W
06C36FpYwMRTkiNn7vzHlV6AgL8MIS3NMzkS9hl9CxOU3jC2sIGsUS8WPTYcbnPZBo0bUQUrpcFv
K/H6FQECEpPIHJP2MRe2RhumNeSdclKUO5moVjf3i9c0IEzhYY4i3iopFRF4vJoNF7ZjmCCSd5qr
9XEeJkKs9ENR8cXCghEKu27ZPlVTBVktEHP13byohqoOUVLEWUj+lFZAaBxAf2feiMpc718UFVuq
X7K5K1IKKGDm9DzRHe2PbVrFC8Yr7f2MY+rO8BstfXElSF7xGuJ5cd3k+BBEvQ+arsH200SDvrHr
F3QXeFwXhdxSDki+BU4xcjvT5gshgbXe6Twg7Y0NqR8tvb8qfXqj+hTVZkePPvGe8ngNBawi5bqm
OIXBcxF+ZLGL2g/NLPorIl/Hij6iyifulIbECFoZS01Ge42D2Wpu9fX6Dqxg7KbTklHsw/abuXKK
Dr09WGtPOht4lTQ7Rf928T4hfcgrHUDrMqjbGi+qsOKxZVD/YwhMxZE1vJkHUYk4L8aEEy+nv730
ROz2wnzChAmhGJZKGx4hnGV5K0uJnjl6tCE/BM3OqZ0Aj9Y3EpBIy8ilcHyU6GjtV5z0CnfIwjs9
WABqpbwCkkARO1gc/RwXsI/eX+lFl9idY3vKRnLa/rTAsncToP1lNm7Vifmu+MWhcCsbALAPs+gj
XwNU9Jgci1bCLIJkwDBQ2QNPJsEIBG4lZAjSamApWGkdL8ycRFYku2utxTi8WSrIv9hgT5eT+oQ/
bf4N80VFOsW991y8pzTmNJ49T3t5WT+WaxyuapVh+FSwM76jeWnUr7Wer/30LV5xiT+LAsmAc3IQ
2VMv778bOjbddgavkhvPsdR7q8K+HPfKZHZfrmAqsR50efavh/BIxwohqmoEsrbIFW7U8lgoviRg
oRxIj5y/ljXpoScA6H2zb+wt3HiTOyMqJhUrD8hco2LCqK0XkNbTvPlm9hGk5Y9AX4CfuFgZg6z6
bzjiDrxPILoo/nzKqVrLUDZAMt9BW2HNHNbLg4gCXRLQQJqMLMCcemoRU5x6+mCwoN3om+3cnhS7
4v297Mn4DrZEP+HprNdX2qqpOJQ02rZ73PoTd94Us7N69gFnzrRaXgBHii5x6daXWFTaSnH5bXRm
UQjj/owWg2VhnfYFg554qqIC/WU8wheEj/tmxTJ7mcS1/XYFQdumFihC1TmNxJtnoadv1v1WeVb3
VTuhJj6B8C/Rg1DA2uusu1mE3Jlyymvnr786Mww3Ld0O1Jgp4TlpTEdGRBy30PqXJSuKiI+HUX2/
ErBuZjp6x9ljyUzCbco6z5tIo0D0dNs2mHiXKqefAlBF3LlAUeSux8ri9NJt5/QUZxAA2h/ZtHWr
QocPDjvq2bNpOWHJc6itd2aaM7ohUhybYOw+SN8SGtBMm/f0gwLQ0YapD3stSyXYfXBtdqpnl4uF
NtH4X3Sv6Ed6M3EayYdjvkhEcoyO4UawTnFcpsh0UumYPq3N4D9riu+BAPRipHaApTL4LQdakL3e
57WmKncnbv9dpx1JKPdPzJe/G8tYvJ/ZLlNP3xfWxiE8r1N3eO8qR0+aSR2/fH2VOebt/KrK00h3
IInBNvgh+bTOF+78mqbftPV/xIpVH3m3FDGAPdKLKlS1o3dpRcYFs7B71TFJ2ePDK7Y22GaV0AYo
jfhamwub3Hmc1b3FJXEiqGLh7h6+GoRsqMIYhDmwEa0Af46DzUDttJAOHpWlVaGVNR22vWRRB95C
+ZMOYod9tYhXy5045NMuZJ8Hpdw/OHyUlpOmViUH3RSSHv1Bu90KtowH6OgdIrXbiyIOiuzqUWWn
XA9DpcjsX2a96f74ffCcKYe3aeoTHsk8/izGJ2oCU04vU5ZyVXoSOR5eE14UMDgBA+06HUmmVWfx
9xBErqiKfGjKC+hRjgiaNj29A+lP8qJx9TnvcGCS93UGkRf6kSciAPVGYqOJI92TuJbYyLAY/mMQ
72viiMib4kQDKxpkkMApDBA5+dLBQmxHfWbi2Vytg/bv/W1lRpn8+8k/fF1xitg2/rLMBQjNmGWO
xXCM4vYxRTHtoiCiFYfaLB2GeVPcUD48WtbEmjagL4R3R2l+IQI/FxW0sIP/F+q/A9ZxuogyAbPI
evrP3Vfn9Uhx8/HKZLd+jEww4rJIltnm8iu4ZBeHSKaz3Dy53lZQ9KBXMfgt7jV5CxpS1KZssMsB
qeQdlONwKE81pLhoHyhuMGOFvVvck/anaeRym4GuMZnIi2p+MOvTLsfMoeWImQp312wIW9Q2Ie35
yvS/AjATSrxUbsAqL34PAznlWWkcVYUOiNukxTl/+Xq+fqbOCzaV4YcnDCgXnWUCu3YPQnTt/KI3
a6ThtidpEkagWIU7Ww/4fgNwHSAax+Th1Rf467JDNZ6MDM09VgtWLCHbDhsfiXzkl0CyKSNMD47N
D3dKp7WweLRjSGLV+oZHuMoYq10bSXF9L3pYTji5uQwPbjLjbc2XMd5hFMp4jCWKGyycEgdRLYDu
dhKovMuZ7fZLQM20E4GvMUN09KYZDS3xxjAIUqxiZ3gWgUNpEf4jQG+1WgmCuGkpnWfGqJLRqse/
m1gwRzGof7DLQ31EqRYhZZAMaIq7/B/QOqzuZ5hxBVg+qN0PSSGkNbfF7IZfEKYs/nni6PUpKtET
WUnLWBKNwkHvbLGM49Q8GXHxaYjn1nZMgkh/I1H3z8+3aa4r+l3GCiYFPfGIwwzpWuIxefR5saLz
XAN6RbFF7jWkUix9nyuwpUMxWh0yVbtEJ8zAvx67Vf5Pi60q98DKrPSysviOcDC2w+diVgwqZ8ss
CvCEQ3cm1f7Nd6uFjZQobtYVqjIGrdYdS12MzPkAMCXoUaY+ot05f2pDf20gkVwCJS9KwHnNjkhU
BUFaFQktb+FhsZtx1Njg5+W9KBOqh2q7qJyQHdcSmlUc8IS4tbU4ldT3bLEkEPMMs5kVUxdQU6H9
H0uaVvwCbE6odLO/04XUok5y07gR6sSyz9j68ssa+x+7mH5clX7MqjJ97HKm19dTyniQ4VydaV6O
eckggelNgyum/9vsRWAKZ3sdhpDIp5ijUOzogzJImN0LhWTkuo4hruZMj8pVXGH4jtULUXLtmCIO
28xxwbEaUmNxhNQ9cat4AzpboGlcxbncLi0qqtYc01NAOC0b2dlTJIoS/LtUqVrYkh1DdgvkTlHK
bVkrlPbl1EsSLIs35NTSuyFYrpL/QJYbArOKdHVEQ7hO5XQ8jMiIvwHzsfyg49yZi5i8ddJzFARb
CsgL1sxXCDGZ1u1jGwvi1i1KhhYGJzuEE4G+L/5iZUqmhOJY6yICRYlUqQsgXBto9dcbK0BBjDYV
Un1GsyhQwxNcwcE4Ih/McSO++iyXa/WQrlDedSmAqCFSBjEB+TxlTifghha3yFGexYqEcSc7RaP3
svUcNM7ktPYTT2tZCdpV5s8pgTrd3qCM1wt/z5t0bZIx0PVJb1XH/pTQv0PSYxpK4XHjxP9shZ71
CN4aVEc8bHmm88zGDp1IJwFajU2/kq1wxU8kfugb7jt64C4heyc+dgDNErZshucnpc8ifvytsNE5
a0MKa7cR0HfdH/N2DlqskSTVdyZPS3YjZhx7kpfXTMtpr3Pi0mqxv+kZRljl52z6cVFTUfVA4MN6
5hjteTBRshBWBV8lr0LSDwx1z5q8EtIrIfyli1GiFTUlmpMI79BlTln2MwattTCU+OqmWpCg8z1z
0o+kI+xPWu1NmLbA5h5p48i1zM8D+rmlbJcrhyVrOqKu0AkhOABRJvYaCtonowRlek0axAm75RrN
NuAVB4olVxMpZLZeIN++gdj2GkJlpeocqaniz7VvvvfPnphVtGmoOTMZia7vZyQLvsvWkQ46nXzy
whJG7DqzfVscwAIecd28pbxfg2Pr08stAktXO2gyoIwDcr25IwXkEyS7PJ+5U7s3XVq5edglWNyq
zLgJbNAdD+IFy+Aaz7ZqUZZSE3aek6676EgDVvV1vBzMW291/rm9pxBEot9jldoZ6bvxZEggqcxn
dV8xlCZxNXjuNk5yZyRGQ31/fiLMqWM5rQUKZGwRNhCn7P5lSzm7kV72+n4dWXPAkjtc2mLITZPV
BFGm3OLIP4copm8bbhIDz1IRnFQ5PiwPFMFxVgJhPLMpZPRSyubgNukeU9lG0OVJ3fx5e5zpOOBx
+U6atT8m63Tv8lYkT6Z5gRa0YFhXv4P2KhPjygvwOLaiE0Bmr4/K76MdATh+U/v6NYAmtBgRceq5
tB6POPgpm0GSwpUrJBlhP0xXE7+y8HfFHEVVYKSrpIUGXnJNSTB/uvBtt73pL42BliXnX0az8WP8
FRPcf75DxQrHYl/BwuI4zEtlUHbZghTLrS9gn9bTBeP3agZdoEt+muK+GiqoOb701YhLmIwaenzH
cynqWxh/787ZWSlgHM7NJfQdAZYJGhb1Wk2wUP9X4BFetAesrbH157UaeNC7puqjBbsgAG4Wdn4y
4WlgMXsoUQDkurL49Gsz+5FLNnSEhTd8Wdl69vcsrbiqzzVmVGhg+Y1HdI4YehfxrS+JGdAHHoaT
Vx5vZGYtHh5bN6v2bfcoe1bA/QvkIjNCOwuJif3IeWaJx90C7uTgj0XNHIt5/hJdYBDpRuEx3sts
Rq11fpvX33zynw2Hx1RuP+qDqrHGEvNxMLxYmDnhXuQxmIEPiYOoUy8Rx/h6UHyq0zCPxkWPfIYE
PhrNILlo4v9nWy+bIFfPKDondx679goXg0D4RcMAtcFH7YI/xrUh+z9ETBWWFJlZ+eFkuwqy1DFF
+sg8ouq+czfq1C9hySmq0nHW1pgFclfmyWlUpacoFCmHv2D8wqCyoVD9ynLLNeXZWmIfDfr7AKH+
0iyFjt12inZUGN0Qx51jgvRfBIjgp6ITKtSlrSANDXCbBO5elzbLkz3S0n936XwtdSQXnUcyRXPt
zTuelxzBlG/Lu1XSCM25OAwOY4ge64pa1Fip3Pp/wsa82/puf91m3IDLcXr/OYkkhuCzSYMXMEaJ
rRwuwtiLStrwDeSzQSNliUv6TCyL4GqYP8FznbSH//kK7l1dJIYtenri/BL0RbzU99iYs/SkVBc5
DtlIZTReZdChiwQx4stv+wDyzZ1UZrXTNXKS6kprI0WSWl1nTYPasaMoD608w+mKrl2qh59l9Zjd
34P2FXSJ3EgB11HATi/fNk8YToNwUJ0N6N/HRFVICSRFquUnUZXwP6In/KrO8/nJqcYTK2FVZiYy
rZ1ariGsg29BvQ8Lz+80wvuQGRqj99NwY7ubiFYyEWcq45JyOw+35lx9Ubm8ufQLj4BuV6xg7Rwr
3lNGM7hDTcweqwNJEX3sOl2T9Mg5uRmZnlDxC43zOFyVT6aRv7IQAK7gQOGOStV6RK/LSyROtxBS
+ClRDD1gFZgR2q44yzMWwmoIei/gDZBweN6m2Uci51We026Twao23bkBXClCo2GR1S/4yScEWpwT
T1Bt7VfyVicltfQiQIvGN0z8ngDLSKTDa8LbbrwS1ZNIliZJ9kalwtcjSIiLZAoYBaqnZcZKMMX1
4+0TiWL9vpZyBNmMVYwozIe1GukcK1m+ToQL9S0mkS9mzr9tSE7lVS+4MUTNWlbiTYlkxiQaC0pT
x6YhvlWo5sSqpNaWVb7JHeQFLFW4chAxz9TE/J2FPLpHUtUYaMaPKwUWoRfq4LLz3ZsTF2Ju2/fR
X3Ys8EeNu61q8p4xyVl62FU4s0x5Ag6nLe6AW5K+Ws/BBz3uuvcMbCw9S6EhOtNSOOQJwWb8PxOg
9Aoyqgsnm5VLvdxcEHmaEJCLxvoONvl4Vrjs7U88mKUhpu/5IptXK+toIPFIHZOEttinLlKPXE7W
bkC+3Tn+pzaEGi6fMjqGeeUIJOEMekA17b14y2F07/KgEGsjZsnQN4PVyjCTo4KXbxconDI4Vusc
MYdEAxFo/mlMkIfQU7fy5w3d2NvzmtbBEINJafS4Vgqx89YVxF0qgs8dA9e8ieReRJu38QHJGYgA
iztqZKcvCklG0lU4ZHNCFLNTyiWEDHUceKSfNJaajaKllfkmHCx18wjYFctG6E+D7OwJKCEASNy+
k92wNNS8bABCQg8ScW+nLxk2MsFLihtv//PNa6YLDTyFJhSoDFtb2beCtfIUDZiPk2UGWFBIXI8m
t3ZAF+ddOEmzOLHp/VqrWAbJFMH2hb/POeAYwX+bm7DMRU8kK7rCoyTMMEPQbtKqFXjHes1NGXF5
Ue6cZ5RHxmdsa12//u8FJ82Owdavq6d6L/DV1d3rzvapMfIhefXotokGr2xeho8XSAtvVqbHHbGQ
KlvJ64T+r0eeeZjj4SnEX+j6QinN6BPHxqbsVokbQ1DATpyAjZUzUN12+i6MpEZeNYFU3xw7DSHa
mYKAo5ylTHFVrFN0Nc8XGPhAA1V2xXFYYh4CbEpPlrlPHpDlpzpsHsM2Qo3weKKMh5bj8vvGGg/A
/uH8wdqKA/w3A8rxwKzUfk/YeKHiS87nnvuauKfiO8+lVtq1RA09maKRU+WjCfsQj4WgqTwjO9Lt
osP4hDeahFRC0luB+g/K8IgU+KjyAq1X8no3cDwfyeOHBgKYicVRt0O4JyNAgtSaP4PWiLT8vk+8
b6gZpf1+6yt/nEMcxnn5/Ye5AbNE1EvRrDSsor/yTjO4iIZjuMb4+CG79vBTMi4SLi/H1+XIbmBy
02i/PMZuSDC/XdqkZRdOZAPZV7WVwSrFrlbrufcdEJREt/RSnf+LWQE430OAAM8BqI5DmGO9WHyW
tD6LIsmsgMA7liDh1IZebi6Az8DfhjHu5mZMi6FBLCD7/ySAduifR48wR/rwZuLdxRB+TuVZUkqF
/douOeZfW7s8W2yEQZa7z1TwiySsWCUvseWuCCYAO0AbBVT8jMjef1285HO4dQAycL/5NviQbCv0
mT5/5YynVYwst65IrGDCRkYbGXxojTZTTxDZf2MdvmrT+yl6LZCsKK2bwRmyNQ4O5qKivruY4NVq
umRubmd7xZC7drz101ALf83LsmdEpHpmxPbzoBj+JPQ7TJTvGtRmGTTMug3TvFUn2+2/fBNBSvlE
sswz5v+H4LzEB+gLTnPwlc1/ixGcMTrBEgyDftiHVtxMWSsVy5fP/zhhYhc910vliFLRdYCVrsY0
xUbF98OIa/M0xcbaIINeoxqWcTVj4bI1ZtZ2zO80SIHv9OTHfyX4UILXjMmYqPbtGKSM8WXfSEpF
33qOYmxOe6tWmp9l7eWKi6LV5rA1cEPXOw0Hq90GkEBKBSjXsz+lXrlunZCuEMJZ0qcJloOGT1wt
y3ZaxeeMgn49PMzE56F9hKX5HOIlvKXsq1K2m1cWz5cr8qC+OszXZgm1OW5hEQrpBEVBAkGnGVbN
EzYn0GPNEqvHxPaGvc16q7zAQa1jvSClXQiSncqiT72FL6YxYUdUvweWXg6lU13xBkYmP9X3PZ2y
qFf5rYfp44IVacQ+VvUpDnv1uFabahv9MKAYfV042pr8SvIkHXHYdHjDPnmR6VmCxuy3XZStmb++
zBHrXqDKPkRS7TDDf7ajNIxMqybcc4tx3PlFx4Jtrtm8BxAtmN+nksylPhmi8AGpHqGdIIsf6l3t
v/0tEmR96Eo0lEDDC0WI/pqJ/T9n07/jZGCJICGTqIrqhtVIr9rYJ+E1ev+76e3FZJ1iv5H5s8zk
d3QnrUqoklXC/N+xcqNSGDt5LyGDYbJ3+Uaez6Fx0BTqK+z2Z9wnFS6axqqai6k7mBaJpwdNC13S
pm/M7T5KrJh88uwBfkerdtjrLkMAP+kH0oVZZo5QQTqw9yNH2/blcJTVquGm2RRz70Y4V8f87zVz
BmjKq+WMnN45bsI8D2mZRKs2MczGUVA4Gbr0CZaBDbQQSn2/jGmWCv8+IcW02b02mVK2VZ+gWYKn
9Zimfh1UFLSee+x8CECpPD9NaC8BhDJ0MVA3KbIVX4dW4bJMx+PCqQXOTiKeT8tR5XlGGHXtTN+5
3HSZSDxCgh9M+sLMaKG6o1dfNYJN/gGM3WUEn8rGdFDdktzEfUMSQ/8dzqrl9LS0j730L68L1d3r
z7aS6S1Yl4VvnZYi1MZL8MHaCZZuORpLouIEf1MliRgl1PfPGOhfVq2Iv1looQR7ALXTKv/P2Zjr
t8/OXE6Nh15tgtP/ApEEeQTiZE6nnqMRZMuiKJAE8erftUokcS2w5/ze04AcucqVcKRFQaQA8llw
5WWlTP8Ol2IbJg59tWYRuHAGTtZIl3j0fh5/r2K3K54ASyl+tzSk4Gmil8j739oWN7xzkGFkg028
3ZbDzlljf+DZmgCTUOD8OWRwA+zGW+ATuCvLGWmx1G9YlX+arXotf4DPeph5FjCuC1etHeJP8o5p
0tteE+CHoG8cgA2BYje2fdTbaOBdtVGHlTnE2pU7YH2DCy70H3mZXbWA3whYMbYy+he+CdqLsl5S
69YUYagRIHw78xizyc3E4eMWbf9jNcax/R7JQb+YVzZAuV5apn0n6hDa0NUn3Sddo9CJ/v1m+gnt
mf/qpGoTjbNpJaPRvrk5mDnyD5QlkiXyVqV3/XViw5aRw5rhMCe9lX69MF8I9otELmuFDpIDfSMg
oe8SuSi4li9XUCcPGHxvW5dUXHJlMu5odZ0TuzZI4XoezCcybUC0/SEjvcHF66/BG9Cqa2tUosY0
R5zRLcaGJiDq1YuKTTptJz3y++pxjS0jiSXImLoddfdmHFLFgIA253PMD7FSW9rmPhAk+WTGYKKd
EHtd6tExPGb+vGrTa25dbYWvI27X4Y8YP9Q/ey2y4YnIC70YePRGBZqTzjEAC3pgmZae3wVE9+KE
on3Q7z4OgWl3GmNbQ03Sbe8/MXGKAUCo3QGYIFzvDoOMLw95RYSbNEbXeE1s4wzjyoiEjk6NHIc8
V8jV/pDQzVin/jWtGMse2+JGPs7hDIl9IOkQ9sEcBdVnlwKCz2LQfiqALEzzjYZpGBmMbq3Xhlvr
GGmk847cSoUkF/zmq3A1czupuj+p+h5ZS3mnfk8F4BnuokVfuqJJW88sOygp7jAUDv2Jh16u7pE+
LpL2FxF0uT7MEW2kb2tKUXUh4dFgNY1h6UV+aN3v0csodrgclz2cY536kdv9hmtMEtXILpCvxwsW
jwG+N7FBCoGjSmhBId5Ni9M5hPkWBvvqwOwLI+qsMD/2G7Z+8s7RHO0eVE/Bqs/bsgZVwjrrPwZY
QIwJxFUTHU5pXhmNrzDi8CKuKcljFdNiUJQ/W9DXxlBwg1Xfunjmi6v3azHz3NeEsFU80aoUyXIU
rwIW9SZGQbi/GrGj7EDXZ9hbTHje11sKkSC/AyR2IPJh+Tgoy0+6O4CSlxC+axIDp0Epcv53gfVA
9msFbU+sZUYATwDTOK9w3d2+WfXDcctLmesRXp0JxZ7CUAOCZ8iArXhtg5d8YqQPbWHHLI0T5RT8
ku1wPwFboydWYhM/nKi1HuBgo7CtEX9FiQVIl+G1PYhkN27eYghrt1g6l+kDVb8Y/4Ldat1Ra5JR
NWqT0HxbxQO4AMY8I6VYgiRFvqS1RUadF3N79eAxsQg0MXw/yY3Qxs6e2DYt6pZxSmjSoQHz8woQ
zpJ3KFwF9yz7fYTVSjPZkqN3BZG7FRkrWUaMWxrr+eLJ0EcnCfqdpURbfHKqQap8cxrkJG1LEOHC
d4SncJGWkay7bcbx6Lq8TW9DIBVsv8bNUimXQIthz0hczDY6FyJkxxfiVA8NpSXylsEDULFB3VgW
52lz/ruBvhuWhVMiJfqADJvFC37dh8yeTwdWfXw/x5LOTKlakiWT4X4OPUc6Ok2s50QHTIZqhB2V
RiWfOYS5pGdYGasedK+A1hKp+T0F6ycLgNeSGzzlb2Quid64n9Flt2uOHEO245l1TLXb5E6fapgN
ExfavDW0GwmyCgpojlGDQ1Y5bpeI/MfzJlAXNnxwsrrrOPpnEMwqbcZn2jhjFRJ3V2DXXo1kdk/B
9B1GHX+wVfuWlG8C/0h6tPnW8F17c/aFhDPMviFNvyemEOTN1DB0P+edbcua0nMi72So5X4+lFwL
K/MgTUa8nZC1C5mJI7pDN6+Nr9K3vXXO24n+20HNVMXnMem6UkqfAd8eRyY/SlZsGrNuqKze0ZEN
GLq98aFGaPMnZdaUc3zFgxpG/7oLZz9EV04uClfOpZfDi2uhmdM5/zV3bzYvCZkHf8W+nNUrJFBf
dPom2upsolKKnTEDKYNrvL1wKXvNfBE+4DFATtiYMTrU/TSEksnn1tnZtRGNFIyT23p4XS6+SFTI
2HCWkbr96fFjf+I5i/yjGB1VPtRjyASSTxiQvKsyuBEVvuLYWjSlEYGJWa089Jdk6hXGFofIgvSJ
ceWygqbfuKxDLUS0h33S7fML8jBchuw+gVWzbves7IxFy+SRstBXHTrvYSE1L5/kjSHDC1zrv4Ia
7E9krIbZrIRjpVsei0ZLip6UIe7A1Nb7mOhmVan3MwjdX4cQWMo99oU/6TfZGFjP3u3/wuUWoIe3
N7pEZU2jB4K8TAzoPs45c1etj1i7HoWmRP40ABxjDomXC6pt0fP/Vl4beTALwB1vAdxBleUfiViI
AlJpZHrmVfK0G2/fER2LmQH606eq4XeeeM92BBrizqmt76KkEdSr7ofer8h8jfkpuh/F0nNmaCxr
yRM+jwSEj2bz6a8WVXk1t5JdsUsSqPG6WHk7jRneuSEaSP8sigxfQDuJfSp/K6FMie7uz7ocOzG1
NggJzFjKUbhTVUSb07w+DCl6avFen9CbIE6qCfn/XuuxfHNdlbFyWwKcApDui7zcPpjm6Cd7nfDn
DcKmWgsDvfzX+0AjUKSXSiwz9u1pLMnqSWWvx58ImBDxsHezLrXR8O3vGzQQ85y6A5uiZ/IVhROu
2zLdQwWXHTdTXCQ/hRd6zLFRrLZYDFkOL1l2z9Qr2oWAUQB3PhTwV0xdkXHdxWoesoncCh8ahKjC
kLgtIBHE++YRmGLbV45C2nn/q0PI7ZT3F4Bd0zoBcE3AMPa0da1hm4ogUG0ww+jl3EZ9tJIu/YMa
V9uAmZLa74ddch1lz9mBzc3t8dkdGDzV+JqMi2iBp8CE0vkW1Vkhz3jC4VePRUcgcF6ccwPpEADB
YPkVF2wBPpeBGAQhrdE365c5HhROsSWvfi+kIqZ6ihhI/T8ctM6rqsYrcTGqVE0TyLjyyEEMeEEX
5UfmMAaO3E3PDAr4TkTbmBaiaRxJgDKYA4R6pbphMQdNRHS2TGGJHxvV39l/dgd9jX5KxND6Gvwz
UagdPUGD78t9Ov1txglXFb2eRhkkTmCLFmfvxFPqGR5aN7rL88RuyscbyDuQs6W+F2P9mRHL7DwY
4Vge6f5StjZvsBpd7hbyeCHjf4TJK4dn4HrgEgoHWd8/XQfqrkunymL0f421kTUaG0A1RX4wAopB
1Vi5O2CAZMjkp6i+QuLYmlh6uzqauEVr3lx0UME4ohcy24hP1rU+dCKJy+vFXP1sKU6QKNWUCZFW
YSCz5A2on2wWlHm3ATo9pHX/utW4kdXWZBz4H6r8Ug4wA0bZ9Gg//tJmjuY12MnbAtc3d/vEaZJ6
eX+Po8eP/nHsnYuT0+f6+YKJEuzPHqCwbVdvmsdtMtJwCrITD6HI8SHJYTBlFB6rLpcujhdeKLKN
TvCr5lFZojmwE6+cDxWxaON61q1gslUvSiEEi1gF8RAAE7yEDaOsFSAxhqp4eNoKFZimL1YTWm9l
VBR3+GTyaBmzy3WI5z1yM3C437VJ54H0669MaOdCedIw/NOgCS+DiF0yjdGA17ZNC5mr8aEN00rN
VDF9T/F1NV4lfBJ7e017WMxqEMvuybdKo88+gapouDsbR3JI+ml3vouMRZKTQ8ervfQuWezgrYlJ
w0HFAd5hIgk3ewQuWbkGbZb8fX+XG24qsFuIMciNww2mwDDMgderBUIbMyTUktHjsDVioEbZ3Piu
lyvxGh5cDMRoR/2KVo0y5pgmE+bRy/Ql3Jher3ZiJDohVPI7bu7d4daNQNiwdnd3kT7sC1zqVq+6
IzjatW8E0XpmVlh19CV3Lx5R6wbBGTJoEfZkrKPcOO2yXRCTG99JXzxW/0mFLuNDukG3x04+yEfN
3qmocqspXMksEx0pW39S7/ddraEMn0EKsvlUF0Om0X9ZeoqyKboSe7DcuWMBIkoG2Rq7cZDwbPmB
Quw2NtQhTC2Z8fGZtLTD0BpFMYQpwFFJdrmMayJkiRQW/XkiXsTvXqQeQvNzYj0hb9W/9WY5TBsJ
EzQepS4RfHzQVwNNPTmFSb4NSUJ9MRmvl2dhp9X+pDTUM1SpfeDUc+pCUBF6uxGmjtGJth9N4zAr
KK4pl1aP0Gk8RvQfY4dyGPnZBBPmVVMinuCkqzmDFDfK8RZR+UEpr/VUaQdH7q7j4YriQ46bguqD
fqas1/o4WfxDzN4+zLNgssXcg1S+nB7N2Ep9qVL6sa89IqWj5JM8zHCUyR0FnJfOdnRYCR52ZzED
gqZK6zH+zuImJktQTA3uxq3CyZdLa5ePLw/NaQqPi3p+2nHyxJl4d/nkwrFt12MZks5Sx9eHxyiK
cuRYKRf4jhS4AoiZoyRvVL6cWfO7J7VUmau4BP0+Gt6MELASuMPqqVr5lFm6R8Nem72+lbbLwga3
vcRWHzg3zJnKV6GjtQsLQ08q3O55/ko2/efgabrzsJkiZPaYYXdovjCEDQLR6WGXGDptH7Mbm8UU
DWQdGzEnrYbAxRE+cY/szD4PaMC5YjGoyN19YyhAMRo7LpXpOVyGF+6s2bLXa/vjNX7F+XEg1e6g
gqW2cpZZ7b9Qb6VB32qDVgUlxZ7mXptlEUAwWmiKCK4CXRJGc8+VkiLKjP14hBe5fznCein80NdJ
r9nChrTaJnY7itRqjCqJvUhoKx2sXmmIbuEuX6sLJrF22dmiD3kyHZkXnidtRS41JoWT3W97/D0f
JF4lAjZug41HAsfp6klJoiGsFc1G1BbTfm3vaTxvCXcJQws1t58Ue8ljj5W0mHQv0+nXSfOnwQEd
tlQWUo0TBhVu9p3xFLOjHaqTZkkCGduUhqtgG5sZBboxMbCHqV//frFKJyKTI0swBVm8RgpHbe75
VNYbOOA2mr51MhYeUWZinv726h5xCrrNxoXjkB7YGiqCB6iAYbMgrC7e3yl8/vBNtNaDMJPnjO7m
uIbmroS5RA3du+vhC7LqNI5866pG7lMLKkg/+mwroaWGuryCBJbxc4SZmhX2sxhvEM2k9BViBoPN
wA7vi5b14QUHp/11QaCZk+ehBeHFebG3X/NTFRM5TLEFw91dXGWLFCbmJ4S5iW83scyPVH0TZshE
vlPb+jS+O5dHpQBx8ADtfQRus1wtewKz/yd9smdgkKOVMv8bOReXIl2dZYja7fBNK6ggqCZmZ33e
NGD5oYnUOpuCLf8Drh/qqcE64YMhDn00m+d3b7TejDMCa+QKhBkfw+ntLGhCYnULWLWvHjp2KF9R
2JYI+A3y69UHHfOEmoGGOO1wrrn1gFI4g29eBBhMfEYQFvzsPylSr7o3h7IFQYXGONhtBiX+IiR6
b+jHGeDbUpK2zLQREaR3ZbmY2kEWAFFOsMPGMmosIIMJ+UCfNCUd+EuDFNS6S8SeAVpuWzRIVBGr
ebo4T5aD8UcQqRZ7K+E5tG4qxY7g16KTkKnsz+Ax8mHypfQs51f4wiDOJJOz9BDr9/T5wXawnZjo
HwXmhrlKfoXS/2gLxROEUgNwvAGT0ghImZYsCf6Fa+4sT1Pn9oxaDRV7V9++kefZ0yPNvdhQEPEE
hx8mC7x3e0pbakpGjVI7tGDIikF6fWPV7I5JlBOgpagSYcTrOtsG2BFFjU9onKwUMFo4I/QUGQJ2
FZS7l/zRlhOFIIROxCA/1YvQKLRDN0siHcUL4RqArGUdBEiXOvPqlW4AjgMEGFo3DfzGQt+Ag7Qh
sCNMavyielWHTGSwXtMZPeXZd5fdAVML/4l38BJ2j79ki3Lz0C0keWTFOKhEXzdRZ0NhbPORAedN
CosF7V6E+wOhB40EzJsHk8CEjAKNXAONJ+J3PX4CW5j0ytjeEMpKyoEWBnB4iZ/hqrHqCSUQIPaC
eC5/8OQC35/jyED340XFXbOjPpwVZBqxI7uGJR67xDwUq1wP0czJrnl+pGCL05yddyrJfvqV/vlO
0AYDjQUP9pZVoCoi9cmZRV0IGVaReF93Upnqt2svhOqt1eQ2fPTp4c7AJx1llbLHQ8q4jFMWDkD1
n02BodMnLC1O1Ozrt8EX1QlGddwwc7ERFRO10cK86zxQvQYISC1H7Z+osrputZrqltvF81gye/26
foGedoc8kA8eBkPfl5SP/fmyFsEeEVBM0X8CMl+6j48QU8mYkcBAWglC/MkAlYBbOUqRUQbFwQmN
QJULbU4UuqavMOBKd2wXwnRLnc5/vL9F0Jhdb8RRL1oeCW4neA2T5XkcHQLhwNfd1TYwWGisR+6q
D8oc2t5tpw06/B9TvH9MXN9yFYF/huVH45kic2+K+JsPIVJZnqNYQVce8ySd7zn1oXhgXs8y2RPj
tz4cB/Ai2NqyThQOgBvhMU4FeRZs0rr32Uk/GDp4f5HQe7POww7e7oYgK/vcXtxG7wrWQXePvQdh
RXzj2boBPMVdbR2wsIl+rNfezWBhl9r0wbNmFPwz081TJYqAB5JlWcPsesoMcLpOLxMGjkorpqvU
3nB2FUX+YcV01IiGuxb8Pkvb4Go3hmFua8eO6iau7CYCt4zxzC8/g7jq4dblSJi6XqQU3a95yDal
3He9mwD+1Xw+aeFmBx9RFyuD9cRVsnG8tSi1bRJoL91UmaerOTx26Rm7K2a89EJuwEOSC8Sa5pWs
dU48Ukkx/GJilT68awuStM66yLISQKZ8LeE5fUOtK3iuWzYI7khRIzVRCOWFP+aBGCWY5Em9G6Mb
vm5Rkr5Vo3j6YfZOhj7GPrAaeo/BRKidIzsyLXSTgehclpSnFFf9f3XqHQ34jOg1pMkWC/4zEhTe
oLxmWZ3/P/MJCwDmCA8MBE4zC4e7vIAQqo611Gba3reF8/y1zz7hKQVYDcwwiyCThdtOa355owKn
vPU4RwlxafS/JTopeTWoxZ485NXZJpx9X8f0j94PXdGwtP5DG/O2Oh61pwE3tPafCJpBi9BUQsCs
hmeSMosGatRWub30j8Fyj7w8VVNbOVoLlNAl6DLHK4DwZ+YlXgIXZctyUgj/Ei94uNXBLL6wN+T2
47PlaLMug4NoykWjie2uZFJrEnkl2BgWpL0bYFDOXQedicKi6RKNq8x/ewvHwrYkqJ+5xsZUVsA6
G/1D8D+qLEVZ/RYUAYrRBvnO2GqcAdt5wFi9aGsvWqrT3ke/gb7N3alQhEI9FIDeebjYLYVKhhnV
sD7sWMGXB2y2pJaxzwhokEMiKh7ERV/ODW4mLT7eee0+yKAfJsPAdFs5T3TkugpIbaa0j2FhNHOM
3QNe5N4hTxJOgv4AgFV6HB6aHRrhIzU06YhMUpGrR/mK6yNgDAs62Q6NeCoBEnOf//KeXjJBUZeM
UFFS7ArKivC7w3mNCCLbfvHQG5dSEyp9pnN5IPzMLks944hNzYkfyaqJHi3A2zbO7zoauCb4UUD5
GpM/8Er7jVwvHBIGQBKt8u9AwxbU/jaxBh+zxTevKGgY7xBylKT0pi9xyenjjz2bMzKYi7H9XkzF
46f2q9MkQzi+FUIBmHFGHSWen54YHkeEF495wzuPshATAwXXLyftkW2j1ofYvHbAK6H85OIn5R4F
IjZ9B3mUFbhh0ipPC3njReIeNKgKBOx4Xk82LirxcYi9W/AHX4jbr5q4ZKtJ1kYj30pkEyq7Upa8
Ej8AytpjgmE8/bY8wBWJR5UwvMvad28uRBwgl9Eu43MzshWn6IGFFiQY8oR01/cqR8CqfP5jgxk2
LDvPYIfUIgGutDe7SVldQTwrZIlSyZ4gp5whItV0nwS4PNJfu0feOaam8dZu30vr1i18D8gQ+IYt
rHBtfChB2oT9DetJyUM/wgJmtH5t2Zwo+0Ir+JjdYjzSx3J2H42gPC5By1l/IkNHOC2E6+y8obKW
ALHDcZtzs3FFZOl/Ar1qpyOXrPqxCXfA5WwwcUl/C3TyFD4KiHddtcJjIEQz3Xi29DQ4Y2kjWr6r
o1t0j6FemocJ5oFPFWmGN77O30yqq0uQTtGg05NCWXY8ZdSh1djAG31DKo8mUj+EIYDo2bkhlz02
gBP9KTWRWgBmPOaFldDyfPzWL0yVTqW7a3mh7hu3+9GyY3z7sBHuSV/bHUl8EzSXayfy9bXzLLHu
bMjXMC0Iz9SMRHrC34tj87mWiZR9d5+eLJFiUcoV39OQ35irTU57XLZFVRsV5I17uwPaPnClRabY
83zNVxNUuZ6HjhnxMHd9DLd4wnYE22T78nqBafHh2qvd/lSZwaHmWNhp91Puv8esDt+L+Yn16spM
Q0cpmuycfpLH9EcRE+YKYtxJTIZKMecwev/cd71OCgOwohzz5XrAgDDIFzuRQp5r+LOB3oTBnZ2w
c+I38u2xkyGTu2432YcXU9SEO+w/ohVtRJwl3+TVpbQs88AeCPnW4ynFv+aQbPi0Jl/HxDwUMNt0
/r4lvQ49nr07PeT6Q6UZsL9lSWfeNzhLnY15WC5MlFBobiLmgi4iRWD7VzsOjk9jskGhPbxbSTzV
YwP9U1fTWcIX0AcXsPJMUXq4NQsMh9M4jbNCGoagO9x8Ojnl8g+H8SHkuIntyo042x5CWw+y/N2s
X0YHiGqTIbgnRdlw8K4AJVSOj00WAi9CF0Ja5Eigtgn3meCAYH5H2s60wTbIGj4jNP7rDGmpzkMv
Qpa/GRpRJ5QEquoNtZyT+CELTd/7scOWv5z+Ulu4FiKIAQzfkkFnLC3Fnb+G3i1RTlXXbKOrKze5
7tJHeglqRlZiPfsSzgZayChsa8997N2WLs8PkEBrS4sso5KfD7//69y9HSMng+xNmW0XQFxdA0rn
l1HTtqcWTemQd7tf6V/2+TsIPqQf+ETqhseIymlEyf5MCfl/Jv950orVwGxxs6kSUFUUOfBiG7TS
CTh5LRVWYVZdgi+4v/24UF0soVMVj/8cT9XhVL3HCp+SxtwQfL54DbpOftYawoQOT12xyj1q1gGm
9l0W/P+zCIlxT/a8tYAf64ujsbnamA0N0S0tS0k3rNc7fDcYCSukj/v/0sRoLDIfveKsZSIdHGrj
/WbJ4DU0GaIPf/nIKGFvBCVSiwdWrxG1VrZtRfggffImxNKUB84uX8vHRAqC+8MXrS43PDoIDeXC
OTyBZ9jiQuW2dWh5T5mp7Z6N+g/gXgt5P35NyoBLHxcjO+Cdz+5g+/UpV/O02jFjTuCQcKIOKpLe
R8V2Y+Jyh6zDz4s46hw34VkDqJ8tzKivMybaeSCYORoNPCjQTFJ513lE0qaFznXSSyoqH4cpSHV+
wL9P/z+HkhNaKlbMVQfkpIGpqwxS1Tzos7rtTqemrP5f3szQrG3ztJWhJwgkGjk6wmZ95gY7i1XL
Hdj8lD8q6iwCMckDdUo2qiDtigHNCBquPz6Q28IyHspEPqnuR3yQU+WZOQvz721ySLUdHH2rIFHb
rQFijjJzzfTVbkCwzPXnyW/XO0nCPJXxdCFLPRJJwKSTdrt1ZxkDtz3tYJ+Mj1TGjePSNgrdaUFM
FohAK1xby8HARpFu8mtZHRqdr1/vHc/iXsUQiQia4CD8n5QEmn5vXvwODPKonS1YRvmAJUPhYdbx
3tJrHrp51lmv8lyMEqWyhVDTSOhoShbmDw6+PiJtgoUU460RJK89DNLn3cfgwCSwccZW0lAmlC4L
u49dWB14FohldmYjrLRZHwIZRkdOD6YIdR3lRRLzllz41gl4L9BM6G/EEautvz0yBFN1oqzxOODA
nU7PGqOYR7e7Vm0eKIqaaaFAg1S+7JgHPqm/xEgqKM9QJ5ANjSmcRakgtmem5w1OqPbPrCd3AEfe
ANZ/eg1fRGvS1Z9VbwlxrmhuK+27wRrlJE2LDCrYvZnskfvHrFTkr2wXmVed6lcuY45F0hUhIEAF
x90vHL2MzSr1FS1gPS5n7Utm4U0ce/pXjj3F4Ys1SyJJZrJ1Wsdtn8kel//CSyyH7mBqBHyBvLTc
igJH3Vy6IZ02doqZ/tAhHB5CeAu0qLxp2XYnZgUKk2al0Spdt7r5YOkNGvYJORU7Qe0XyEgRc6d2
G30voWJaPs+eIrjofv7n5pw7t6N49HQK00qDpJIcC2YXOWQU/Bv/au6KKQXyk/uhIVvuAOWY36rr
LYE1hYlCEh4xM37rSvdvUkiCto4ecc+BksDvlL6/RFNep0qIG+n+lknHUVH+ulvvbBk/oHsPTn6A
o1P3XgEMjphrDDWe3L1YpviKYHPVAOuqHl/iMb3A0uyXiOHxvBrh3Lg+kvWRF5U30vHHLCFwohbm
jes4EWE4B+BLfxtza0udOrHmnaL4VJdv71JTc6GtRBqWe2xY4S3WvqYTO5l6dAfWOg4/L4cNBmZs
tjnjkMO5gheAvmLyd8HaGjkfM/xbTG7HrZRSU81+DUkh6SxemVUC1WMz0eDZF3nWQFb6y4sdiqKt
QheCY2855UCitHLrIjvW+Hd4brOdwqHlfhZPxG0jPb8aOLdPn1vOUfYPLopnokAcw2v/s8LCZvFn
s5gaOwB1LAitZbJBwjyLXcYpvx7fZQO3jf16gVAv9jbAJT5PqCYiAC1B0jD+zigS+YbzaoUekjsi
lvmPntKnty/U/NBDgl4Atp0aknidKB9O3Q/u6x+C0NUOchVyBLqK6TVDeVIQ1oM3W4MenZN4Jhoz
3yoh2QwW/6nTJYIxSJx4yRrhy3srj2/I1ZPdDAOvTFArPDNtn9Y+AqUAc9nv8nTGoAtmzopxIP4D
ouT8mMe6tKjn5AA5I/n5deDjOs6zaAdlhRtCwKFboS2uIxAfp0bs0P4u53E239IQJ3voNdBrkNoB
/BP7buVF0mZUFA/Ti8tC/wXJumtlVg2v/iSYCQ4NlicxFs/y2A7g8zlHcWFjytpQEkNp3wpmD2p3
AXLfEGUWUfnOOrZiJIe0QUuBjJRWct9tYITFGFnSNdWmVizuInscMBiii4dbSoPaFi/DrGNRvoz0
DtdyWSdR7oIkIP1zgT8BwdYNw2Pu6b0fT14n8fmnACqr9UnVWdd+B+dtwq7WgOAVX4SaAx1fPszV
6Y80dM4SLguSLy0hZdE6G6pDVaX50WPK8sM3CZHMWQXrF9ISRNVfRg3/1PToVNouC+YWZHf7GMY6
n7aff+/cUyk55AbPJZ59a2b/+xWGE0rZKRftHTypAiw6US31mYv3wSUtMomIrrE9YbycE+f/KnNc
Chcm3MFPyNdNn12rK7TWv+OXM08wyyEIGGqh0CAKOKWnUgRZmcUu5zMubxza1XXlKCw0v5rfpNlW
NWsTCKsAplMwJ9EoMaKTU0XHx8uf6MJPXTWCYPGvcHv42q0m5B7ZMewGYOx1FVOLvR7EQTxUNqqG
yLXM0HlNLvYy1VCHFA2e2vzDVNNy5q0ocJO73ClxZw+gXjeIfrl4rmQVziBW2FZN0Gw0Ipyq9f73
1XVBRcXyYGl8c6aPB1xA2cEiFnU/LJs76uLiB4SZ7JPb2K+XNyhLvdCcO8l0OMWqSY2o1dyxHeYD
vA5+B7xI/VsbSLIwf7KoU8JkhZXWDqn+lYhGGNwq0aOHRhBWWKsOWa7F9tm/dg7jHqQCtJhx/X5c
3yi2dx1aOvfSH+VWm0icK4a/d9lf7aD/y2gfGaYEIHWGwfgNadwm/d3s7zfd2EUCdviHMAp6G08K
YPd2hG+UlHwH/I/l1xZ96JpBeIZcH9IPfn/bt4LM9ONr1C852U+In4HQOIRG5dGlGpIvdpfjU1z2
cmIizW5O25s5N7ImTJzaqZZF6rjKjrNWGHiP1Idkv7kMF5+kB6N3aY8uuxVXYepK7IXIFvtrVNd6
th5C/w/vKVwrsyQKc5eAcahcgQ3B9+kBh07XWGzMrSWth4tUG/ObCHXRYw/+8GRsdN7F2UV65pjY
K9054OSh8iorQ9raSWOq2GiJQf9oYbV/xFFvOhxINYfsIyAlXnGvoW/wC7YcRejeOwgFC0fkjmeu
8TRcJFiKf+DPRssCMWWBQSxC2p6xPNCF2XgTP6rnFAMF3RMb1heYQFEnYdyFWVyGpQWXPHprmOyC
WmGVSbJkh9d8tftss5OvsCEiw+JI4jylU4qpMtlteBHgJVww9wVl9evp3p+KD/R7zmX7C1H3vRdN
poNYkGMpEB8bg4Gn/hu/hHhacvaFDJQPrS6c2RK4JYXLZccHLuw6Sh04wlFqPxg8H042niMFBa68
2uLBKEIW3e+nhFPpD0XbtQgT0f3a2fQ0x2whlik1Q0D6IHEbd+Z2qpNwE5iSgG+H++JaklqF9qQi
N7pQeGq9ksvPmotYYLULbfhP8MPvj7G5U4+nHOPwRFUfhIKYXT/u1+ZhGoF+e+ts8e3K9zHeFHUO
4wF3LXi2idNkG9C+Q3qUuzZonc3CQ+BwEVNVSCxMRblCSZa6KGvCWsld2E7Po41FwgiJza1ruY5r
xMHxJkpKBzBSk+MGDrenYJZJM7SlD7qb7CK1f/hsGUlzpxoDX3A5ZleWrh/HS7XSVnnQUvWbKcWo
TypGH7qrUyFwlO5Boe2qrFFkg8QOVy/0MfN3rdlKVtwt1/lGTh2Rzhr7GttdQpiH/dgPx1AQHy44
raU9sAoWVlVeAbGxRA9wPnwNK3E+xtz94Yl5QodWYQIhr+JP3DNWzrAgnpAc1lkOStj2MA7Levdv
XvSsct0XijfAooCjf67CvffqK3C0kGqr96u2c7BO67K70LYqhibRIoBFIBi5vDJiy2rELY7hFNYs
rN4thuBlYLvVPs68qzHvYt8e6xlhBrP7gc1dIUlBfAOZ55xy24H1vo8s1cJrXNRtUnoqg++EvuBF
DsLl2slGSNaXBY3IVWgdgH6QWYXepTyng8ETl7zl2nPBofiOIaLXtfdDKjL71zAL+EqGmb/zIQ9m
gPrSewb72/Q18ul7iiy5JqzxrhzAHsmALR7IMkw3LapMEGzh6h1Ic8hBWgJlqQhU88Lz3j+uNgJI
26PxsiHRr2xlnCljdr3FvafpmQOEZ08nG+bWgpYEMA88BnYwjw4Y1FNLqabQH3Z2+QQU1JFN0oeY
qcPMRl7O4Rr1rXKCiyw/qNWTigFSKKPuCCM9qgvb5s+hqJdllqPlvZ+dVSUGRyQh7qncV3eC84eC
TIaajFaNVHOhojwzyw9NFA9EfoqIGz52TxhkvqIOBoGzumrTQBCRB/ZS74MlXb55DFRR7Iuiny5U
Fuhk1zyKDraZU63FgAqCvQcQyBLXME11hHMDtz+XAE8jx6ulegRzD0OO8dUBaNcyQNw9vlSGaBDy
s9G8pQLtYGDhsAE08gYClDsyKAQ/2HQq/WXm7T21HPUR9G3mCo5hghyUqyP/aYQ1i0VLfIlAlxF3
54OMjT5tDTtlH1snmgHWES7N27JsmTEj5T+V+oiYGFVbPa/8GreQ7nX0cOrn9l8hNJ4NK9yNCgly
mRSuFMhKx0EwrvkP9vuU86nLJNsjnvegBHNCk33t05kSTZNF6VKYDNmIgDeO1YzEaGup85k69t9V
BCFFVA/WcGoUXiD2E2faQO4PVMuVtu/Go9UbCD93P4Mtj0k1Tk34zELFhqeCiPaZSosJ57ouGDEi
lMa/K0EkD6j0Jb5MyL1iSk7HzUWfdPG+U7ksrjjjO4ig5zvPs73T+XGR/kzrGcL7E6tdC3yzjQbB
1RhvA/0IY21+4tZk2wJaY65Y3AvPnQmvJ7vS/NGBshmxZLytI9PJjBk9GJ8pnZ8qphlDfvAf+Bet
+kkU0/IlER8l5LQxwYNBECe57+Mb7TvT8Vn2UdM27PQvdEoTPFZtMRXjcy1NnAMy1lzEh7QrZHDJ
CpMYXrciDJF0a3PGEJ9QfHIJc3D/QSUWYUbRlkfZ3mftlZYzndT/i5BcsacUB5sbG/FWuKRGXV3J
CZ3XQPtQaV8+/XaZjJvSyh9sVhIvsW/Bzvw0SIDiIsSn8ePbWbQOeQnX/WWzmzBKKujkpvl9oerO
QZegouyUkZeYvNcok17+H8vzCcFfbN+L25NMsaIMGsLhkmA8NQ6u2RTdbmlFz0S0cp6TiYf9GS8y
U/fnw5E9qG1lft1Q7ElO8o93YQ5lNfXGV1TodXZmhnDKX2+IEM8/y64xiAFzTg9RVj1ga7/Emdwb
VuknYmdC40YJPSbmfhM5QyxThZ4MmBAxxWCqmlWw4OpsB12zf0MAepzRkuPo9+uUtHuxoiqQsnx5
dZLm7ZNhgO9zADbD13EgDrEhwJaHg1QhTLBhND7hwj23qN/P6J4mnYzob+Ih42VdpnQZGIj4wEov
6Po+NrvVj7XEpqUq0dx6XIL/f3ZERJRXaZ/ucpOB6vl34clU2qspSK2ldlNegkexCm7IdiRSMK+u
2TYsMrQy8MEuX2PLP6BJo0s6kib+xdklotr3ByC8AdMu6kuynNDYeJh6sTbhS8ZwZaSG+xQo1Uk6
4g42qgaxXGL1mwAeCMcc7lc23Ctj/EgHnfKA3z3CxADL0yfYMemuLdFHWQvJ8tBiyleQvCD1/HWm
38q8v7jvkkJRO9aZESVQRP4hqznaWLsB7G3bYCkWUW6qsfH4iQKn0skbQ4HlYrgWfN8eWaXxA5wi
1bTnmR/Ifmp60XpLrLBmDPlkKftoVmPAgNgUkkr0iBVVsHQJPKZno2TDQJxjB0NSxPQyjh/mL0m8
e+dWRnu7QxJMz7ns0vdHHzkhD5SgNJtsucm3M34NGhqDMC4yuWZ1wmrJ0ePKqEFoD6+ZU1IC3ehM
2BDLRiM7bEaiVjX/0vMg3w+lq+5ixC8wSQJP/QfGUVWS2zRZqfLLBecBI6ycvG7XSnIU+rmYjTmZ
E2i1cvCqtAiyr91nCbeEdD9431TzM7KoE3aZi4BrbMfcKUDviasOByKHQbeyVLkubMhKyRVKc22f
oS0WPxI7GyrH3BfHzSlp3g6bZMH14FVv+x/MLsnbdZlM1Dk6/CktjlcCd/DcMvkyneUKhXY+mRUb
Zjuyox7xsTiWMVQJwZ5xXfbze/TR4fMZ5mvvgE2tAQzHRTIS5xeNxADGeY2YbjEuQiA8ar3iVZHU
l81TZcjVREZ/MZVOk1iAAAXrRjv5PrEQoiuUmpfe57ohQgHh4pUkuVhuq10zmgjVPtjiZI8oq68s
D/THc4+BR3kt3PDZ/yfXsjm3KE/OJaQkgxofQ1xrd1xDZaU8064EigTDegtkMOmzidxrjVKj2B2s
yRiHX95QevCzcddU0cBECo3GDv0hCz3Im6ZMTMzxH+kK2WrK7WdPV00PXqVJhV7dKFdIEbBoUHmS
HUaOmRBWBixxnUoNTJ/VJW1wqDZ36ZlD8SOuqO9VlGz6TsrzfWuK8NreH7yXKdPwvz+WxACbN6me
GeQ/0g9FewdUF+T172cIYEtQUOzTmqUZprXcOlGRCDw44kTGmeAmUur4yvJDrX03DmJQkF5jF3as
+RSYQ1Nsh988sqRSoSettAayYHWtRs9kxLXOvpUrnYa+8+mplzLPiEZdpgs1f3c3u01ogfnZbiVo
RiJEOb/e/cavPi8jaR6z6rjLbKM8RDAVCVnOFsJkHuUp+bbpRKFTcQLbt9ZXEwFFflAq/EWtLVwg
8sirWnbstFTur3rbNimLo8/I2r71uCWM19MsLzSSVNlkqBQePB8GylbZ4gIL43soxYk/R+t3uV7a
a843dSZWJiIA6218JtyiiP5bkdJJlpiKSJbuwzzDu7eDRwAdNumc4bZhpXAunOd+RQiOMBQsM1U2
6255lqLI/g0Dl8pUwhSqCoeUPkAP/KraRAdjb4M/Jm537iEN0sXwGIwU0tWOH7CGKwijmohFAric
GMNOxjjdeorVMQlsBSQbLvQJa2GAhB+3/AmJwVOg4UJ9q5VxerGn+2/z0dtwsEhovrziUDuJRgQn
pKDutbBYNkVMAhSo033T3p5L+Gl5ffpqxI+uSKh1eyefSRZ/Wz54l1Ky3EDaAg6HcmW/9Px+HElh
faY2r/Ufyx4bQjkdJhtZcbM6A4XmlnatDd9W+f5Z0Q7V0A0IKCTprK4JvKdIy4Teg/Aj3AITXaSo
ta/TxBPnR3Zy/DFjnUVMofBz6NS8XerjvdItyd73crs9EY0GQQLIh4El4OsyiXkfs5bgHrLi9igZ
Uw2JH1475LUJ4Z6ulBUDtTIda0xoiz123LpH5jIDHey36IDNbvNLEJlnJonURUin/LIYYZS7a6IL
Z8WXx7dWDuyENvFSG1oPuTt4pbM7cyeuThRLy52mHUF+vCtkxPhnpGpQT9ebt6axelc+qBpcmE6J
RlasPY/mOuAbusZabIAQnpBso6/t8yINg4HjbjoCt+sWQ7XOBhuHJyGOFRTNOdQVyJ8/kD4Zk0hG
GRs4je25IJ2ytgSxwx6QY9svGNEaYqT+VooSceu51ZOPY2r5jqlRPKqucGTDQYm1m4eTmHtGEIDb
tBeUSlgOlqwWJ11dGU5Ru3fOGZY2fIEgE3Se70et8F+9mOm4ldPWiFLibkL/QkgQmyc/Lg5sAJWB
m4ZUgn0PDUxjT5C+8xD9JTK33g7181vpXeqS0fjNjyuGuTIWNSfZvO75joujK+NnjyNc32AGqZ5h
OruRfZ1bhQ7OXv1cmzM3br6yQrWC0kqyf/pAThYMHjVaefvI0PE8x6s9lqmPX1V9XKOAUDGGp9P5
iztngMkZK5j6shwU5ZuxQsKsxJ3rmuIiI4zpeiAOWy0kuZzq7f1z6UgFygOkVsU3gEjE1nLxFaZa
Keg/biTexd328DeehEfWVH9U3HcVavIrM5amSu4GJ1JNsQ6HJx1m82d1/23TuF7ZIbftdAlMbKFH
58CHgBa8mfYiRq/0JQrfTlK4izQqK00jTL9LdxEs8nfbyBjPwkLbBNh7aZXC2aNUetq2H4Jl+ZW3
EF8IjGspDZAq3FrWdgRdQxgiSmFACLi82o1q0WjquKjLU9YH6905T3adsTQbc1jOWLddLeBJ/zIc
DGHRsevzPU52RpopwbdeTbTT4FRPmjmgiw+eFMDxFOuLTLHHKJGZ4cMQ380n4IZJKhbTjoYm0oL5
Tuh31FjQJzKASs0VMqMRLoY2/adumRqqcJH+L+OR5uAis1YqBX7k2heI56bPsSapPVXq/Mb4HdjK
/eKQjqhvzRo2cAscqd3EXhxML5qfezoLSsfP/C7tTpvmJYFYUsSblQ6XGrvS/VA9LKYmMRImljHv
DI/IyCjfmbL7vnNuu9DIz6nqL3cRMlJ+tKkBoxnkg2gMhb5sKjRSJ/JZ4gmJ05Ef9l7mvbhqzBsg
q6biOclXaFm2N6HZKLKDmB4I/VII9WJndyjYswl1uLt0fHclNwIPda1WeU3yjj57kju80b16ezqA
HaVdNIzb57pk+Dyc54kN9fVba3tIUVdjQgmQ1O+lC3094Jb4nSfL19pPu0vmaXAsMV3bIExVc0SO
58HraKW1IciNQ3+LHEvg9NX9+8zIQtO+/87FXMmovfBEv5AHr+fh6sjsvmrDZc3jCQXK69RUDePE
nFSSSI39BzeW8YVjQlop7z33TS75ek5h0JsjF7Kkj4615Y34BxeEQdbgn1uiSULDSHPu7u6GonUY
W9MO8q7NRQ3o9XottczwJCtvlEmmTQuKZ/ypekYSrkijmJ4yXA+abE8jQp6n+UqrWrnlIqdEWlwN
rx20kMgLrUvFBnTnEoBNrfIKv5AhKYDsxgB4CiJbrFmkV+SEP4W5gyyp1YFIZXxOwnBKH07PIDZi
KgZdOuDJG5KJHqN+LGXdu3eIUEkBQWx2BvdR2302WbXYZnUlr7IuctLkHS//QLtO9JcLnk2z4FxR
BBgKl2aY5zdeVnm+refI4noxj0+8toTjw1y+gcGb4kRalgllyNiesrvUz5KZjtxST6DrJ7PRR1vp
OYXEs5W+lkMxyhNOM+o/6N1Xe/RMDaYbd1lkJ6LUTr4mZ7PpmUbh+uyoJk+TTzaLIj34pvdZ+OWk
nCgZHbISKV4OtR7dVBrBfozuNBDgpcDDvpFi9K5eo476E7kYlw6U+/UYUtMQ/GNqJ3wS5reCOyY1
KfGP3EmukWQeYfwfOZHqUjSa/Mr0InOquPR0nudsrfQLgVEg0u01VWkDUJ6kUsE+CaHAgwFUJZO8
j9kHfP4ovzqViC/2K0c7RTnLY2IkIFUBoD2MT499Aqi8Icmp89YtYXLkFQ6qBXoN0yzjM2om04UU
+p1J9Lftu87Rk3NgECIWHIh4EDOERB6l1coFD1qog2VlyhRkZe7mp/tC65R0MbZxKYcwv6zY/fMA
M4Qn0KPVezHfDBLz/AgJL/H/hU2vLwt54e2yY0OMfbWVs0DnblIbAT5qYxhZFtvP/JbP9v05osBt
exM/QW4C9ahiil+yvJGuTj8yN5CLXr+BloknfZ2wB7jg1Irpv/aHJWGk7fQEHze2scJauYEHe9zk
CzR1KXjLuD9MAC2e+NZUMklWFEX17LYhiCjq0qowGsU128feV7FJQVLKfg/DS91zbjAG9ulV6xf1
yta5IoKpOVphZuR10LDdoU+KLEEvevveypWcXmSIr86y8QC6KemmyRV5iRs+VKy9iJ+9bRwlZFjO
N5eiEuAKT8ehAMj7fsYMlHHH7LcZxtuU7M/LW7OtpMVR/EzjC+huu3oT3YwOawW5WhAJ3EEXgWv1
sxFfvawMj4WH1hzq5yonmtuQIil9ZkvZKvxJcFjjxyYmLUqRggRCA7IZ2L6w3lTfj1g/EB+nUnnw
6ApfH8Dmd23Jg8Xpbbt3nqFmshcyTHCLkJQStyM7vHhD9RWj+yYOeZhXMRV0BKr/QKWzBXFJjnjC
ToWoQGgsfaJWlccZClL8wGkCbkBmGxXMXhldwtDB108gcCSs4QNqE8ayop1oXYnXRofP6mJ7KNxH
jcVa3Bv5nqVARmDUBYCs5QeA+eMG4FU4KpkA639xmqDHDlgiTe9HuwIHm0yj+44O7sDraIzkV+zO
UwthRCSqZLI7f2j20Pzmbjc7qs+UpMB8v0gHZDVluGcmXiHFOxpq719CXeoTe3a5V+FRkXi9B5dI
qPhLBeofvCV8XS+lqJkVV3c6KFyDG19dkMwVAO8UqzR9eEeYPatGyo9KpRxux3b/7iLce9q/uC35
oAEK+EOwUPiXB9EXfGE0BGaF65DhZJocxhBXW5fA23rxXtR2XdVQtPN+VQivhhc8+6IkyIbtTc6y
8s6f6tZz8ujAkZ/+XzsizBpBGu3eAda5XjUV6F8HNnLIV5SRbO2w4Shn6+/5GdoYjhZTkOhL5a58
DzLWr4RM3aN9lgFRM3BluxhOleUAr/rTo03xBMoG34+Au1YyNGj+6zHh1SBwP8qRkDVAXnOuviHw
b2ECQcs4dK1COvaOLZUkl/FypCrRKc5PfIgj86WnnEqjbeHGvvBNV0Wv3uBAQA5uD1uPUqB7zaHb
OzIQHTlWeWgQsGdWkIwGd4MznO2B9inubRV7hEKmfhpVJLu/iFLiMZkA5WmnKqKTueQXTWsKw2uM
CBO9nwhKMWexAnq6b0SGj4u/6GxdgEliHsvcltcVMPibu2S4e8mB8dxOJ1FZG3rohGMobl+lQqSm
7+PDOfLuT/ptpuST+1TtDPeCdGoELoBQuJ/S3oFg4CH4/OZ8SCV4Xx76qkfIvkqSvyZvBJv4aFN3
pUkLDg+aPp7sr34gkZzAqASBRi183KZAYQ6vknOyMuCjoLT75vimjZLS7MBXq7FOrdfRTiv3cODz
5H19w0ihieu+gNwXY4l1+eCIbNRLbIlwRxc4QaH66fuEOyNmQbclIaj4Pn5F4yOMBT7ullUzzIKN
azcKZc3prYaaoQ983lvJhjGDZ4etzQfZ2c1ASqHSArgbIBYApb3IgiGj8QY6jLDVCxOVXxNPPNT8
gwVFR+BTWwudo5XrRBXZ4xxJek70cwZTKDgSpnS9ijCNCM6Fz8Yiquz2+nosp5vDJqjiN2GFF9C2
HuJU+pQwP3eS46DQziEUifSTsN6+YEHGOaArZgTQ8nnlYfGSTVazZGLCfHxNI+wkSPPD78QhL7Mt
yUYCXEroTdQvRvmPPyDP0+NQfgGvWx7OG6nwtWziRTX5rLzF2tbXHJQRK8WZcu7c5ZnFfaGSgZKP
mN6MazFmwkQoi56x2TUSSioQlx0+squP9M9+cOx5lZ/2uKBLSXBrAcS9mNc1cWfWR5/C6e4QFLWe
AkMJGvxFNXbF9UwV7xwjuIDXu42XI8Voxm9ECR+mPD2YS61l7TFRcijR/QZdPPfu2FrTFowMmYW7
P2e8otEWqdbmzGQ0t3kj0Mxy1X4FK75pbL8ZDu65qhLm//9vQTgdUcbzAiDrHM/QSG4EPX8Nj0Gs
aTgztfhXBUA9nzLbKq9PcYJb15348ifdS0fa8zG98HZZFINFrdoQXrkSCLlTrGbSl9TFgcJ39Zrs
Mn55adDz5coGvrj0yJRKn6qtyngB+MhpjoOES1prTDT+UXN5hgQ9fqLexo5RjJ9ztpl1AjB0zcK/
jU0bVVI5Q5L5dp4mQ2RUetLkJCxN5V5EyEKbck77dfoF9MCqcjifR9v7SIRCbxElhyU9y6YABgsW
k+ZGX9KY3ESPcZy7faQelEp0GE6wvT4SgHS/bkRM3a8UgF3oKkdrtXtKHKx/ncLSfItVqLw3L+tZ
bdaeYbSZb5IHCDKOczpRrzT5v+DSg0qFkLlSHAdLJhxbaZUoE2pv4vZ3k5b6bEx+RNWDv6eST2uS
H3xmURuVRRjVXF5fooG6zJ/hvP/yj6bQEvvMCjTWtb7mKKO+eVLTE8M1yVLkInletPYnilz5wiaC
akM7VVjoQReRmpg63vE2eRB/brXINoedPrg5C35mVbxL4BOzv+79g8aLxjZNVF574jBIiz8rZdnP
FYSp7JcGuq84v9ed7lSNzGd/5KqkG/eWkaa4AOpYF0+bTK66U/2bVFkCCeLTSaUfcENcWdrBkN9e
UfhbTMWGQfFIm8Di6n6/rdFHRwpKDCa5PeDg8ot1YnH63qbTe/aVi+gf9D+d7HCe6e1n9vTl+CjB
Rq2K8nUSUISz0HHPBHStxr+NpVJYqQ0SgAWbOR2ilYsBt+0apm5bfODI3fQXCYZ9DA+6BwrLWVk3
16/JEIDwX6pkiAj4dAhJ0nEbJ4wJfuw4I7VGckwiypuHwPqDlPbQx1ovURWIvItIG0fqvNnrYHlO
BEM+JmyfwZdgj0JUcBDe4+1SXR7cZIYQNnhVMgQ8c/MK+r54FzugRgm1eedgj1DyELHK4lY/PNQF
ZiVH8bsOKOEUK+MGA18egLxWTyXthdLpQKujp274G3DQXP2pC7piXrEVGy23pQHIwq9iRlnTXCCC
LkhLGneSsHIgjgJFt8U5U3a2nOraXuREWGGQKvIWcNbRV4G3geN7Y1XN/3CW2FI+I3olt3DZCJL0
cZRTZCF5Y92Oka3gXdx63geNSW06DXNGAlkG69iK1EVHbnnMZgDITp7cRlO2UDmrNJhtmGBeJzCk
OlLYlNlvG+9+lQyoAZV1pFQJvRTaPVZWda4A14JgexdoLd6Frh5l+FO8RMg5xTA7D0f3E9HS/S8U
vjJIBswvIA7VO5D7QDkLpdB0xuu7vn0LYWHw89Dz3IFhLecCszxLUd3YJVBc2pgn4b8dXcs+my0R
PpYz56O0PbEUh8dJFCuS2lowuXYk2ppy2SPvHS8sW3VJGF201MKO7031ijBNe6p0Rc/+4Bbsuj5b
gTgmrZloqa5VaedMY8WQ5aFv0AdMZ+GVmBWNKPVZ5aZipmVvLEHrYy5exGoMoGGM+pWGQvK6rTNw
fOyphD7YkpHiUQFQDZLtD+oS3B4bWWy2j1iXxo0YdeHwF2PCRQcp6JpvFzXgifEIKsvncsWb+Ako
UjuWYD9J3uoWsUC38d7n3zPPTUbNJB2NGtRzW2967lFI/Qo5d33LCU0cjb3+qZgDyMvQcqtJ7i4q
anplmiRSlaaljNC/J7Y55+94CDdcgCfIcp5O//gXxF5fgwFl6GB4TxxesN+K3Y6WR2aAiZ/57QA3
Leya+uulZz4hjPpYdIltK6kEKhdmGdoqYMYZbQ2erjd07fTiyrxcpNTWqJgXBtpEiN16OIcdxSEP
cYRHlrA3sPr2/+EffPAH1lbixapQUHuEnfP+pSryZTlSTcbWhHn7Iaad9Q4/mkWtSMARo4TrexqH
G+WCgyS4KHjaXsI/ilztOAV96+1R0PaiXY72d0tVrP6Ap/G9pv6rxu4WMr3SCelYgty4szP/YyS/
m8iTyb045adtayI3OlGVQsNE+VCQ5vhs/nG827CXGPElUkoQkZzZrsNT0KBM2beIAuiU8x8IhnSu
dLH95C7pBvDVnrUzC3fPphtWcoZ0FMqua8N1NsgPKMjo06TDSM1syUr/uOLI5BBY397FPq4bJ80d
+ICsv2xiXFgZwxaGgPswkfDc6VEL6weS8nSx/eKu6DRaxqLq2gJowmY26PaMaUCm/LFGM0RJhaH+
N0xI0kgj0NNMnczr7KV1VLv2Rf/6lqQRG+V2meUaC8LjbkwRGBnix8kv8lRwKc+t5ZRHSJMC4nc4
TsSKLQXb5OjBz4VYL+rMwaJJ86RQGm05MTZhMyLrwj8s8KxmztUfvmeXVS78smCxGRIGEMcsqEuW
c97s9WGKWK1VvcdCU92oVQYBDPZX9M1+oR/nhBNjhqR6w0baKqn9uVH/7WSL2FBW3JlTkbtd3JPq
4mIA6tFKqSCnVMvmbEfscnea6oN5R3uhqaiVkJf/JackZIK843B3EzP71oWgV+4qhd+gSzNLKuJD
4uivRaEoVmad6baek3xYN0hA3MUd5nbYTEVEykOLczaF58KUHUVpbSpeRnFRwP41ketLWtlHd4/e
oUVDRsO7SSbToz1yr/VhqaU7RCp6mwAq1ODjvxyH0XDH8XI0ovusn0MenYwxYdEJ+A/XIHTjLMLH
EDmPRMGCAM/Az53b34cLkiKccaGcOgsdVUh1kl/zcZpzzBt+3Q3fy5C/Wh/6i4edXspilUDgkOx+
baF/S+uupsuBnWFIqjYUPGM80mE4v3/xEQnRYnMTc/8IjZLY+ypfkWBS954UB00JK7ipdHCGp0cx
Xn0KZmpPRKxNrrxkWpZlW1cRieNsV4LYzKznfJT82EFZzbAzlIcDvItSkHtKo1mv+4o2QW9ZOoQr
wNgHlJ7odNRWj8lapGyOrLjX5vPYxKepi4eRdmn020uldn5sEjgOCxnguiOL1S7zfFu/RkgQulaX
yYWQ0kfoRNOEKzJbn9cIXnQntvQQZ6hO/zkytRtR7ycVSNi8a0T2Aezt3YGqJWC9gQP5xvrCCsTn
ZXxftse4JgYvb1aG0kR3g7+s/2W6ouxn0TCZHoWx4LKYXNplflu1JC5gbdN9pClbbROiskt9DwAi
FE+sB3j+vlHKy/dAX5qFC/PRrpiP2CNfa6JiPiJZw6sYOvwRxxwvP/FwYtKp0DojoTZNiM3Sv9nw
7zwi1/3kesoouWzejQiJw6amI+BIl8mU1qtv+/ZkeEKNm2zJl7Gbvap5MMjDhNvTLk1SEM7JSkZM
VC5yNSgogHAZyabza9uFhg+D+jR4asORahQFpse5KdSvHiSt5x4Pv1zuQFugRS+lp/2T4CskcV4G
Qo8ayoVv5R8vydHy6ZwiQiPOTrVVrrFZ72v9p26oY1YL3G6cS4DVGtd8zhdqFyGMpXZV4uUYfiz6
jZl7bJdNo/V8B3G7uLyP69XIh3BqenrwTZneNVTmCioiq21otOfpELxewTeJmQPl5TqFOsdZAyan
MyrjMNJaMGl8PESeubdrcdhb4pz81CciSnw+YgVOy+UOYkWfezwhBFop8O9j7BqFil1RaRjTL7bp
EFKw5NVuGCg2+FyL1PicqvEvfkKiHmI/AOHaXQSG4sQqW+5FnwE9TYPyzGmvV8SwNQMjbS7HNxST
JYOw7dA7fV8BIvmYqEVtuenwU14aoXvI/5+6VEIbE/EJfkvN3esP85zuDLIw/W0upqfH7hB1Zyng
YTOtTJbATBrpJFDUV2FSOm3rm9d2YMF5OMcLQHbRSmCQI3Q243KgN17x3LBktnv5J7XPCCnpxIWI
easgaBuUXFx4oarXaXb9aF9G5wM7EhpYG0F+JTywJfOOtz0paK4JFy7eVNe7jvUg8kOEbzvdmdaZ
2VGPpNO/GleUMoYD6uBU3/EQQscui1xcDnF+DSJZQDG6WE5X9dqOKo79y7UEBXTx1wgDGHOKMn5r
ikTmLI1XMNIPgAa2xOMP04O+3Be5Cb+LMwJ20yO2PBI/EjIoNKhJq4yDxEiroyMKJFrQxSoipjg7
CmX3ZJhr8oUo5wRn8DfDpkIhY3+EjNhDzZyDuSan4Vu9i9FJByZBS4weigums6y+Jf6Coz//+koS
Au96InHe0bYf9k66GzBxZlTbl5Gw52JrG792XrfGQX1JpfdkWMgqazsDL2j2qu6ttqQwz7aQq6jH
a7yZuRFxE52IaADiJrRGburWl49A64t339WOsVwe+IJa9gQCQYoTA4xi9ag+ffsXMjdRYCcVQU8R
U0bmbfnmRbd/YVwsB6sTLF7aWFaNvlm6FwrrUa1q5OMRusYjMci6cFl5BeQ3M7ozI8li7p424B5v
1eEJIbKEr5L2o1ngQ87Hmh+sksa2yDrQeLCQWrH8Vrc2Jq7hwtxlil/niTvlaUkAKqQUoER2weoX
8aj0MSUE7gU7f6eflPEz3F5f8TpFS1Q7Gu7aGctWldhvaJKq3bhDSTRh3+kp1PjGygX85AfHiL8q
fFwdCJyLwUXZEWmMHtr1Hu/KN6GV81BZw/1oXxeY7ZKal6owxU2ygLjiG8+tXNuxoG4ixvs7Kd60
iq7MRTNXlSCq4OK4XJdKhzphaeaT1QKzNijGnukN754ZZ00sqEfqzHFJTudmc+5RhdOfF00arc7v
01ibwId3g162f9pOKy1f833fJ+dWdftTH+d8rPnzk0GNIcfdHm6IrF/n+xzxoQQVeAb0Hc/Sqv9j
dRs50uNHiComvyaUHIPSsAjNaeQM+YnjZQKyHBTcT9Ykt4EItsWf2dsxTjLfPCxB0YDzeXItv0dp
tUcgR9Tsn6uyuF8fEQdGkWDvBfs+ht0hILlQ5RiLfgGPBeKRd7cmyGBeCWm2PdXfDQq3JQpYnZlM
WrgzsY8JmU6+vllNt3aVbSy9OQxx7aAF/8EIxkWWB6YSStMgSU4PTqa/r8r+wC4D06vrznPoBWfQ
wsY424cz0fesa+Eg+J0f0/BFnU1U6XU7C0aG3/LvPl5JyQR7LZ3JgWzrMi47s0xNBdo4iia/tCQA
epFABqTHm07FSpMcRRKg6WMn5Ri7+vI8WurPuPz3EhSW4S+knKdg/cayNr9mfnkd2Zygdbqt5NMw
BAg4GVFLKZNRVfSnXPtRJ+FuIb9uutxvcA38NC04Dh1MbkfscYMXOoc1qFi/c+7Q9cwhMumk/Wnn
Ps0hICDsFWONmZzNIZ9wZVNfGuY7TikURBtz3dmEgiSfzObbw8uhBpr+AvkvaqjeKxSmxjDrcXnW
LqjnT/fPQ+6xCYbtXEgZHCUumQGS+VOq6L5QaKv8V2PDX89/o7RxdvdvDMfRCigZwgtyyFw6As34
1t9E5bvYBvJHvmXSLFwLpc5jIwMopTq+3yvwlaU+1blOVpzQmrQ1Gw+bipaNlliG3oEt34uVfEJy
M1TvWo/FNRkF7cR4GbgIwE98vkfORWaK629PhCcsB09gCbF6UYP7hHaJyl7E9XL/BX6FwPrzZLK9
1LkUhu8L/+s+dHnFf3TTkltILY5CpltUWrwZbL9dMr0u9Tf9i1wB7URdr5H7L9BRBtnxyOQWKZ77
KXv3fCOns1940zXNGfgnnvOU2UR/2kly6THpF1OuGcuY6BkLNnOKBgsFhRZqmHp5u/4/I1NzYg8D
lfEInpRK092yAC/VLnE4fz+9MjTwG3pUfco+oZuy+P0Iwb/OwExcsg0ONgc3pBXtqYXNjJHD8VfE
BItr3gd7PJ8fiYYAeUHqg0uIamtspR+X9bBd/E2zxjjcnnW0RkFQagiNJ+KV8brANCemDKumBbo5
cI6UQRkJYAy3PFM+x4ETzYhR7FXXLTAhNh4a0Hw69WpwYbcScGhXkHwFxp75V4Dp4bv1UukhAjhV
/oWKbsqqAlVDhgoETUQP1tF2OOOxCyJCmyYWkwxFpdc0cRp2IjT3x/TxvFlKwfumyadpM/FLxaBm
G1U9mgqD9GVNRoGsEOyxaSeLrX4jifMMMM+pfYzf8mlDztc+Jrtki8Zgc8YLiL2ITJQkYGuzUj5J
DanAtv1DrSdHBDHOQKAz6WLb56NqeFqPwkk/dyuvG/W2Dv0CTfxVinMSWCmntKGz5YjiqCVP+SiC
s/lLWetBC0PIr1iBJIynSD+AiRWSK51iqtB0mTHySYhEvRx9qimHjbo0495oJpzbthUceHJZUpeo
UxYEyWZa/dZSYYW9wzQYK/cnsGnk9xYnrRVuECkLpvqE6yH2f0ZbSYkIGXO3c0CTd3Ej5DDyFIpX
jQ/V9YWNMyVswiJA0HlaQXXPQM4bBoj/npXau/l9/9vnGL/KtWOiRNpiK2PIv84tgGlnTcoYhs2w
ONs08QVrEOXxPPhd/b0u+hiDJr1Id7mdjpj1+6J5ws8uUMSjybJzcygK61Qmr0LuhNuNkwGv8u79
1syr/xmEimKmAZULeja4tNXxXVHHrfQ2bzKybngH6ZC95Zm6t4rRpq8vUdEWZ2lxYcsrusHOizPE
2Elh8v22b6DGrKD3MyT/vd1lBTpwDo5zm+MAmdyUVRTSaEC2N6jHe4gW9cYEX/w4rNHW11HLJ7Xt
+vKBXmYG5azYRPFEn3cPx1Fz9+I3bP5pQvxZ9ZMGcA4KC+VjibeIV20cRAVGC0raNuHfTlfIyX76
BGwFUmHzQhoRcsWeQMjTmhwEFL+hak4bFKxN9Zm45ii3BMsUr/lzNNrLqqARyNlFZpMr38I78KX6
L8MhHjvveoh4LB+KEr0ghdAH0vlbTmHJ/cN3j1WI5VkYW1kDd8wjI7Xz9DskwDQrslj7qWbJ7rBY
06iCesJYSB5ENJ4kPw+2v99Z1oVWpYCrBWIpY5QbpVzed2REIxSjmRe7Sbanb5/4iDgubhFLbmw+
ylb+Z81ssDjDny+Q/kmfYduNA546Ityf3cAykwoy05GiTcTp09tw6X3GYyLphpFbp0Ik1JWKnCHP
xJo2yVte2iZnHxyJ1CYpfwz67WLJ9MmQGRobDtT7277QyM0f72yQ4bv67X3cPPSBhNBK/jcPkmdf
QE+us7MF8E3JYbtTE7YpZblttHoDPrIyNKV2i7NmvRGccmslrKUNghqw4xeb1MkgoAgRbGpcR8bC
wvNMKDmB1cShDwgSVQG0gXTCj9He8bRL5wb9B3TECrD1jaWQvIsBU4j/6Ad0YCGNswQ0HdDkuAQZ
yzfWDO+F1uQb1eFuujrmyjPOu/7vbg/K/2byoWW5Yt3gGOv9zftx0sFoDaIPcWY097b8rT2FeSUP
duwiEQHe0XhRsmXYh6got7vfxXTg0zcNojdQA7BC+4ZPkgwclZ4+WGz/CJ6qHoQCr8JvJ6U0HJJ/
0i/nRGwWc3Wlwi/uGOwPzcOgZUO4Fb5echxvyooJ2gtMj05pyv/fDfDsHaS9LPOOr8MdztN+Ct+P
oArST50DnlFSICWbMvUpJ7ksRp+1nZ3ul7XwvvdBQ1AAZqPnr4PyOIp6eog+YREPHv3/OFo3XiLn
v/a/UyDiXOkiXEG671s2b59VFoU0forToQwrwU0XThPw0+WS5hRggN3Z9PdKDDJ4ESLA5nc1Uz2x
iktlr2WwDH44B1Y/AVLC+s6dLovc5Qminpf4/23bkNaHZf6tTtxVIttL/b/VNj2HxcoukP1QSlwA
6lYwnHHdoa0C6Udl7ioMT9Hd1lligWQMYvy+wjs6mgA7Cr1oUQ5sKsFA9zxNNoGbfj33yXK6btXQ
CXJ0ln8obpEdQ5UKIEsRCym1ub24hhRBCUraFlsTaQudoVgrWBAvzFgEFf/rI7bWEmDZpa1wN/0+
VQxw4vNuyXi9WlX9W5ffWAbaIGSTgyenCgXjhiBgyOOtKDrq3+xenRyA+xTwN4Avi/YcdQ0NXKRD
CZkuVX1EVZ5/s46owQp2jZm3WUXEyhZljStzxPVWb3qPgmFpEuI+GbUf37W0cr+jWJSIUgY6/gkI
6YUKldZ86KM50mKR1S+FOpzh+52so048FnLHkbUe3BgcZmuWl63Ip/YM0sa/TivZ6KmxZXfOdbUc
u91oIJSWcZOhtQduT8xFeqkXqV7/o2giUSm7tJxs77o+zbQwaZF/J70nHW9CVBeU6nPAKmwLjSTQ
7wAuefVjn00VOldthuyLxU933B2dMoN1RR2sUxjffSirRmS8SpEaiUE+dDQn39U2BkqKSAXNjSnI
W0Ihcl4kBFm1uGPk3/PqJJdSD4U7Q/g0JIIft4b+dYXaqnay4RJB88sMy8PiXBrelApn0/zBuAC8
EPM8Wlrx/l0CDIXZZ3jZyEyzJhVptOzh94tO4fvqaxQ0kaPItw8x5jGGd2PDTKXCI5hTY58WYK2m
3NfsIpkVQFL92eLZnMQDEa48+FFZddX8uhw0M3DO6UE7qFwu5YfUdXH3cDn0p3+lvRk41wycjbje
Zy+05QarFkN0epSrahRCbH9b++oECXhnmwdfNgDXCHk6qvj7EguBtXd0k1+FHDdZkAHksmZ/WKEL
duJvkuJKJGcIayBfA9PT1P8FbHv2g2Kubx/hsWvmNlreVqzu16RMpPMicczfXNfHx1EaM4HuPm9U
zMftv4ep0mdCgZEvpapR3xIN4zU54LSSjCl/3CxNiZbivpDZwPsLWvnbu8vXzi2d0feaSAUrzIeI
nfYWZhTTwLbhRtJbMuolMCOAbiRrTud97Oha9nXGP6gIF+dH1WRusuu74mpA2J5Q8ffRxtO7Ceya
8KXQgReQldhdrx2LyDkfmMhfM0VUaH9b64GyF32X1WZcwN8sbJksMDK8Q/3UiuRBYayp74wgV9aX
L2vCbNC17vMppET00f1/BgbeKsyl5ee1sK6on6MdSfwxbpa23HHfNEj2isqmUiFBzUPEc6qWdSXU
cByoYFb3sT8RLps1wjAGkWGiXwL44axzzQ98rBVCzc3ajpoKlGLABOCMP6mXvOeKw4fAVVNB6tgg
uB/0UCg1fNvsXcVLVD0mBZg1zGXrVMoxmd0KLFd1Yaqm9K4fdv85nlqDgARzA+qWIkq5BbMm3raE
CTGDHKWShXKE/vGECAXizm6ULMKtVMZOO8q0aLFdLcD7iIbEtBP9G7dNZEIjBRUhzEMwaeLJWm2q
0/coFepxwEgtE0hYyZ7IgF+PIHXJwsoHiYrzpDTpFRIe99pzVdRWRoxxUuFhbTwUM4nQE5BW+xFG
SUTdRjCiYFcgspI8VqyW1sRbQe21Y7mVO6L8CZ9OcNCGwuA1fy2l7Hvgik4KgR4+y+8ilRJzoFHJ
NZLGV7Fx1O0GIBQZVvtk+LeExIpKgdY42ZTXARiZh6XBwGXenIRyRBqBYXY4bh0+sBFoSvmvqO6T
0JiL7BDozZYav6MEJSA5wRi0E9xLe5Hw5g3c3ne/fmh2qQdKT0+xMNtds+YTLRQ1Nj2qqvDh3SHq
RWBhpRwKvRXaigadKUjMDKK0nEQoEvQnS4Q4tG1DQqnISWgXZfThwPYPW6g1kYU1XnoVNSv3DLiT
uxCwykHZjSLeslx0zKLn+qVwfZM+GhOboJTJdWA3XyD8sggjiRbbdACeqa9k9ccBlZjRwnGN39Ik
7aWeWWgCof7zl65byIvmhar0SU1fvmc2/RoNtpr9D4ws5OaIPtExfhZtpqbq0iU0O9LLQkrhQ887
YlXWpWc329xXlv5bo7dInIn3ZJET8MQFfmrbW/yt7q3vym+WT2lBUoenKbGu/by8YJxrltgpvjwC
69vEJR2xB79/haGR9XcCkE0/WAH+gzQ6HP8NVc/rHYZ67Y0QNy/2PAAaga111ZCQ3qpum6Eq0h2X
6zt/BYA+Ntftq1ML9sNzTodllnbO2rlyWFLXsG8IZiy9UiJtfRVkJASYRlrwzA7QehDMlqti8s1e
McNB9CS/X3pmMnLxauf5UNYk0kTyBgHIIKQznN7aqmQzKzF90MiFryLc7/8CxgEWJIVSpNBWJgvd
WxhakBhkULFvcjlALly01FNP45GmscD43fTKBcvxzGREnA+o5fl0idni9fC0uO2sMFTK6AyBqDJ9
DR/w+43HzUlyYTZRAN2PdT8YXNsugHOfcv4t87EfYDEgBaImmSdhXUck5ZkX1n7CU5wI4c+6tI4s
g1HunsOes+0XUSZU2n0kuSKy2xG+dsGjntLAkayoEXikhav8XfMScTBOPjPMHHnRQmp3vP2Y4xwM
ky6GHgWCABFlpO818NaWuuQQ/eXJr9Ob+XCZDkxMeOkPK5ho8C6DlVoA6+XADr7tPjG83nYaBF8j
l2lDIluB3Hll4CqtJ97PURbdhY/xWK2HNRXElYqs6Nk0ADm56BNfbVeXT2jXiX3bwW4r/QRs4Cg/
qXxAi8TP4zu/2xQqHunZOI8/7X+weua9q7rrUlX5vXdq+TH08BfM2FnNWEW9NQD820FohuiaqqQF
tLhOeC9TsnfaRTObmIPSXm0RoGe2598dPLMFAU2V7RxvHUBbtdquk9ZBeevurEcUtF4fDoAtkjYK
UL8owh6E7oWj7kaKXjAlcxIA3PdK4pXmT/X8lLPMNYafad8sMjp/otrxP6eI4qbrtaX0jao0AcLN
gUykE9B7X8tUGpcyKy+Yeb46bEh6nIlIIVZOtBWjX8n9pZwhEKizFaD13hRUoVm5C41CJo3YJmwp
zeCR2znQVngIY4aykqtSoTQGaAGO1ViDDjvEvtgY9iw89LxZnCRImYFL2ZEcgu/fHoZHxxz9wCfO
jd7Ef/oVYJSFTrhHcEiii55N1xLKCX1wNx6qG5GlW+pses5AA/trbfnrrpvnq6LKK0djedWGQM74
AabIQdZ4OTlXkLtRp427zZ+yZa/Opcmx89verK8/2fPzn9lgL8fhRq1B+PcDGqzXR36W6L10J2g/
77rTV0sIkBP1yBPjP7vljsxPDsSLmJ0JQx0gBiQVzfuI03VlHva3VrdfFL4eN2V7HhbJThMXkiid
vStJQhgVA5nFQNrs66TUs6b1hBM7cbq3D9LT3I+bUWb4cdazigG/57CLkVeW0+V1nh7juEMVepUf
MZ00XNiPFxyXJ9EcDuiePOy2j1SLantVJzxpF0JfbVB/Tg8av9ApqKV2dD4OVs7Hxd/wsgHFJcwH
w/Gcv/xAT4EjxIOi5zuYr602elN0xolmfWdmIPAK6yn7HRzFCsShr479Jlo0zqlyj0NxgFGwyHLX
HFWrsZxFdYPn33e5r9uiWu5pKPffZYiMpmpaEI4ZzaDTBZA+y/1YrvlXNN8vJWVA6iKehLm2+wmf
bUgOnBXffjL+w1IsVsR+D6OmzI0a2qwgQKJzAd5x7EAeZJx5YTdJWjeTHrttjaLgsXJCOVm94+2r
jzU0g8oce2DbXTxYKuihNyZSGQEfl1vBbTOPz4i5VEWHk9pyhMnEOgKvsQNuFx8IaqTK1gHKmxUv
NAcX2rd/rjeNjmI+o0yt7tohIns8BFdjS//rjel/EXC0O2NtQGbRjfkjCIy7JoKYyzl/YN9NQJ78
4CzwJdvBaS9A8lT5MeNiGiF5l6K0UlAmOzfMQck87i0voisctfId2iJVazrfd/bZ+Y+8uLG6LNuT
0G0EOJsu+5wF9fSzIpJYi/1VJKiCbsIP9H0NyJrSVnRrbEik7bNWCRcJ6tv5hcHnBmZoAYlU5ZWv
uWOFFPERPnGeYymLq4z4pK5T/T36npr5HlllxK6oCeLIpRbezR3TdhMavHlMWbK8rSBvfqFFuoN+
QFMTT5k3dAWmwOCiIG6O12LcR5RoBZKuv4xuVeqr0vlSkllpxwpQBM2HxITgfCBR5KaMr5i7TMhg
hAYIMRMkCAS5xXsYedI1CNOo6MtPs/XFM/5DJcUYZ198y3/J5wgR6zBlrM0xvHF2VgohHM4h/340
uwnRz/pEpJ/G5d+tHyrDgpCqSVxStKVnhC2+NdScW09a63LTCnL4dB+aakHi9Hj2iV8aKJlHzcxc
prnNxLR96nBLj/iySMr62YfmH5c8Fg0uKKs+V/SouHQwlBPWZC1wlPsHYoUYWNPzPY7mNYImLoO4
qRPqeKCTDMEsqElPAjY1FgjAISM9ymblOzpMa0hk0109oUqhsRapx2t26iHCtgLzRK28EwuaCU+d
SR8EbK94YbEluWg3DU+2dmubSF4TdOC1FK170HjNcXZnys0kGycKyZoJiVGV97bFtWqChPML5wMM
PZOtxO0IXUA7KXBjB7EFCTsz/i5cFg4neaGtNLxt2Knsu98UlOteIqzzcPozJD4njid1kM86DWT0
TRkqgIZviMyb96ygLukF4dIHA9OK0t0lZs6Dy6oKiXhnFARga9aghgsJMTD9BCIK0JHJZnI/1GrB
uZrfYJcWl/XCyTv7hfy0Doftj+WSW2+vkcZiDXEPLl6Rzu0vpvfSfpu0nPq4fvcMQwQUsuHd8l7w
TkCZfGStCbeL3wfjrRMWrqBsOhN958AqZ6sGdq/M9Kkm8CwR2+3RFhygB0Amx8iW8vl2jYoWbNZr
eW+lXskvxXDGcT99l4PkvrgQw7UmH7OFmA3KfFUK1VuAxmAfsDO6jVa7A7HoSg9bf+6/I5L/bZt6
BUJRVFAw7xX5xHwIecqbU10mj2hx5GilCX1QldcuiwExQ5nSU6Yo18WHS2MJZhBJwcubN1rCSvL0
jN6tIZQG+BTLxMVV19FU4VfLK/Cr6O+dLEluR3Hsq5r1V5ZXpAzZHK+jxv0cP9jEku21guvZBwrH
XlaMmbOfw/hUnUMCsTpvDmPgf8s/IAaOXdUvz26yzVmpuAHNj+EIXSn6s0LXcdJE6vNcYQ09aYrt
SazDON+Wr57gLClx+9GY1/EAAnk22GdlV1eOCHgS2HZJ3zhB3gloEicHqGnVi8QFy0EttwXB6iMq
VEVEAPObO+osWWkYy5x97P50ZzYUwBL0xv4yVmt1Ik4EONviVkEKt3egmDpsB6LFG+8pPiokAb+U
Esa1IOiCsIv/LpL2AwrBIcnX6d4y4bpifoHF00qvhzX5Lrp78khLaI1TO9C4GY2DLJFHzH8M+JPA
lO0X5I0IKVUdl7wYqiqIondikA7jb+BCh+6YGFrVCQ6mnBJxR1sUCJY0Spo17wUK+A8OYvu0g1JH
oURgdQhZMoyRZvQw1Jorsa0cjgazAJe35DwM5Jw/fVqlkN4dgphys28uYCEGjlhRzOx/xH3uh9wz
wy3ERN+uKbvtfMxful3b6bcCXS3MgzqvL6gnzOW2YfviJVnD1xx6xQv1sG4EEUZp7pWms34ehXbN
6WGErAYei0oW/D1y1e6TNLHr7ePcAOBXAUV6xQWaS2IKsCje8PVNdf8X6/+iDE9sXB9VIKGcE2U2
sEM8Oqq3wl+G61ewO7+TFvz0/vr0B6/QmTQEZbh4RUJveKBAxHkBtE+EMH1BsGRKCByxCHYPZ/hw
V3F0VNrYTOMqte2XLjCTc3tsnjfDtqyf+ri4lYgcz3yhAoiElf8k27cRVGCVd6Cz+ae+kRO5crLj
Lj/mMh+0sLOoVHPlD3D6MeaUQGnf7guuU8iO9GY98eOw2ij4h4+YJ4a/hB3v4A5VNyO7vb1KqRAG
3h2e6VxXVyTVLTbpZ6ZewOzw83Bf8L4OiXjco+YOm6OG3ewboZxZwSrFz9gl5/w/jac9ONts7wiB
c0zx6rIkAgRjffPzJp1DcnIqba8+n5XdFRQJqO6tPtzL/dQn0tk6mte1x/qWnPjpzqlcTijN8SC6
5DN2Hq2i5c7iWu1J0S9yy1RwOexB6VcvyG3yIw6GtepHQydIGKYH0rq3zbXRr5ymMFtGW4g5siX2
QYQmS+BNXKuhe/tBIAHH2oT/giVGiDBc1OcHSFFCTAm535IFPmIm5DhVXAObTpfGIcTyToBCZBe7
VfcNZtDuUVL83ekV09hak/VWhNT4fMwDZV2yDm6fz6UaXKG7FZ+PO2RI5YHHCf8f8MX5fDoM3xjw
CsGXzmO4pTq+od2j4dzrpePQpj/5+V9L9ibiQ3+t/F6BLb+B3gz+OG4VHr+9IVe1wKRikeifD+rB
WDaDGkXyXrPf2ABR9wg0ChAh5RjInJD3XqYy4My3E6us981j+yb1kG5mUeodHYAz1DtC2ahlyjKc
IBGaqYV5KrMmcRdrNVplim+DQXGyPDdZO2sOm/SfwGzGsl3Un3SZcFTGWrdakA4cMIwqag8wLanv
c5Rsd7GknG8getDlBz6wrP0Wz+ZjotBZ+sDKK37ZsKpv7ZwSkLPIcZdGXPZLDsuwM5PN6oo5PKpc
3IhJIVxroz4yjOfgmhrGlPZVWB7VLSjBckCXeZ4n6YvTzpHKm9cXyC34pub3cZQTre2nl9J0boNq
052BcfURY6VYREpLaGAf9hO/2VbdRU+ffy5WuVYHFee2Nko+lquKLLgfZNZvzvuLzSYIoYT+7ql/
Worgn9DI0V7HmeiOVKCIABxzBjmJ8E/28mNeU4COqfJsrJL9b/MnoSr5Hm/LuCFteOf56eqQKYsV
NvXNYDgHe2w/HqTWXUupCsR999p1Us+SYciLgv1XYe5SZQcXE8f0KHOpAXQvP6qGj38QeeyYlFKA
QTj8lJDtLlJCMQflGcpzvoz2XZhvs0gtio1hyR+ZZIILeIBl7VRIrM3lob2Uno3AJTmAt0IjwtMP
P/Zv/mJewywrYHcDHstWd8hqsMM8fztmH3Qx5UPLIXXym+krNxWJlzicWqOSOIqBPdeOlHf7wk46
MvO18RMm4ma8yrUzfbAq0/jyok4HneBgorZs6XxUhHX7vfN0acPEgXl8xUsOPsjbKMc8y+emHQ/H
XzY1o+/kJ+DCKSqT2QzWRQgQCvAFfbAAgTzsivXxGLoN+EDHnWMmAiaJv3trtQ2wt5NfCIGgIAqc
GuSIwlQbzMuO7fc2XYP8opS6Lx4tLNd4q2AsQzvPOmhrDlQmumqO5jE2Qg/8UPqEirDIUdl9lnrj
+3o3AmlGdnkxfVxaukk9JZK5d5KmMcGlsWltmpx6+KqmvpyELWPYNzdADvCck3XAQUiV4M9IWI9W
bN82i0UwmAyWztSwFufyx/WNCuDe2XnRYQO5eziqqzkIwahRdCGM5mdTz12u2i508yjou5xyxfPx
jdUxVld3cHcG5BtddvwZm+VkEg6jVjgsNxjhUCrrUSBb+L6DHOJP8/P8huFZwGe1128vkn6u2X5d
agY1M415wRGq7D6uxHqfa31eYzbwL711clFWqaBO6xM0s/bVrZLNunnhC5GMHF6cgpf4v/W3C6Rt
ZEo4/1oOtFMJlcIJX1x5w4Xi8RAdHfrNyN5Z5/SUsvz522d+mmcbytMLY7WmFjFyyw0Lj8GppqUn
sA/uBjneh2eg/oGscWU8p49/44cz6oYGu6R5+3KEAXZHxb3h1nsn8WFT8w0ZVi2ZKoipPb4HBeqC
s3yp2Eej6bdo7SXul2GXDuVs6kng5olol3QjJISgOq+GsY5sNlo96caD1vY16J2VqqaZsfR5lDdX
T8x8RaJP6t9je2vXXr2DpssBYMV4DvMDjAPhtw9rXjW/ahNFFSIQR07QVqs3NQqmhJ4IERSSXM1T
sFA8Yst5jQCq9B3y7EbybMIp0ooRI0J4lT3vnPA9Ai0JTifSEMpELHKtQz/gmIrPMz6CpN1U0/D8
nvgyvdC36i3H6gadh9xro5mf/vqbNNM3XNUcMf7RuxUmWrxsQO8E956uJXtOKc9ALqaMjYtpw1xU
fgWW3/JXxd7ptekB7ZSg9yTkiTwNMZG26Z888uPvPlaqxt4IHmTOV5V3VE3YP+CS6WzMMnU6arvS
zR/F4LJieSVFlZl6aKHCnqGoOzMsBF4F3eIHMsQx7lCkZK1D6kvJZPaDY+pysbt3nnzWThQmSkMh
LWPmxFX3bmw6ikaXTcabWZHHvA0aFfBPwsDthTcTHODjZm3HaOv4e/7O6lQeRAzYRoej5uGEiM/3
aDZae2YBAzY2DnL2kFHhZ9aNEiUUNIt7hE84mmuHO1FsViok4GJzfkHo2VVM6kp9VwVLyvYGAAsy
YgUUiWWhCvhash2/UkSMUYkmq1Z3LExxI7t5zJ/ktC9WFBal422lpnBHis2APat9jNGLrKPz9sJ9
pASbMGnv1iVC3UcRTEylKRqTMw5GP/N9ksbDHGsFJfFJKjtoGVPd4yCPg6++2dvSQXaLMkj684RQ
xML2/GQDIKt/WpbHZtPnKR197SCbyFpmNa6kET1igJkPV0MKCcR5S/fZ0hXe8RKOQBmpf8tDguOY
OC8HqjKJEcieWPnzhi98iXaCIDVM/X3/eIZIWVH1JYQznjgrcdwkAEFWA7OlqXA+bC080XSsOjzZ
YLXFyCnOaUxSIWxYwd8/Asi8rS/ESoTq2UQeX1inQrvZCIaPeWxrsNK3oOe810TISpEx2orhYBxM
H25rP3QlcUJbW/sVALQfReHKEjJR7i/0enCZ0PJ6I/NOFBTmIH4jAq/EkospNN9t9h6uZ54Vu/6L
zREc35X6HJFy7ci5f5Goncvy0eCMMo6kKhdqs+BuL8iQUXm4Yj2xBfNYQDu6NlIEYDm1icAUJ8GY
uujDFmR4wxG+fa7cpI3/YFZ6st3ZPvqDr1TmroZ8oV9u91huxSnOW683yrReKYt+rOiVReAkVMrK
Geph5NB2yH7Cd6QWhSPFnUD6ZEKqy+Pm3gL+fHuK74kLmrLNp4bY2ZDXWMhj2xtowentv/nW8CpE
e0+1YuvIcUxsL5X07UKanf+/UbUmOUbKrHLkc0+oLNsbKKS45G3G+jO8u/cYrpRvelSehnMyBXn7
O7kOkYetOReoiGCq1jTlfnuL01BIPbJHjbAqrh4EAeKQvPMe17bU2Sekw5ZtuZsQ1OszLGfh9aUo
QsHUUt1urE2sMNrXayrKctdd7NWsWZ5W85JkQMr2rHmgkJyZB23vXcIO2CDVChCxEqID890vTYSv
yZdsqiYnII1R9/9miaFy4eFw/BcM1VdPCvFf9eKwQL5qqeu3O0Q+diE9RyUWDiRQGNd1YLMM0p51
AwVt5r6buImcp+I461kWd79PoMaB+Dti1rfq7HV2vwmyrz1CLcfDSFfH9NO/WPqr1aP3VCFHP06S
mQp/AaqpBNq5qrwJgWGRNr8rZ/GnYcfXdZed6kMXPCORF2IosNDTqWcWWimQ+BCTXJegH1LpbMdV
Jjzdm1hAI5BSkB5JRYxvWFkjeCBT18Td/vz7OOrutI9zNgVxjyyIfo4lbhiLsEItVOJ5vGrGqS2m
yDKAFg7akiAIbo2v/5s7dUfo9BQt4bsM+WF8PBO2vKb7X2Mgn41xoOZ7ujEXnASl9SNZs1USnD4I
onrzalMJb8f29mxEdBXGtBIs4CU2UTOhEpU0bKw6GHiWYErRANnDo7M91vXxrv90L9ziLNMTC5tg
2jr+HDejNgIHyZtUogmmkbq9/W6ZR+8RCCXo9Wf8+LE18kmkPz/EYZTks7jwiJzNXKWSGXv3tSzL
v3Ch6UPf/ija/c2A/vFMvWmTwLsrNSQOG2MYGG15o72Uvw2foTA06x4G16hh9N+cPQLAgOiihRQj
xNymFCMKY07jphvpBVpMBm/xfe4cJDdeBe05QQ7QGATaCToO1RqxxdpaveLcvXrDO/3wj4aN0ExK
dAHLMkI/TGl4JiAMSGReGWOLzwjRfvB5BLr2Y9Yny+WpBaVEnshZXIoWT3DwQyfbPD4aI17Ne5ak
+OUwYgI2xFDswmoUFhMZV/jv4eZlsmCKDQy63vvBi0rFWoVENL6ZKMEIHnPcFed43/waGyQwra6o
11NRdQnAc1+pjV+nFfcVDCXwJ79epbZRnYjL3slf5UBwuoAJGlzwySEtG7abDLdQdEbkjyP2ZfST
C42V+ZWAJyyARhTLd6adWTvI3MBfSJXT0GFxEydtXZUkraowRAsCZucIpWCxs+PN9yRt5enDz43N
TFypzkg/ZV2V5oDb7NsCK2JEaoalrIWpBpNY+JcnmWbPNjYngWy9/kO8qFBk6LKx0LjhTN6vTqk6
LYC1HeEmslclgtaB8SvWLyRk2SMvLNilwDC02OeaBgmjk2n9E9+MCTSvOWUWmHe2He5duchd00lC
713VNJWBfCCTxbUDpo9+Jy0rQKNwy2ZDLOp2JUgo8VqncXW8iQIqqE7nJRE6nHn5PB80ngXFlv6L
YdKPmu3RnrURaWe5aMcWyQPkKlIl7eORrPmOjvHQ6Cize1yRLJOUj5I9RZ2giJ0p8pkHMUpx7Hdz
VnbyH9NXTfG/i3OJe1fHETv/4T3imQQhqTAxra/mzqZQ7elcZH8J3WzPrV/0LHqtTILh9HfW6V5o
iF5qVAFQJM5hIA9VBz2YtWQkA6R+Vqa+kwgOWJcUn15u/XtGNt5cwPY1chFGq2I/0MuiPpawjQ2I
DFxpAsTJHz2DtjuLutdNmwjdD94tPa0+M+2zakjCXgIRpbXDlC7U7QLTcuKyqSjfpsaZdI2DNhah
6bHl8/WEyVffnIGfyDgr4jODyW/NscpUxcvEkYDtF5OvzQ4OglpmXmCPM55tXV4KUi2DVYmvyvRQ
UZ16pdyZDAftxabixJLRXi+lpwEzAKYUYes366XauwJ+3GkfJFW+fNsdZZIaxE25P42iNLITbVUy
SOit+9dm7895PNVhB75vJFDzOyspgXW52RIs9tASZwxMQ0wLk6kaX5eWkv+e1VZ29ujy2DWUGEX/
9HhHoTcOT3+DVY+VkpyQNTmt9ZVZL4oaNkm54rQZrOo9CIynIpOciFIGEV8b5yeFJwVG+HZ0VE86
odL1krUK7SZp3BQdDaje5uSaeITJlPJQvrT/lE5hR79wECZ50pMqMysqF+OapLHIWKqgPcgefrhl
BlzresPSy2MBqd+HzzvMxEnyQKQibeLHjC2c/UDx86HEIGejLBlJ6znz4VfoEr9pG/xV+x1uIJtJ
FL9+PibTCfZsJgnr/Qz1Th4eK0y2c7aeLgMYewHpafO3fpsXvHT2EFHEFYLAzERgWJ7rQ0HDfUX2
y0HnayOzCgEdB2aWvs+TovnggMYky61tRex29qZEEKiKT6KUzOS1q2uRgp372F7QUT1aEBTLRrDR
OqKGtmtrY4cd/PgREQqt91h0HvnktRg+xXC/N1+8tPVq9E/ZVqBIUPLCGZ/CuuqtxhhysrvsGGEz
CIGb4DnpmQ3sP0qCFpCY1LezmS0dawIhIVno1w839PFgGD+SIcbIQU/JKvLpTl/v4F+zmj/sEoS5
6jfzmlNVQqH1jeGLXiPWuHgtKsxHPVa1T/4m3h87llIZkRDY9voD+J2M1G7VdbdMX+PH6756UDV3
mV1hxtCdBqgOpMBnNJnU6VWPE7ujV/DrTGp/eQNgNDdKKMhF2kSEAVcPfRhlQSUaRJgNlKxTHDam
HgVAVbQnn9OSyBY6LB5qtge36SpU9O8awPzfm4V5gWhrB82XiMYLuuYbEhlGsNBwi4uFIFwQbBBu
3y9zJAyHuLFADl5y6V3qpeeyeWUFSniO3X+vexXOdOt8phBXldhVtLxcAxSxVDrKGGrqCobzNZYf
vMizLe/AxB+T9C41YbUNkfxPfOwBPNoQy9kZOXB9aa+JrjxAv5HRXcUwkwIy41i3NPJSUkPZYyOs
/IlUm8BaUej1PavWIU/z64Dz+gZPn+S7CS/ZaSteZKBWr4/qn7eItibHodO8K1iVGNwyOtfxxVvh
wpjk5QDQSwJ7seEjUqedfZvhHAZjdVOppogd+ArF2XhWkzrZBoj4ec932WHo0sAvmtZaLPK6dWPp
iA5ugycY8FYbC6uNgoV286VKADRuC8tAVhMeXxOZnTc6FchyO/kbgEvdcKM1zX/7UotJmzy42KDx
L1oy+dqxAK2KgGHVXEfPq6j6zfp9wmOc8Q3HPKyx3+vtyLrg/XxLyTmIXW0xrrsMT9tc8Z1lbJe6
Kvbs+5IhkKXAhR6eEcNqX/P2AefGtEuUYrg6iSZHV/CiGhg5SjIJkXOAyIotZ45hs7TTnWejnhPg
tfCgZju6LQy94TxMJ0i/TFPhrb3oAc3jqgYfh8cnYUZmUMvRYLa9pv8o2uyNNEP7ImVejuej3Ftf
pEBlI4R/31aBi96KfH01Zzs9Bkzo7uC0M/SLgyzSR2FLa4L9FS1Axvs6qg340nPgJuQeTzDT0XQA
9OiPDILFRXW5cD77nd5YN0R00nNgTFYDhOIJ4xPFMsXx7HgUhfN8qKQYJq93ZMmCxb8lJHGYbgE7
JXHXip1EoLOMgXHp92fQwOz9Yu0da2uq0z8yyhCnI6icmxQ/W/f+M5p+lk2QlXVPMKJmAo4c60XZ
hetKPHBg0wCDJBbAxFjUKKkW+RMZkOuhTceheh2uR9/8ZxOyWNKeaDks2jsD5QyF9Gzy5LO06CIe
zOnm5+Bcjs4T7tFdwuu935DBRjvy7T8lGMfGpymcnZd5PRpQ4+MRrt7SP1mAr2Zct1kNhE5sHxBa
Bec1St/Uyg+J6pquyh4Dy0MIIWvE9nRblCGK5uBhvd5nH2REFavsyoZbQaLGPZdW5o+umvX7FTVf
+K7EEd07QRgR2o+BI1MxRifRn1z7K1PpQo2C7LvY0r6ftd0RRfZ9IEEQ9DzejzTH3zkG2VLfS0Rl
9Sxte+5kElBC9m0iSakD87F4mjlaM/7jxp4V3gembXgHXp13Bou1Q+ACa924VXCks5UjYyyIzVqL
YctnSrq40U5voKD5BwEisEQsfqZ/9j6wZrb2n78Unx0ZVUhXumUtoMxjyD+HZJIP93FJLps2Z8t4
ziZ9tIcP5ZnS3yXm+MqPhuxRG1nozSTPitt0hhf548Hbb4pCsaKY8vaK3OcvrUI7peh2SE9rRuZZ
9onJ2UrPxglGukUo3RUs0fY3M28aabHaPy+wiYXpH7YGo1fc/EsgeSZ6+Af6uywgJAhQdrUtnJ11
/Iw3zR9RmzPF74foU+s021wG0WKZIPZfH+78l69aC0qcQni/YkvCz8ciDVMaH1PGRn4M/BLoBC87
xZAc5FjiYB0+G8ySjSv95yU53qUyjS+YEpT9CCxk1SmojAtpOdQGYW7JnjOXUIZ5brK5Usz1svUb
mXSUwDRxpflO77qTjz9SGUCXpIalv+Q5bxqCEWh66TlHOu/N55ghoadnSbfvHSzFLW1Jn/LbINC7
+X68Zw+Lax2LtLA7O2dSOEnz2da07KRRgXD41MFjYnHSIqWJKl0QmvfM5WlVtFr9BgzV4eC3ypJl
+eqDu4WRkduC4tiU5NQn4TAR6FV7q9tyJNtqgsfiJnX2ZTLn2x3luk/Ukx97TGNdWiBlJJ4GJcVJ
ln7qJTPjJvvRgFjk8R0JCJ4x2dLnLEDDcpPoS/hYTERz989uUc9rp21wGjKUSfYqNWffyT6W2uce
4tS1YD/DleD9TqnavOhy0IjVYj1CZrFgqBFqmiTFO6kS82AuC1/fiEBzhSAmECesPeKAaJlnYfZH
kcGuDMXxNZJWzzGZKZNiXXSJMCZeyDfxMs4DOkNW6H5sdnJP3MwCM+D5Pc9eTLlOXtG+p15LU6FI
C4AZjmUvrUlJoEg4FJRb/Gy59UzjXDD+5eoJ1S871wGO8ze0GphWs16n1ST+wvoZvuSYROML5OA+
MGhWGmt2RGzIRiuqzYZASohbAdPB2gkkPbZk1i5XflxeK4fcm4e0zp58ssv9Td/frLnudP5epORl
OccwLnktCK3WvXpRBIl/hc1Nxc6AyyXLamYwsWaZAGvVXRPW41ZanKx3eYpvDzpNuxnFxJubFR7m
DyoMJ7wKF3n5qN1piQ8TTVqrErqe0PXIhhmZGqdz91xmPubXwjbhsMQIWSMzq4IHGyxrjeQxtSMZ
46CLljQay4NKOky6hyUQJ20xrCx/8yJckO+VdlFywK+DJhppOWYnCkSQHFSnKWtEK1mGlivkD9np
7lMXJDuzNlH/JHR0DunUbSffzlR5tjEBo3FTsFH2gZlWwUsdSGLKHoxK8S0XmJTb1GOIouOQq1Jx
A7SwDohQNQAD/bR3Vrj5pvpljT1IDKv/f9PhMoF15hiwv2mK6EKLGVn+nv70ZO684rBdfk8TKEVP
cLip3YV/L1YjQCOebZMoWM6cmYHaPSX7OwNJu1ID+UJYNz4XSGjoFE1TMM8OkiSmcZCWw0CFpFMD
GzbEmyJZx7A4QajvbSDFp4F2P0p9MqEKW8FVDn343KKSt3Bwn93op14e7XwWaMHR5AI/D3VjbQHc
JGqI39ru+h+4CQXKHQNvsf5f5qV+zTltWIoB5a1NxnvlgVmJgzAgnuYbsF955VHIqbacrxEYAWDC
3J5UFfcmGkAZjDdO7FFbT750u/kngpHQw2XHwjvLskX+/oNgIQb9L/rgb62o6Ggqp1/U3mzZOnL4
S99EtuoK2kJi2ddtK1Uzq5aY6Q8ve3SZUa0a2xJN1gFWjVo8mwI5vmK1eTyBAQiiy6Vm0s1wm+Ih
VrMoiulzyL2RKiL4GRLs3vR7GB9eI7ccMYJB1dFEVspxvDbzh5BxlmJkzAVyToVu3+1nRqAovQhq
kTfYHruxsc4QuBtgFygYqJG43q/HK6PgqjaxxSKDe/40WT8sJw/GXOKcsOACvFmX15OCrlLHA5cM
XoGVtLnfBZC2IAbXJtb8pVjWZYPFK7IZ8k7rp/NM8cwZus8Ra+UM77UP46qUD24n77lP5ps33cL2
q12yiGWiDl0I2qHQ5KXGu/cEWLHl6JTz75Cfzq5tmW0Iuoe+qZ6FkV44OYw+Sh/oxwdIwFL/IrW/
TO4GpG9VhMN/alMB23RyU9VqTi3n99yECCGG9DVBosU1HuGWvVu8bM55m4CFrkSa+Rjickqo9rgl
W/C4vkcaj+y9joI2dmrHXkgbnjjxXU9SFKPZXj1HgctrNJ5JXGrJrwMrFnp5EqZnijM3VH8dynIj
kkeQdgpSs6Gz9q/eO9kUMIgpfyaca+TmBNPFsXmy88Xkw+Jor6bSscibX3vk+7V/uz68FNGGx0OD
b9Thi1GOUN5j78Czw/Eb86L8cvoMy8RZ6UgloXLmhAc/lf5H7qQpG663GWrSn2h6nJjV2lOtd0nC
Anb4PE0roUlXlwrRZIVHpIsaCGdO0pOuwjnsXAoRJvRrY+Ali24riRCTea2MLxAj5vvi+6WcHJYh
CRHRqRVHOiegXjn5lU4CyVLFYzjSR5G3apdCXq7W5HfnnMnQvrVk4YQReC3TUjeUhPuIM3kzuyKU
7Wd+b8lAdzqy4J9lxv5ZEjPDS/0gwRHKPAfM0ZPBWt3LpDRBT93PsQuwrFMYYCzzqoWsRPiO6GkA
MYiWFIpgiJPXym4pLYcld58coL0/MeGjGrZFbllqUg8ioGZku15rxW8Evrt/aEprTZxyZSYcQhtK
gFSV468puBBxGgHMFUL0C9tyyYOck4qXiNeH5b5cecgVs/vA9SA0sRb7vocBsJ53jsTcMBaaGZLP
ojaJ+kQWNEY/B73an2wac0rK6C+fG55TTGDKGnoychd6zRj3qofKCQXUiD4A/c0m0MSOZr1tHQ1V
t36xRGEzG5XrNSR3fmOLTrmLT5wNH+ucRe6tsV/2CsE8fyhwfaAyZgYpSo2g7MocotwD/BAs1WjA
9l8NFTE6Bx8Pf/bKazdy8d83lw14QaPk8opAzzZsJ3ZFsj+qY8G3XwfYulHx3fXsmjGz2IG4YoLp
XNDoiQmgAowAsuA3IivLFL1Nt97jStUTnoUmT22ctqumMRzNw37E3LaslThVZGuxs3LRg3nNBsU1
3KdsM4HRWllqV4X5veNh0+NXmEnJwBFF8ECIXnhkztw4HaJy6636jBhlJT7xZD7NZSvl/8xlqHhy
NCXyPg1xM3vv5bRZvXc4D4sSoBix4c0VTEMMwx3iYDrEjpocT27gfGizrH4r5h0mptvhqoaUNcGB
5anMBGRB6cwAvfznE4EYMRv1Jk4xepd0aG56Klwv/dbUBagYL4e86bcyop/Ezi0qOu6XEO4vi4ie
N8sJk+PV9F7WGjSkX/s5Z5O1i2kEP+03klmiPvK06+hm7HVEf2QBaR4+33BOxbcdA1A0I3J3fKsf
6LDRU7CkQ8lx5Ysc9bBQ1QsTf8rVZCtnvYsI80vqKwrPpKDXonnoE/JuFzdXOeMA5T4qfaFP4Ote
Q7alcjVXgqJIsttu2O/m+x/A8aI1QsCcQZG6d6rZVa0YIpUAF7snuCZ0ZKrp/X6jh8Agfc0siwtM
+5LYRSZ4C4/REzNirglK7nwytVa44KXgDk1NPQMlGbqHeyi2O2Lj9Zq9Ezh7sP1hZ5nkkIHsbSSG
z6S9I9kGI1D1AV1j97funL8NG7F00emy/tlRZnbKFZDwuXruf7W/HDsE7P5wyR6WtVb6o0yPKfQl
u9/dEfGL4JrcTmF8ZRAJfXb9hZ/2CRL8r15AEucKWYHKs1kaUOJtgsd+kIhhTANrxnIUidTX8s8t
KXb4NuQqX0JRVEt0mTmT0c3b47gDFZkg+a2gSMFFQdkg4LFUCv7jhh+foyEQ1xr4ZWdwHZ1E0qg8
ly774D0n9sILiMqd1ieEPCWaIv0c3OaEBugHVdevlkWae6sLb8HahZWNPVFhQCAYa1mFJiwI3R3w
2dqyRXJPKl7sqV0Pcs6ur8vCec8OtctCRUHRFYOBtY7JsQcwXZHjWKf0fymA86qNGxsCKSh6Sucq
NkydCLt6YUhiLiVQ7xqmP2ELUr7oGCecD+fhXgQ0BnDmBDCenRv0y2wiUtjM9s2d5xsWoKACLSWY
JN4kwzVOICF3xsdYc7RgUmOyJ3D0YsQjHCxX+6JQ1EuLqSrYmVyJeD0VYlLdDq5RbSZP0q083XAb
JDJjYE1Os+UgHpTAj/cr/jlAKkfBMKO/dK66TdnElQ4+5NdzkwLLPgXVzl3Y3jemvC5A4cQi+U/3
DbEGAIKVnO7mcVYUM3HpfyGlmgwb6CNq6IMMrJ4ccY/tjMQOx+ZNyEQF9QekjPpx8mYiqR0cBCXz
mzwvCsASOCVLqnReORJUqjgYVvQec5DXyP4310a82uEqW0BkafhEszXMRlArFrfmOwem3gr9WW9g
svlBMwEzmlL/MxdGhowQbVg5jdWpsw2IVpy42wfFTgVWNzctngs8xe8Zhy6JdlMCxVMj7P24hH5p
pg7SH61D2Rs9+ATcIEacbMOyql/hNpCJV5sik1Mm9i6sz7q8TC5PpZ5xQI0QUOjAY0OPRQCGZghQ
ORFmKOXqpJLxOv2uytfd74n+uXMZh3bf7WM9vhZd9eucS3Ik16L+3Lvq73OFyaK5DOGufPNwvq5u
bTKewYSCST59bjhQEFMi5acrMLbmkhh86Vq3caw7eUH3+LrUKMWAT+1DC6Qe1lM1vEUTt8S+6QOz
iPrDFYfVpdFzPGJL7xD9cg/MvQPKYKmbPnqEys0NdmoOHUppkf9EDfIyooakN8EjqXzh3CrsdxbJ
DtIjgsMgn4WgCWFh0tWMKP4Ug21iChR7K+eYy2XBFaIR641FjaCcKnV5AbVImHz6dlJmUd7sIaLt
BZoRLO4qzldAbjjfwB1Nq6nEpjD/vs/d2o4vBGKpqpD0auZSAIH4Ml5+lo6OyvGd5DVseO1Frz27
N6QBYyUKX2IHkyZgJXeKkDSSuxcPzitggMMalJW7m2oKxDweUhqKpBJT8VJbM+tvZniVvb9zNrGg
/G5BmtviX39fQP8yvsz0337K4/ZKK7ZJSaCy4ylYT4cXqHixWtd7Tpdq41lKg9+Mf90v2pnkKPlI
ADKnM5UIjDUvgc+IA8pvh76jeQAZ9hNs/nHIQce/YoNM6nxT5/Vn9bBzuqq+22Uhz8Cl1fwIq54p
8peeRhzspftGWZuiwJ1xEXFEiNa2uAUKTygj/ouyV9jozcNMNSZzL7qvhn6OckTKiBpYapauQrud
Y5CZ5h2ChSopvXBgotzrk1/rDwrti09jkH9uaMCIeFo0TPWvuqFWcCoJQhoPBFUk2ZD2tpMPgLv7
qfsTN105Ob2+4dJVRozBqxjjQeX2ySLE0HZ+QOE+f4sa4m3n1mNlVwZXmNhxz6WQoRIALz87Qvkb
/xj1gvkhmNa5CuTOMA9I6nvwdp3EgAfPTq9Bc9GHqR2EfBsvajmBL81QrG7h4F5XoeVLY58GRv/u
3CWB8d/HZoS4bFQRxAxb+cTCeAURXSHecHCo7QZh2xDFjvbYHf8+RJ7Bsk6b8QKMwVK0c0dVYvFa
Rb000aVwxbPk+4MQNiAxZgtptMjvTjuO2UcWvilutHvcpUPSjzo8FM5bhXbfMhZmqeQ0xTj9C+fy
AEVu8IUfUHUUwwHi/H9FczHUJrmrSufWqX95Ve8Mr0TPW6BCLNWY5vZiGInAKe0X7R77VOHSmf8v
tpkmtDhmwetTK2uTjthhANI3hfIrK7YWzflHUJzXcqPVSH8bb5iBgkOdjqy0hkUufcZ41EVCZJUP
72lA+a3pdTg4IheGtywmwulCrrIcBVXVr/tuZjvIcWHxpY/KW7YI7+d+ZtxJitPbzAUosWK8pnqp
8QpFFQQr4oAFAAwjoE8RmTLhTE35uL83SUi4B2doutXm8qgXAouvLnEWpYv9HjJkZ9NbRHsLOZ83
3M9DgcUN/UxwMmzMcZ/5Ag1QaCanhdGoaWQkkjwVVW7Z97gMx+me51YEoiNxrhat34I5Y6Rz/BNV
DQNXmnV0CQEEyZLxDBIDjwXQhVTYF7IIQGnnErcUAOU1tKDNITPVftdrazKGdYIVZT1SIhp0j2eH
/ZMLgvuq8U9uXqZGTrArbzhiQLV9tvXotlG1R1FCUWqIW4wB1uXNYtjfwxZJb3dtHLbWdNsfbW/C
W69RfDDoRs0E95s7xA99A9kekA5lbwtkwuFX4argxP0Ipt/JEczqNzEpeeD3mv7WfvSrtl/YwUzQ
IXPxD49BlXwqEQD1PhAp9qu6xEZmCp6VQ42oKqbkKtsIJo5Ai0Zf8fWhiH9pqhK5qAOUOtg0Cd6z
NmCzjlKm9OmBZ/LrggqOTqRUTa4qH/fJ+RkTskFibcxQQM+Wp4O6RQEtVRYhpPvqbEbXdSn0RaP4
94W3ud1IwWLeHPNVuuw0MCRsi6sKIwv5RHJOaXWrxmyFF1y2hmwkkq9ENTrPkfbSNHXFBc14bntZ
iWliur9UZEXhdpXbGjUdAnQ1Mjc0q8+ZUecqRNrdgrNmkZ0IksOrLEne0hM3fbsZ39widZZI9qam
+gAsoycomsSJMPz3yhQLpbq8K0r3PsnQmo35L9kLMdLMxEP60nSfggkMsnHeSYnsLyOVe1txzm5l
T+xblZ2XG2a/Ujql6dVOI+PD5bY7Pg0vQh4K7hal+62jPHgL7L/kgEBqXiMrp8t3n+gpPG+peeIG
KVTw4/4y8qwJAiK8HKf8Gf8a+LAxxLzfHMOiBd6u9WkGvkDTtOATtIMeJ73M0BEIdq9sRFQww9m2
wJnauVuKK+4gXRiBbrJiDvMlPPa3XiQDyz3JUXR0wAfLqciHVXnTTR2Rk6f0hmsEPO/tnIZ8kNDi
f4i6JLSu/CN3us/BGcfeHT5rvEYpPIvtH5lZLqJSZ7WI1tbxxLjqWMmzbzjIWRfiVSuQsHav1yNZ
lWj4U3OlLwiShRmM8jNC009iXP96LZ8V+3Ih7VcPpC4Wbn1PYRFMk+gt2PN/Tkk53mx3NCNm5EB9
JobqLD/1XcVl4GBKCNwQCzskC2x1C4y5vbQyMOZn0ABXNILYPUhmTZuG7ZsLAN0dTQcX0fzFay/O
J6uiIqqi4Vxtv1MWhufum+mdjLpufi+SlZOrj014MgYDP6TDv9tM4eEMj1TzwVNg7IQqMaC5bRGf
40vfOhoXJiOg/MPjx5C+VvCTdVAaJlcNrrLe+Tdh2kqI1EUoCIJMyfahDswlKhCEGuwnOlK5sFcE
Xn6Y0FPyR5GiKTkFCEiasW1VTm2R2nvj8xcs4oCDCQLdvZ7p9Pzml2090zEcIQwmnX9pe2jNhjsi
IE68ZcdKiJQwR3X5k9v+PLyTrrdKHNaRK7j3IOVRHBPrYMyVxIpHxyXk1JGBzTatk0AAl832RMpH
HZ6z2qNJXXXleJvlMFPaM10DbIqiY+mMBN9nHGi3UHNR0toLHzvIIQE5PKFSxPa7byApvgHj7P9C
Vo6kTm+hBr1toKClwLrWuG+toz+whe6C2BzqhkCCX2LKtAw3eFxyeh/qEhH2f5o613ZrE7UP2kqA
Zap4DqWxtAPU5+hsC+Pe8TG0OrcpV/7zAllXn31Teo44K5+NJ6lCo+zMBaMazTZ2HwwXfD4dopul
IIv1FHIvTvJFQqVFikqk3qYvDV7BXRU8u716GhJJ6sxtKJXpzasDWcxlN/P6mI7hsAK8J2GmODyz
ND4uJaHmyzUVvv2jkuKjpKVjCNimM2U2KQdAGKR9f3tpxCsvXupvqEPuEIP+5CSdV5ItlNyqckQG
Ut2opRDoPTznAO4x959gQ5Pfo3uqvDN1swKkamb/rAzhAlt32CX6yXvxda8rdfBqO+GaCW4fzpXf
RNbxapfCVoUbpfkiyDHIxDjAIq4Ca36Cd5ENV/79xe0PF2vq8LwWJnAWbx05C0iRxL/bgtai2CZS
ybwPpO3Eiqx1FjxZdaPr7t4fMW+d29FOCrZFiiBXIUxMHnP3AlLMVeVgMfNIlbIl7ZYQQjZDfSUA
Z5zpDjenzTusQ20tX9ltufdhDjbK5dxA/LoA/brsMLtWB6lA1SM2Zs584LVQK2MIyLqdgK7JhRIE
s6fbqFZ1EWS1kg1cpbMrDZPT4sbokCFGzvnF5yvopKEfXyBcUWGxOe1dy8Ep6bsTjH/7hqPsxkDp
hP7/POAXn7xzkYA9jDqTFN1pwBWC5iC9SA1mU3m0ACO1FaGbh9WLni46+t5qr6E4lWqqGPiNP2mn
KKR79nvGbcrPZHQkeNJSYy7meZAPdOlt3A80OB2Vo2/fhUC38aGPggVHQJ43/d3vfkeu519MeCMR
ZytwCVxFuZXiEVXzIr0nh2q0GcFjBJXKB63r6lMKcoq7eJdBGUWYJHJEtVFnDq+0gD6KO4NK/umG
mmplRv5muQ6iGKFOqFSPfjdiJUfJn8um4s+FJEM5bckDNnAsOJcP4Z21PfSBoDb0xzvmNER5rah3
5ewfhreqoxR9OsFI4kgUxSrdkcRxDOcx4NpyeG97cGDgJdi4/2t7Fr0XdqwFBN+T7CKkksLcbzqb
ALlYI/1AQ3DXnbyPO66pXYX09X5Fw7jMgNhcBA0QdFZnYAxZWLU3s+QEihA3ycjUlOBp5KlFbtXV
z2+RpxXNyo0Bcbi2cFrBUHf/QRRIcw0FTe43y/vINMIHNUf2juqkv+wQeVyV2YqCk40in0w1YKo0
r/CQKq0RVf4HqWAAI7VtELNoKoE1YdsjfWRvsWNTA479Manax/Xbv8zcPPdFLSQ8Q3GTggwLZXRj
2nhAOPyW7cVGJ7vca/UdjshHEy070Odgbr1Nb/CM4ZVIx2S/GDNpB6eeYjV9TbBRyHvFnRjlXQC9
vHlLP8mx4oa/DYh/lxM/jV5ZgUc4ANslp+fxiNv1BV8gn/BaEpvq/16Yt6jKphCUGIZs+S3Y9QMB
EuxqmKGI1OGDk1kcWldPWFELvoL2uNdzUqH8nyXIhvcgLaPTQ+X+/MfyeBr3o/1IOcQRR3FTaofQ
N75mY4lbiJf6IoOdQNjn+HwlJrrbGYU1xOMUKfINSKwo0u6T+C+Tkb/3aiMZ/xL57Z9kmSnZ0cnr
/fPJtslE2LueGVhHoC31gRuAYywRWoEsh7rArlW6OVDM/RGBzh595aDtX4K9eX0K2YGjtuAM/ghM
Yh5eK/FvCdDKe1auxCNKe1bHFWkH5Pl/Zih5nRXzmkMQbCXD9jIL8TCoX66UOaoRjbwdTW+gHiIs
vk98P7k0GqPXkUy7XIQ1LGcxyweQGXUo49oyZvWorjDiI7uBhAYPBwARdkT3jU+AdKKlMKld07lS
f6Dz1LEW7lo/y1sJlQw8j3T1tU4p1bdCQ4hULC4rDGIrInyz7KqPrnKBVnOxzdWFgsyPFs4z00kE
COdOIVCGg2QZAFJorldVLR9fgW8tstHS9TMbzh3ic5s3F4hFBiYK7+hpfd72o+vP54Nxh5lx6CVC
yKqf4YeKc/HkX0eBZ6ITCzSETXiiY5wiLsMk8jQCxYEPwU8nPuofjVAa+wOcrP6OB57jkpc1Q5zW
+PEQgKbOV3+IWjZxV7rWJjnAqskUyn8am9KjCk4BwcuuJW1u6i8JyRGdIS3JOEXAYvvajvm8rE8N
owkFzRYsnsCwxqGLTaoYVg90eGZp4WKalidzdH/rv7IA4YvyqeBZd+dxSrau14wva1VULO5dREcA
t2zu9q8pUynGv0VpVEUUnL/o1M9GsJsvRxvYfPfZzJE2OCX1J9qQDnMvYzUPzIv2uGrkn9fgkbAN
hy3FZhPNmFVYMDTOk/z21GUt5NajMnmofMiorD/OgMB1zyuw2PCoITkRbFKj/ekgA0X0LLOc3j8M
eEFmKdcOpkVL6nYRXK2yHW5/BQf+8h7Fw+7QidkSA+COT5KpBKElJCTzfSW2oCkivMGejlHCsmqk
ViIllU7qebeyHP8RbgCtigutZH3YJLkf8KNV7+zpwDfb9zn3GUEiRvXktZY31BEnakRSxHOvnl9+
6qMApLpL0OH1Rf+q0/oQ9f3t7awOuYtnbolDhhQWy8wn6tdSBLwI5AdT0n7OkMjpv6Kua2c7NTrF
w5xvjIAcvp3+eGLCkA+xNMNxKgIqif7WebrbBqVyBJqcfKWwiT/1NZzmUgJrdTY0JJa0FtmnqoD8
vU0QPSmUs1PZgRuzU4kjIkiDIu1pFuHQR7OJCCBx4S3BBV7mXBNz3WB5IIVHephWmql9Y1xirfdy
St3PCeGNTeNjQ2vHCi+LAaQaPCugy2lE6/V1eS1l+/Gpd2PFQMlrw66beiabF4aeuZ0v/gfV/SHU
2Y6X3Sf3FOi9UpRlZtW2rEbaeCHeKoTyuuAf0PSj+fmnQSjb9Vln9ztR24RdSdB4B6LhlYZhrzz0
OQiwAIucckp64pJyF///rSXEK5TBOGi0SfSAvRaFDpiBLm+MyQNKBgKWGZXCYE3JL5FHtQRmSd5h
OmGGIUQiHCUSSkeL86nxcsXnQ77M49vJPW/4zCcR/rnSBTJYK3wEjPAKlvnn5zDZg6bafNJqkWkO
FF3pzbf9D2+4MPF2ccODDB6CoKZ+pTq91/OHruU2E/AjF7+Mki5C3dT4jiTN556T3W9mMcJ2mq95
oi3FRGylE5S1y58Vizb9UVcbQ1xl8o8N2Rr8IN0VBJR4N3c8SPmcHCSZjPA6MF2f41tSr9MOy8tz
Tv26ZZcqeQpuL4oabSBTJOuEZMsOIkidWEYk0pbW78Mlw7jcq+5B728VSvdVJJA8Vg2VYkiPc/0i
qeyo6iDttLqw1KXgwnB7AaeNrGR7z5JuQiqRw5NJJqT0AoLIQaGixA7UTTVAcMFppGNKuGmBsOpa
2RgBqbzFI9k6TPxgbQlLIzrSjkRvqkt//oqGRqOFDdc31ZxfXNJSxcPGvjLL43DoNplvC+oCYhUV
FXDgMtv1KRMJlLqnSV5Dt9s8yuu+Zl8dZwpMQYE0xTTAK0FIwPZXyBUKuPrivukPHYz1HmRK2SKl
7VV1+T2cqrWYhY/jaK2gs/vGB/m7ijGcahwz410U4K6t92r6gCrtpOny2Ffxz48T4tCgjKJt7bjD
WZ6UQBNoHokOR/r1HxjrHxExmRWARHavMTstDFUGhhUbOXYlOVp8oKGeIIi9czvXNoO60h/A4HqB
WDT8i2+jJgyxxlWS0FZXj9hRhydym8BfY08EQyJf/I6B2LArRgvJ7222SRG+GvyrHCf5PKRET3q5
fpPSAbA+Y25UXObZzrzslJsY9Q78DbXGb2AddQwipdc/w1k2r0NIi3fbIfLMgWZ7qk/NXCV60MxW
/CgqByp8Dh7HvlNgDCBwNUvk2CAfUFNNigLVxJXDqZSf/JUniY1KgfbBGTvaRjp+IMnsYOmCUXnK
jZAMF/eIjt4AW+kYuBNovuWvGFpPJeqcn0PLdv1NTlm/AnuPGkLa8oULpx/0oMAipAO8afRsBW6y
e029+IgKqkFyMORtWqR9BAGeMVMpqIqpQPvBBhJyFX81b9bGfGM93JmjlA3/XJlRQX0J6gerobG4
k6YBROUQuLx/mcFete1Z6PdaWskQ/yZ2tB3wlf8bTiUmReItLKA0omo5vHaefTNRBbA1jPOnI/rQ
M39+Jor+8TwubdI5GILXysorXNWU62bQHo/lYvQmE844m4g+HOzL4JGINTtmQdTCM93Ggm3A/Jyh
vxNkBiaCHPywPhI6gfVVbV60vzdwXumdBxuhUxz34Ww0sGcIn7fgskKo1PJJbxQnGWYKYrE6rXu4
YVl2EuencsgFWspMwQf6RoPQaZ/BpxzcSwXqCXlVR9D5JNITwRdTzOS0mW5nzmAuU6ox9wojnmId
xrQT+BA+X/vpVCNM3RnDLRz5SbnC4K1lPgVvre4HgOtNMLvUoE7dDBEdrwgVSV5/vlaotFCh0CmU
kdOkppVuZndCNMRM4d2sf4/uibOajV1Q6AikQVjqiUbRX06ILbTzk60mrtIz+VRpX3FVPsutfTkF
L9HfMskTRDjPW32/Dt8RgwaatVtkdHcd/5We0zYoq9Izg2u9Wezj7GVB+/mnnsW/GLl9wG+ziGrx
KgXWfA8wCOe9Yh6iMhMhcj8xOBBL6Tdna4vDWB2UrWNNudhqPNFZpHw4qQ5ppg0MXTJNfyj0q8BB
RXs+rZqM3Yy2pJyyLr/6q5vX5CwpjBO72ewUqOPl1p7A/FXxZQSY0NFhkbf8FlwJAojq+iw3NXQE
QCVdTyQMapwGETsqdE2IiHUCwS2BKMy09CxNfw88Vja8MfOSlbP1rTN9vFHmGgSDpOywIKUj8GzJ
klOHVuriIOnoYCmh6bTGzN9CsvjzC9xDgQGUhOPrqU3dWs/eEIODHIAvTFMkyoehFkjV0vBB2taS
IM/K6Up+wn5DLxnetaTbHM2GIJHA8sd4xZaa2fge/6Xpg4og1RtgpsF/Nd1ucYBbnRv6qZnPpZvp
5k1xi8Uj93xgfJkqly6zmvEzsgmEpt7w30cd4dXffGQMNBut9FbqKlFXLCFkVO5o4jCbdVnecSKA
jqlWMgvVldeUbzYM0ZQk3uCQh6gEGQIo/no9c8wFhd4BDA/aUQKegH6JbPPHlDUFcwOC4bXxZ+LC
SHz5k/kVxBaRyXXc/i3TdCn13flgCkQrQwqwhV1tC1hgBVKs+DtHapMqGvrbfCzKkyfDc0qwwjxj
LOLmGrYIunTBqAIiv2nKS1Tgd4FWV3GwE59ngn1H5Cci29FCOx/yucIi//GC50EgZoxqaIxLKkxw
XCJ1P8J/9tHVEcNfXoJSX9CAiYmk3wsQOyyFfR4uBpWj7eb7iHmr65s3Ud56IrSx4yu1QrK2vKPe
3lDcqoxW8b0C7wYUqCkUDoLnLYna21AhEZzhtiXGBonM4j+6diOj5m6EIwgj6neonkMxk0bGdD3+
dsLpPXZs3Pa0ibKhcySD1G+jazxwQVOxZvSSGktWy2yBlcIoTErQ1gp3/fTLm8dtimtxYob5MQ6u
dx9mdSDDiD8FZDyvDRAsImPpfiSzYnhQUebF/gAepuIQGSumZYUyo8ZFouDH50vjIRL0knnV9Tth
HD/wQGbIlOkKWxIRjANVFoOLTfg093cdLBhyo3ItM5Ql1d8suj+lDwV5hpiEq+mcfTlHBhLGYDWA
n2UcuLv0awirlSkIU0nBj+VnhoDgg9/xjDLvEVlRU0/EQP4y30apRTIiW2KxW3f9/KOV4ybr4IXy
eaonkrKDXl67q3+7W5OWN1f3aSnu0h5EkTY9cR8iJbL5x80gnvYNVVxIsOOY8Bxi7OIw6fiYUkF1
yqCnKIw3+fi/Kj5u3NokECXW3yVzGRfW0rwIftvyKW7X89TAmjtVT8nsYGjGk+jpykRsfQII+w1K
9QI+BVj9QFgEL7DJ2ZGcMpdDcbDHmkOiIPmHm+iEwnGicFqw6bj7XDNNCRtI3wXXTTJIiO+h2AHP
fnwZ0jvKPQFfnkQVGVfldJw4lDygNqAADzKd7kIS1Qgr1gKPu5sSUGfeKGpBfRfJvOW6wVScPj/s
VH/YFLgRYsYYrRmkbR9bAX8yDQjAKZL/HIaBiT4pGm21H2capKHEaRWxA2ACZ8GbgSpkmdRlObkn
22ScHr5tC9S0Z1VFr8T97hAK3R2RMx8TZSfmoQ/j+rYShrb1wcLT5HLw44XXIUmXVYyjWc/TFmmj
DA3zCmBHVA4FlxqEqVJHlR04euKHppJdReLx4aNjyW8E4voJKu0S2cXUfA1Hf7y6h3sbCFcABymc
qzMHMzjU088AuK3sL3HUCgaYvo4P3PqqbXrN9NXPSh2DJ5eP4CB9rMDLzCGxXW2JfcvLHyJq3AUq
+ErCqITya2gzaWen5CZdf2BfUym/NJ0fSXpJq4vrpDGWacYJSoUetzhFNMs6eQGzIwhSDaDMGSvY
Y3iuNMwMPdDGx/ZQnBzOqOy577m9icaLnpyat2FmF+7LqXqJa9XAURoY5luzQzdEKj0yZILP8+yZ
9Z9cLSpqJRckajgjUAVqT+6eASh4e8rGUj21dfHtiLPNnjEO3o6XpWY400Ex4kp5SCY/L1r+O4n3
d55tWU999yuvKNt/GFm7P4AzPTLkycNDShHforJr3p0iVtm2IMlNakPlZWQ2s+F79zGKBDXqX6ge
LYBJgp5aQX5cs1PRc2dLWkBR2EJZAcwLxaolsxmIQZ7g+K+Qli0sdr8gg1dfOiGckVrUEjFHH3aX
e+oCh7Mu6S/x/RaksebqiB3JtH/Es6B/xTKvF2USPh2vQnpJSVrSSX8rC6cKJ61Qg5K3K+Yp1rBC
brzkQBcJLLRL3SthXbNEznLyAZzJvC9Y5H3oTGBu5q3p7gGBWEVWelFw4cnq+gaOOCiV8BiM7ndG
voPhTC2sWkvuN6WjEmgbJk099NsIbJnr34jl0FkDJ3lJzm9gEgC6eokx0qfxJBf6xrhd+PrXHFWK
JGE3pOqeQSCY++t9ExRC0njNb1Vv4bqwJp5KQU4x5Qh/utJDqR4GihJtmGIYmf+N+gBc3NgVREon
TGdLNtDKUoJCy+PE/kArQErxX8qr1nMNog/Ed1YAhsLlkbm7EnplMUngelK9S3i4GDHj7bX9DR1q
22y3aGWfGwpC4Kd2TVcC5WyJJIrCO9vCsTjxW9BKUmUABmbDkCObhGsbUtsgrbiXEYiBc+PBiIpH
852f/kAXXRUiMSh0wm7xEw95/mZFXDrBUzIkMwnelZSJOm4f+p12VHEjtO/xnXfBEv8R3E4U5TTP
38g3lAfQ6t+9g51uypdFl0/ciFpj8D3gAusTwxkt12HIiUWJ9FsJtxyEkaYPOCGzTGTBrueDo1fk
0KfZFccNE5kqXfqSByrsoQxlwhK94tnKfgS/GgM3yK95BXJcvLFt2gm/YwyjOu9fJPmkGsQbZGG9
Ri1fMaAfcuJLatZ9Hq8EzDPfmAZNwsMFkohvr8SRHtFJOIdP8g8tiXABy5eoFIN8qAo/irLXdOLL
M+wiMlTCFoW8yqOpBIiyt38ez+KJlis8Lr6OTRPlZpHxWdufnbuVmPPeCedcY5nSkeQYVjSzX+G8
5KEB0IYyggMXt53EOnbrtPka+yEG0COk3FqlXUjV0v6wAW40DYW59pt15zmgKSGAT1kEkBp3A6Sz
fP6hwdZ1PZ4IcMgk7pOSOEuogIMJJrMZkpxhLD/THZIZYSZioI0sxQZX7F8Mqz21zm61qIqEjaO0
5VNIFfPfKzCNyWyolo1fKvfEXC87hbq61VUetEDLmlxtmsae38NDLykyVexjnNw9Dg66OdcdTpQ7
awNQrsyMTDPNPiLi884HPlRc6w8AZ/LvtScgKA+yMa0PW7vI0GkTN6PECyyAt0qzq0eLTA16Cq6g
hf2XPiniEKxKXAjJnG/UMo4/HuezxjXxed3pZ/o4WI45ljI7uu8g/QJK9BKPb4/D1JUHB2Dfb357
2ZQKkT5cCEEALfuRQ8YEDxtZfjKD8pH9gqR33ehJRdVB4aKz/7ICvIoGQRASHXLSW457/98Qkh13
FZini5uoo6IN2xuO0NZUsLWb2yHtRowGMquWIqTVuod6ElwdHYU9MpSeA/u4qEqBsTolid3aU1WT
rxB/u9gEUCCZAsG4YUdbSHfLa4y+TtKbQApKrIiBwUMOLjptbGBb8ke3w5LN6F73lB9Dl80y+mMQ
pfgJUA3yKRpx3koKg4FUCd1Os+gKAc1y+3o/NDCJv64NnTKGpYZE6p7NB0QatQuoORTuRvxnUTz4
DFUVuZuqMiVA3vQsSyEcvoxAxqKVsIAkmhlzvn/9DRU/6WNrqVx9UhMY6hjegmccFSusNZsHOkwr
+6WQ9hwGV9iMAInuT8Nr7jbgbarVYplYqR2aasNcLxVELhZ2YXD5G6CfoANGs3oc2XbonXJgFt2D
5WJLO5gnjwYHTL85ySk0WhVlQiyhvWG4De/1v2q0hU6fjhuwV++5UHr1Bed4oa1l+cZLcTsFkkKy
iRhlEjZfpXA7enQq0FH0/9NxusWvwg+fJ4W4RKmlC8MPIehvP3XKD6b+bP8HdZx0h2m20r2VQBbY
8wKAxXDKn+cFcqThTO/5nI/S282QRr2Rw6FdQBeg8jFuA9/evDvsEfdMAv7sWNDvPVGHYQ14EaF7
OP7YHdhxZgBqxiCccUQv4RYWDNen0E1BXzbYWoJoilgKlpSa2nnO/kSeS1nPUBKD6nQa91AdVx8q
08lZo7kodWkexX41vr58wPPegD1um0XifRUiGEzZZgeABdTZZ1uHpWjjhTUhOGhx/FbDJoYKM387
mgT1fog3XVHmPEcsU6vunK0M5tImpnoye0qNj67Fu2nuJRV1aJqWys9z3bVUo0PHL4CNZsmSGsrn
jHaZ0jZR9y8Qi5U2pFzu1RDGlBR5ayhP+gvWYhO9Rnz4bfkfQPqnAx6idrvxr+S1fz4ZG5lLhK4z
V8gTI2T3z5DoKYuO7vH0+KijynIcE07C0qchSuIOqG++MLZE9+gfSghiocbQ60wlueVFH6JzHWps
z2bTIKrRVJaOX1+zEAITuXHyVdjzdl62xq3PbWj6aw7Cf+bXzw2X4I3CrlXkBgb833/d2s03wyWz
iZN3TtORZ4WatC88qQ3t2vYMWuuv+atDfUd1scEu8kAawc8FwEKdXvDyJa/wwqritg6pEvbuN1Zf
OMbfcIriX8C8CP5xKh360NCypoABE6WYYkJRcf31LJpR1wg98BbKPQu4NABqBe9YpiOTJKztylBF
4FMoqEGU6ZFQj9iQiw+ciGz932orv4l4vrv0dm+zZc9cIqnDugZ0OC0ZC1L+naieuGhPKlH94Eth
E/ze9p36zmtV5xKF8qEO49Yov03bwTIvWiTcTlJktWgkY6ugW/2GsETE36wV8dShDCUwr4qvvrD6
YT38KBxbW6MyRdZL4poL3SSDFRPI7EcLzQ3BzOfIUI0Z5Yl9eMAIxgxukZBwWO853ibw5F5Kkbyt
7ZqvNVaC9AWNphoZyMwzyVl/LcHkrrgyiasg0t2qwxSxPfAUi2H/Ho8N7HoKF/rlGU46dQ+4jnb/
3sr3Sf3wy0WLrY6L1PWdImM3LhApXTJT70k56O5XIlBl4qKZMPVxtShClJl3zgzgXTOTBhMuc3B8
ZbBh8Pud37dgOe9x9O21WcgFNnRlrHb291m20pzc5et7K0y8U7Z2dGFTm09wdNDxPZJ5iDoacGkg
FgF1RchwQ1cfJmPzovwoS42NFxqs18ucg0oe/EiJmO5CwLPJpxQF5svctGnim3g7LvnOPDguVV3B
oRRShzDYE+shUVyVCUjCaSSVZ4BtChQq3Ek5lKm6eDjvFKk9UOZil76JxWt2MrHPZ0hEoMm4rcFq
AJJPoMbnrF615cVocwv3cv/EY+8RnHFYsk2/Env4TV8tx452yf7aeH5qYVAnDnXY7/fYgoNf3d+C
h7IAWkHARzwtXF9cbQg8VSQ77Ub+XqAZAirB9Dm7pFyeXZATn8jQT4b8CV9Sw6NePvXWBe28nVGZ
6AWhYTwXjyr1zkZdmqG/A4dQ+KJuBl5AYt8ep/pD5IHNMiIP0WsIOuNjcQrQQ+O8PsBJA9BRliaB
/TrmDRCP3hX9tJ8fv+GIa5KHyJL5fA2aKCb5v8EM2lBbFIHFrdrPbu7O5K2bhoAQ1UbJzVUd+zB1
3CFBF28Xl/O5pMRMLTDHH38iflWsyCQsPHv2+fdwrZFyvBkhxPvXxRfodDH37lRThhmiWUYxTmnN
BSXMovD2k8Zd5naZul37tfFTyESJCaMghXKDOqXsCOFl7OchVyfrXyngqneJC0WtO0fc7htcM7ok
O+nH4pviXaCpdT4Kksk4DvvTqmQ1nuTZsffE1oShMsEb8515vXKHRXSc/aMI5PVSxHX5Wf9iu55B
G07mShB+Qimbo4NVKmrLdmB4c1wyKQiWlXZPv8ahXmPa85VBc8Ie9K/mx1xvaG51qBdcwQFVPxUL
eBvgzKJGOgzRGiaQpXWkSvOe10//Oq5f/3wBYR3sfRhC9DGMeG16gi7qthaJHGPlTv24MpglM2a1
dsFRZ5KOFyrpWvC5r8w+cdo8UaSX6r2H5hiER6ujisSYybqQPYRzE7y7iwiKcB94Bwu5npidv5qY
YaZplD5aD64wmswtn3GJSzC/OfwATbYf75YtRUSfJPdSYMExNwlnQrO2/BKzl4cTFgjZZIIgRHMr
gnXBnvfjLE9veCV/GD3nju84wNBS95/QojAYX+Eol3EPv7IG8IjnPdNSQQ3DrX7y1Whpj0Fj43Jr
LDFmM6byZyNxKi8f2xDdyTnv1Sk+yHLgRCoBsuqq/N9q/vKapSAe0z9mTGvVrCEiK1OBFNjjP0Dg
oBjQwOyEuGo4K09N2sLP+UN2XYWwJlAYzsdkLlicHWw/IOWdFmgSbj+uNepUmvDPYvRKxRp/KJmL
0H3UO752WtnuTaNARkbh2024GDyO9vkx2JKsyuAyaaa8sFrz3w0xtJpot5HzEBC5/I8QKcCjNkHF
VfK6s0mricSBVip6IHBsCrpc8PXMyhOolayowTlg6eQn55cYSzEh6aVzxucKUUoSt/bTUozN1wMR
zKOYhdT5tLk1Hx2S5mJaUIIdLzPlJZtXOIboLuoqLGZ+AWjxu3vXbVvbIQ6UWzm1YYz8lGDGzLkv
REwJaUuwE3GdFpGbBARx27NDD+Tju72tM2mZpmYsA129KDsjf5XyZQYm9qinZtLryFZZdp08YeP+
SicQ2u0ioA4qWQRzwJrHIJGh/ghxiVgG7QRKfDHGG/dncTSrCbYHLUBDfCQFpzb00RXE59veQ9f1
iq54nLtha/7+YF126hA8jc+eliwt257vukU5WR9UDvBzBGu4h8eU/crek/2QzXpR0Jakb/FV87+t
DNPF78Yw9uxHXkuSunwiuVtlTbl6HBH0uzQIK3T71HYK/BWdsH0EgivCD4asneK3hSRL9xGbBxp4
0TOgK3rQPmYo2RL0inG3agEn7SIWKQq8dwsGgTizIYgdvYjpmywox1e61wgQY/JdFaSU5glvEEet
MOKr73KqLJ+K4isu/bF5a2ROzcCzYEfj+I2y8URcPaMGAoICL3d7+rjZnQByLJzv8Q6nFRPHRYq1
08ccZctA3lLsV4s+COMqivo3ju2Vn9J6vCRp9+g75kxZ2wtPnfNFEqrgjVXBlXyYWh8TBBLk9z7c
IEK13PCxPfVetoTVgi7on3Djj2lvQhCbl7PaDyTTZ+S9AT0wSpJobyvar3hYiXuVgk43eEC53BHQ
MxpOHJ7OOtoXoM67wdKRvSXHzOsR188YOMyZ3i7jhkjeUksQOjBoO+O89pLO9sdKCkKIb07SbngM
xnedHjPQ+JRQsSd1KOSzeQda1Qu55cK5JflN13JwLugpFLj2ll/R48gD2tdCQcLjsxMAHQ3wPq/4
StGVlMWjKuqioQj+q2yZ8bF0vOtn78paYnj4CClRx2vuHSvkYFvOWF/8gX8K8+3SoMhgM8V4Raze
G69KnWrZe2zKcB5n7cul1oWhXwxDjAcbHD9ulobXDCAS8uPqpTPNN3VlnQDGmGYYslmisnenDIg4
0cCFvlwVxX7pgF5oSjaQ8KxboPtYgbtFr2QNz9vUWHrl4WniVl5E+5SDfGJzi/auZMF/DD77JdCh
Gp3tzsEef5176Y1qIOrosg+CXSBEq6z1U1qomc+RQNh8VVjGPZqkrYhh5s4oHRA0fiwEjxTUK8Gd
Wx2Hwvrr4ZxVbfQk/sA65HLT7wkdziCOZoN9kMOTpPgL0YewngESJsz2SJDBvesOyigjlvcIIGNM
xvQid2/mm4CFquT8bZqoagZmurhdQ1hV9fuiOTrRFaxze17a3gNAU4of91i2CxbaQYcoHWfpeFyw
O+nefJSwqEZhosL3Rfc90iQxIqX5cGaMfZLfa30Iv5IMqjJr1SUjiiIecjfXdm2Vz0Cfwqd0qlSX
C2JWfGF/PdqjvpaMIKfzy72MynQuxD+ensFvBo9PF5ipNgBWKUevy6OQzJ6Vwby7q14qkwHWypm5
cldF3S3BsSWaij1W0xkKvDmN7t6RjWHApD9TDmT2oK4mqdoQ5DU/KXCXndNmX0BfN6xYvpOqlrPT
5gwM21QqO+z3mgbkwVPYAsAnKOdIYDDx2qewHGYJCZ7wGZmZ8LXr+166YuMt9r8wJDd2ejKdLkWp
o9aK632c50Dv06QF67jOuu53SDEhnj5etSYuCEWqzyZoNWraFvY9WY3GsjWOWBDnrc6Tba4I0q5d
pipx/m2YOSAM2C1P7EV7cHbhrcQ9JZF1zsWvg37o3Nj4vUjPhY7W4I/EBXigK/SvCJ0zKIsWnda8
vY+dh0cUK8Ge0CmVbc+Xq7WPM4RUziE7zVfZ/dD/D+hO1hHWB4SubBdDXoQHj+53WUcA4ITcmGfu
ksXMt9cUhM6evqPn6wBSizXoK/8juvullg4a8MUjxokgBRa7QwniMtrintyE5fbYZ62qC+kC0/ex
ils1PWU5k01ncnbHrY1j1Q6SWeqfwBK8FDnuyMPJJvNrVYVum4V6gdEGyAOFVjnc+zLUoM6BkhFS
+d/+kaUgj4CPFdX4U1xibzK1aI1opTJhwosOwseXoSUH0gXGWvXkicbf8ob5Qie/aU6hmjmIyiqv
CKrscupMUwMGQuDMREIlAZEicAzyiZvW28ljIsA3F2zW/IbClg/LLl3U0smWnUe9/LRUX+r8ZHiD
Xo7264VkfKtVlNMBOTttJ2LloLfvjk4eaJdNu2aPMuQwsN9t8D7V1tk6beqev60inkcA/P4xuTa/
ZqxQ+4NGonGcARIsWrHp+92tUqHIslw0yzWBlzvAAdX49uiUwjEvuf30hfxGtYIQVlqbQaiaaI8B
6vKQu+bd0dM0tY7ghDI0B/S7ABbL4+Bnb1TQt7WN8XmIdHYfP1KC27X7wxTJEEx48T2looVuYpS9
JfCxbHY//P8Q+VeBjrza7TbnObo9H+9X3gGfyijHxe2lS1D+ppph6D+g7sXdrV/cXfSW6fAEO014
m1Hmn87DyPR+zahNvsMu2DSc8th2dS+pi7GKwFmy5SUL6XRVDeaeWKVmRBwuS/rK+7Wl/OiZj+Fm
V7mYcPbW6+F5dhW8+8KhrE2UJnHSkSZL4BRbY8/xOOBRZYHswqgU5JWsRPFJLxpC0aKY2wmIK5py
TsK6tiSyly8furB7Pmiv0ICJV+Ct+EEkc42WCEkX//x4x9+g0sBkJsHHrtWqE/xL7N5H56LOi2d/
aW269mKBU4szQFt01rIC5zity9FjaVsHxC7eGwD03yCB6GlfBpt7yzbU/Zftj08rouvnp9cpWovj
yqM8NewWgwr5jAZ1h5N0idNZ0rNVmV5AgBe7BLn8bfPC5DprnVlVPvE0ak8+J/XAn+x9Ciafrqo9
HwoEfblvTrosKyttOSIwVxzfWIlIR9g4SGASnzkx8EM9sde/oTYmmkualy1SatIEsmO08658CAoO
Rn1zcVw3yv/tXutlg/GLnWdYdY9N7f8OQG8YbVnIByTe4AmnJJ9BSdui242VWqCZ2WwrJk7Qvudf
YBX3wMGVxD8Za6geHifeA9M3oQaB7SfzVIsNujlOdBRhrnszZUSLh3BKzS6X0kxmo0+Jn+C0f0Ux
BnaXh2miZGg729Gk2gbGDTLBXlaUURKmralkiXt1kIqmG0Z9L7WNQaP9Mdya/qsJ742e/t1kqq23
Tn1YjnmEq4HTeHzpB0GfRCztSzRyRLoL9efW9DYb0ZWOBVXVn9LL60krXTNa3ZbY8VdqiLtR4pof
tx6orhwiQg7HxMMlykeTP+QW5iuhBo3UByknoozv2MD0SpgXBDntAfxpv7WX5Pt8EiotWo6WHIUQ
k3ylnLxS9KaoaihSSlQ92IapkaQyf8iH1jXO055kdL6jXaQH02nk0it6TpMEcMXEwTzYPxEk2j3W
IIIgkJdQcqD5eJp7jgkIySOOdeEXNCR/MYCnxxwWBsmjV6QzK19+ebl4HkDpk/7fRGH9uUbTOdXi
YlZOt5CIzAI9a4hQdoqcsN2i29UkIFXe2rtlYpokFcWXANZbD1ivTE+MvSKXY/t5RpHloW8Ay8tm
equS+9UXgzjKBxP3nfOHmXYHo5H7PnQiS6lATjd2Vq3v9fihBe3IBz+65BNiM0fXVWAEsgqHCafq
KaKqCIMSDSB5Po/OEmvBH5mD6ZKtJyUx3oDifL0yg4KuQFRqxDyktimN0GaMKMX00STxaL3lK+Bm
b1o+D2mmqGW4kLvQhq4B5hmKfCUTDwyaQvUXAftQxO/g8Z2mts5sot6LEZogH+dMrjF+nTGEx6ix
167zneCzuLcFPyrKUjc8xkHLE9UmF7LPeYAJscqZi6Oahrxj5ukMzbY7JLP3/S0EHOunZ4TDgBYv
CtpDrRqNL2vD4qhjT/MMI240D+4bYBQrG7lVLJFpnMwIV8YZqJWasIvzOFXTAGl/Cgv/q7qol6cA
N0OINbgp8W1v1w0lZFLAtjH6/MFEb0hWasfBWYVHeSHGkKN/thFWJ46YKjh82dSxmbXv7+Quee2R
v60MO7y0HAYXpwjn9s97HXHgl6wBdBxwj3PerKNhPP1LYSzgauQEO8stfbW5mjvvE/FE9Vik5uFT
nQhpZuOcpdFomcdSr3DEw4pgAbyI0KAIuiISAdyai+GlRl5j6BqBv21qI7Nia0Rchr6kFKtMMFqF
GKPnVELZms4N2Dg43pqH4jwZnspdKJGXgv2hIXPMXWBnEmPEkXlR0M72KzlcvIp/CuCSugjaecyW
q8YEO5CZ//SwVj27bGfp1HkcrmoVVNTM099OP5LAHlTBwemlOauRJ2N4Tx9rpkSmpYkFuw/7ZSZH
fNDEkdLo9CqOeO+QORITIa8OpVtEmyDwBYGFEsy0fWsNWIz48LyQTv8GKsWwJZIToFFdVubYLYaF
wl4m3wTopHgxZbJrPxUJeEMN5Bf8Pnd0cGS6C+pFyruNQsX84fhKOmMwda8sRcrDYAbFMegeJzLX
UmCTZyY9IyCEYSkA/r+Wm+FSO70pUXPCQWGnJ0bWEfa/IBi/O8QVQws7TclEMDgoR0BiSfjewfOD
pK83YMmDvkY1jJjiNGMGAh4UyS2Y17RGjwPPArYXcZmfawD7MaWjZIn6EruwSTbga4aFjfG5PZJz
DzIZvU9Pm1brIqHMTM1S9fsZfuNQMMbfjbuNqL4uJ5ii747yv8poaRSINsQ0GCfI+iAtULsMzQZQ
Tu6PqWP4XMAoZG0ie8QjpQ3i+uaA+FB0hqRkG2VZ6oileWHxK+SFA1HBaXdCyCZvZzAgsSoMcvmk
LVL0QjcBKHoiRd3ay0LAFdjncFgW2lbckK0GfpURRlG3X2gBcqPuwKID18eBQwBDBrOKLTGqDitU
n4szA5obaFSdrxh3vRQ2p63ijSea/JpjUMukaaNpbzsqo6NLihXXCaWcYwAx2lKNhRKBPsHXJUlz
Hsnyjccpb3eliseLcR4HekT+K0+jds3SydVDyqniOljvqEiV9VQd2cZBoNGuUTvllpHwG2T88lzh
0nmPLs1CX0ergbY2g3PubZgPFEscWaLSSw77B1A3T8opO7BLWn62mEEV89eJOdIDowpDz68TW2fK
wcYp2nFbJnoEmoXd+tOCpA96hJr+d3dCY2hrMbqwpcjJ92kQkLDyyUZ0PcV+xe8ojVW0rBgWJqIb
o2WbeRjU81FpdOkbOuVntCPrI7fHIYRNg8HHPpNJ0xiSRHQOZi72qWGLCaB0qsWEwN+J+++aTyEh
eDZ3pPQiagHZllVHIwkgFazs/jPLrlSHccta9iQ5Z9vOa9DE5Kjh1W6WB28EC5Z5cNk/fybuXKuO
juvh9sLEe0sXG5yi3xqs/3/ytEsgGNcthaIDos6AURIS7ShWm9uQ8Ow9DGJn1kaAAdEFiu6b5BBF
ysYko5sQFjLaM+5pL99K+1YIR1mcQGvNhm/N3k3Z3sOnsdj2YQRuuF2tzp5KA5uPvMgys880HrKw
1FC7ZkbO3BibFVFxvxF8TUe4tL9/l2anijBdV9IU9YLVVV5/gsuLEJissWeTogGvRU0ib6TkPeuG
YOVlv/xXJLLyHrDhriQU3kryRbxtBuivVwfB6BbCXYgITbxo1TbiD5w3wndtkI3Di24mAifIqb51
dCOQWtC1/UML5tIawGvCULKPL/0ZcFubELLGv596uNkr4kyMTyj9rIf0monHBIrBF1ECZwarasGs
QFyaxaysdNX/FoJDlDeVdM6aAvCzMp45ctzNeYWlq/seKUX3QwlRyEafYu92qlsixXl9XROqdKMg
Pe3TVFV1ItanDjety15/GuwT97Zjt3tz2eZCgKTM8Yka28O25kzrIjhXpwm+4KjSF8qHOHIZQxmN
8dSreBvS5iP+CpCp9lHT4y7O3UOoEveAA94HAdPeejMz/Rh185G082Fsh+BM55Gyq8I4qTsX3y5e
Octsuqt1XOsQQyQ8jtlO7T/L3Q4Zb05i0ovlDe8FYNNMmhDFrmKPjV6W9fmccAtXeB4cG8mzBwun
xtH14XjeaGgNDmOXev0uIjOYcpXOhSzdNUbs7yS4Nzt/o9HxyTVRG8C6rBeHmh/+PNQLe9UgWs6c
g8yHcsQI2YVOECjwW1ZdqIuzVMA+8Mmq55s6ftpqv6gA3mCrTmK/IxRiLKxR4miN+4clnJRRjfkb
UE9S95cIqeVyf4XyDjgpXo8xpNoqTquFPghfMveeGdJvp2TiTsy0xOYn+/c2aGgYIsP18yEmrjqG
CRfpSPU4QO0nOfmOfjA81FRdz4r05PbH9oP4ZxzwMOAz4nBTOAOJOH4H0xVzF3lkVU2Askajrxca
SsjClCJk9OQ0QdFRrTTro85aaE9TcGcQI+shUlkv3zRAgl8rKYOruGxNRfKujGc2ZtQcuUQ3tcFi
K1ehHZcbTNxuSMNP0q6kJQwp+E05HKRdX9EF8EpwBMStQIMcVPUK472Bo2LjMVxr8fcxatS9IRfl
w2lO7NGd8ddcGOCJAqgYRHyNgZ/cN2aqI1xU5Q4gfUFdjSkKBRofXb3Nc2BeYHCy5XwkhSpn4NYg
3aZ+7GZDNlfTcDpefXxC8eRHkLSMNpD58bqx4evrnWDk9aPXPmU3KpwlP3HZPvSs1lGLi/6xJD85
NiRqxPCVJochr92+m9DfHxCcWaqYqw1v1lUO+kq6AUeFHWNeoqLkFMZvsQo9jGyK2cAM1sGhUXEY
LnHKJG/kb6NOVYbfZ+nK/wuPq5xNgIVgBqZrV29wiZjyubJsUegZb+tYvYrJQR8nKX9wu7nRy12s
jBfQfoAPEaKaxXN1G205dvTRQURKiRBZk0pe3iKt02od74VaUbXuVc5g/BBAra0Vrb+fNQYzfpbR
yToN4BgP7dJXoCucPcBNP5P9ugrX2rEbfmOW8VDTgPn3P/F7A+Y+YXaFZ9iEM4PauYhtAb2+Zq0C
wszNIdziBzx7PZxVuaDM8KFBv+nhuGlPn4+V5+VTkW7MuSW9zxAtZ27aCYSE9yFUK8aS1aBpJ+Tq
cDPiVmGEdkaINjzMRT6qhwO4+CJOrv5dOlgzJ88i1UJCq509rYvMnO3HPBfaNe4Fpc3U+W3ZebgN
WNeeR2uBdSGnXPgdqRn3iV8XMEmSGNahS78Tk4X8ajZQ5n2Tlr8o4xMCeLHUVAROVQb0SmGRyC4p
baEyEJ3sYR0y0IFPFFesHg8/Pj3DUXY8wvI9fIo9xFl50BQ+CsYFSqePQT+uTO1Or+rIiPj+UkAX
z7+8tGIzdpk8o6rKgy+oTdTMUvQ44OldLlBoVWOYPciguAWn0nXt0L9K7UjZI8/ltHYWpE2MVnh4
HSUq40yRhdJj77un4aSpCOP6DTc/vsBeX3KuA5/ev4xWlMmx3kEcl1L7LoPSGMAoh8tRePeOlwzP
3bunAGt13n7ffoPKg/FGnec6mbyFcbgolYWXDLGDI5lQs9SaKzQno153e2KQTwoGcxInwuBpb6JW
zEu7LbUBKYTc52ZpEJxDclXUmwIqTDWxQciq+ncbIuH4yAKFkNCYha7PYvM5B89mXkk3goL0uU9C
TBK36jtjnRgkckSVxc5cM/aUBBsfqMCtT8Qiw3uDgy6PsD35HIZ69a73KN+nBphF94b34tc+whF2
8QpXJbdJg5MFCsEYn/w+6sh375jNkV4gsJggss1dYsoD6K0kDX7NSUREB+edmliViL3Ey7PPl7Qu
Fj+UwsOeGlprhVKL38cL2Tp+6c9FhuqfbTCK+g4/0ImJcDSOZDMrIo8M4IwfRy/YDz567vTULSR+
r9eQmd8/kNM+Z6/ToL91WqKUvc99jNvHTt97cRkltFIrYLUDgwQi4joU8creq+fnrWZ5INJJTPNl
trtHO96GowqMy5ooXh7RzwB1tTukylXOpKKFZ/a8ocv+XtLYIzjCP2mkKRS96jH9lWQA1CKGM+60
hAa4KaOYSJWXCbB2ZEraJ6owdAy1pbH3zsSY+nUCP1w3Jjo48x+iL6o3Q9zMbq02f6TR6mOi76J9
u5a99uQksygw85wC/tRyCufAjHDk0kvimwkCmCh4AvpcHfHsOocsqiUpQ3rQRVuwuk7W3eB/KJMM
FpeAWgJ1TntVIghxxmaNxES2HKRgxxEpJzq2gYZN6DiZJBPmtz2UjDZ85IphEZ2agCiNE0iK7pKW
+lKPv7DUM8L9DHk5Zvypd1oAXWXbSk8yCsdCSPraJBou4fuYF4bkuwiV5dn2KlXJ86kts/ljSk2u
Ic9eYWVSn3zLz3lMRMfvFiovKOUuXYJWAMmcChnzUaTEZOsJ66CTj30JU8g9aJfmh1DLYNBbPGGg
865pTsLizmME8ZoChhjAuVY58kfNd94w5h1ZfLNeIgOsC47GV1Ixx+/ugvrapiEh5XqxdP/Eki6r
zhFfpCMXXqdwdsKB+R1vScPVH0sPvMFenxavOBc0IRZmnz0nA60l4UPQdt3v42IEw4Gho8jtUeus
gIzbhikOy4X2u+Gk9Be9mBC2Z8/xIewJewOvdpOEdXIOnqNip9/pchBMzj0eraEv/R3/4QNN2MkZ
8iR5+cOMozGZ30u6E863vb8jfAKrdNakc5qHSXMIwG+yUcur5L4O0+br1QVVhrigA3qTPBI68uNe
uySawennSjeGwYxour+0SvYfz/9UbUD2Aqt8b1mS5XL62gRCVygaAeGYStPtdwPvczZN+/uvoAXJ
p4muHqXFtt0ZrsNNnvoPmU/47PvJdJHtKSX99CD3Pd0f2MNSnVnh5t9fchn+j0m1YinqmgBh5PEy
bDNgo7zvatP9uC1MrdRXfTUHOI6FsS11cZVDprHeht/S/rs3yJKfZJvpbiLuBYKwooYBlaOlLQkS
zrwOdWs4belsM/iG9lRsi7bcUe2l3BifS7HDyu7Y5jGN2ZbEzfSnU2kcqP71y0SpBajxVHiDqJaf
Aw5qItO9UYwQOhs4g0+zlXaT2xD/Oytcqcs7mUQ64PSHMOHQuOTgee6LPPtvosyUfLVp61bNxQZS
aUzgLnQQTtp+wslV8uhkleJRkT41QCJNWhQGYvXIP3OhAv3ewNCRTRIioJRWtOISnspFzOcM4Sx7
TtNeml6cb34a7jQq9/erIbqouYbVHYa/AHXlGo3NPLXK5/eBqo2XgzO4rpEqNGCv185401Qbd7UB
tGWYlEuRLFEK1tB9LqJ1lZ+fcjGwsTMqnylGarIm+TuKfpbYusQBTXws/lt0SUu/5X3BORpq9d5f
3fbso2FocX/QWDJVOWU7wzG0ZogqM30U2QsWwK8nXb/RfYu93xF889WwBwWVkSSU/ZswGbHK+6CT
B1MRX9R4JyMedIfYsfDtrNzd1uvuVl5/qLWylVv7hu5Jmq4oxyPxduiLt3XHOBbNagfHKxxh3M+U
iQfPVtjGEa905rK0XvPpnFrFfOk+QWpZakTyj2qJcsJSFxxZlTE9mX7EgXdeyeLAtufvu5gYwZEq
/WJw9k+gicgrsiwfjEDecs2Ky/zhxB01/aRmbzN8YVIocvuRSYvfCjiszHkgIVjZaGq59zLZq4GD
dSoDSyb9U849v1CKZGoj/whYuax6lAW3MCdElEF7JIngaIqxPMtTtcwDjYZvkheGOQKeaHtn7aOv
RIUvFogFQb4J9wFI3AoBINxNPKCIrFBxU3X0bBLpRdJDbYWpXJjPPHj6jHBdUhcyaA3jAG2hDCeR
+ZzXmIzWoSSbhUozpaUarjeAdMdDm0/ldVvyGH210juysTBixgj77AsMzZLZlu/tvUGN8cceyTbC
cJ5o4BtEUShuLhxIdGHWfMhfyME+AAlvsb8RF0ENbT8A661YHBo9snDHhOsLWybEv6dJQDr0gIFn
dJZUnL53emm3JAFfxDHA5+r/XeKvb3MStR2q9VGfhxcE/t6ouD3aN2xaQzYIWcF/EeIi/Oe2JM61
WHYt/KRlW4NF6FC3T3mDRJwAK/kvE//e1LCxJRDnZxAqQCklF7kfVWLHTaV7YY6xKPsR/llhV3jZ
4WzRGuKmW4uf4qkfFBjw8YT8uKm53Gr/uTQoN86f5MwC9rEzHDJRYOYYT7nN65w802bplfRfZ+nD
56lLfGK/mE3XMENh1bzle9YJZXGVfeCJWZbQjMeeeP0L3rrkKnoj+gDESfSKMdjxRSl3/hC76NKI
Lgksg+SipFV0rvM1aSQSOo2l7eKlh0TjhlfaF6YRb9NOu/CZ9jepYBO/dNmxXnLxSN32rdzFs0Cz
r9E2NdDbwfZadiKpfpcjPN1vY41Lvo4aGGqY82xT9I9wi+RGFqLz9jy42pD2Z+5i8CZwcZkyUCp5
6OlQWoxV5tcOKycYaWdtLZkChHBnQexuTGqv0ipTEgMDbe3Ss5ddBBoCTyY1m+mJ/N/LpckJB8oh
d1hnXSNTP4VIU2bvZiBXo5MK1TZXyzvjoGCSg2Hgzws0d0vfIovKUIl+h1PmUA53nb0EWA7DFqxi
Jt1uLl5EBrEAw0sIelarVBKn+RG1Pzx+/NEZPGk9/NHGoHFeDhiISlZM9WjPHDwTpHHX27H3GoZx
fJxXtTpl62hsknAS/duoDTm8jLzFhiCpldLU0kIJirOyX86mDbXdMiH+P0wiw2p0+fka2l9vMoga
UlNnxRu14wPjuJdzscbqjd/wE1V4SnSS5qlab1yWCnU3OYWJWQTJmPBDmOOWvoIXdCYjuBcO4+W5
g1TqgQitDTotUOyWIPpv0m2LPlRIvvLJLafZB5ZxkuD1bbNvr2gLMSRxviutrFkkoCjjRr/iqEf2
pvHt90wHzzj0SJct+VSnTLcLEv16FCodo8Wb7IfYKM3h1+fEfNDv3PbXIOSg5hwY+BK6C8lzaon1
7LSK3ecSjkDIkGcQXaaI8Y1bAvVSy5/+261J8X3dwpMeODMDv5RX801rfRSpSXfdCppZYP+8MZ68
ZFKlk52wNleyfDXpPoI7BWC9S8gMa4rwk5HD1jvfI33tVTI0ioZQZiDvfukYvEKkLhMpPW5OypN8
nlU9/YHIXLANfQ0DqLw4d4WRoEI+0ymIcrPRVJXTPr65yrjGG39Jbaj52mQb0RoI2aAIJRTrCuzO
pIcol6BVOz7D6Knu13yTPutgaz0VTHTsThxD2duopOpV8eOv/kdFxIncapzLXzZjn69gU8Pxrmes
7Kgl80Q6p8mUiTu08UOzY+oXAD8SWRFRBuDUrlBudAPnaLo/beeTm+Kd/PUR/+CUzMNY8BRMvfuc
SueATMhNptfI5q0KBrO59QzPsKCCOQ+4odcVeC4nMiq2Bd2VDmr9I6GHeNikWL8bGR38LLWYt4IG
MRTWrDloOatwP618v2iMKikmXlwXCIVJpnglMRJKwRNRlQe0gIh56d7X+TtOZ0FqSotvC7PKQ+UU
WJFIjqpCNH/6wj7g1EuuuXvqDdNWFPAQSeAZxLd/q04/gRZK7aktauZzoY6cgQbO+rFiyvVCPSRC
dmTZ+Plrdm6zPWmfOUz2uNIN7w6x5By1PztfvNnwgAI/2eXgHMRMTEzM3x1BqP4M5uRzuWAWvldZ
aDs/gLAefBx1sWjKBs78NmOjaxpFBXXm5i7odDu0rbPFKJn6rR1JH0jJU//Nu/Jhr+f+tEJ+iGYL
cpgO1qUhzASg9DqFpZP4E9wbB68YNwooOwr7kfFIiYJQYcatSFHed02F3bu0cNHp81IfqkiiQR4I
mP8KELxBxdlKRWBLl5xiJ6/S/fQP/zz3KCTP1B78KHDVD359fJ+Lk2RtxgxrilcYlvw4k7bKyVNQ
0XJp3VEE7NKePotMOElMB+L8MKw1EAAXI6stnLl9OABPW90LMEx4PMm8S3Ymv3rFtvb5QcYlgxmT
BJ6PebDo6ybcd5/vpdwDnPPZCw5NOnnSSFxKrf9dLmRptO6Tyl/HPJK6+FP+3EPUZe9JQrzkaZao
j4tPBA96fim5iQ+081ydW/LzVFQtONfjOsjYJNgGxWrOlQh04rSQDx9Tz0JMQp+Zi11dDPOGxcz5
7Z1GdPYJCtxNmwIFSnuL1gFFiUPah9ECYmM3g6uGAr8H6beUJwQvvJbcDgG59cZcVZC7vzwfzWCc
N+IeSDazJheFQAV79oG7YgSGgKLifEhrjoBPOnLuWzMfaLKvIY2VTL/QqXBdlee8Pnbon2gf4ULu
idjAQIg4nXfIFytUb7A5gfDQiC+qLtZJUOJLHLc4ZJ8WpjjjCznYwHhVlcpsOkJOGQC4191i3uo3
PRejdpogmO9mzCeuNBx5iwKlENndnN9tLr2wFb3/D3Aq57bmZJL4eP4A27v8ZbRvhyMYlKCZQBdp
AKBjmR4k+F63zLCC31CbB+okL3HoJ6KMuAC30hiipIGm1l4jcYPux0tFeniCOlOZqjHOp1YKZhVA
6hqAHciZWc+iUz0Q4ktNdH5h2dI+bLyM4l3u5QMrT+EcWs/2FWsujJCrGhAuCxqnUIfIjGTgHmGv
yYYf1dPwYgh44IGq8MN8EdjUZ1AlAEC0uFH7B4F4LdEsyZGhpgkvAff41UFcbxSS5Llmi6ZNa+if
4mmxWrmgfYRgcga5keyX/oWmWhkdpo5JRlMmn9/WAWOhOoBSuuP0p5Zq1zBMsDttyNVTQ8tx1u6Q
5UKFNOObFKyJqYSWOrLLjpaAmAsubwmRoZ1oJPI2KsGhEz2Xn/0xhymQXfNSpdPkwCe3AQuKBONZ
x2ygz5Gx66pjL0Ihe6RthIOkjI0KZ37QyqlvlsjoSZsB1ubTk0nEDqjxBf5sbRYw5P0XAYLV6FKS
9Y2o8Yg41fjBdNHbJ8eeNh0dOOQMzSJfMd/3P6sA/x7QNBSlxPyM/8mIf7bL9zeADG6y3c2tEhNq
iTRFcl8R9fU4EMCA7W37brbmM3seoTSGFT67gLMIokVQNwZdW0OGV2lBQqbWCJIhW2s0O1rHwe5u
LXUmnm3OxUV6ss5BGUdx+i6bwC2Pmsb5C2bhid4RQpmbHTykMf8eWdTJeJWNvGgAgUQ/zNLjh7xh
2kvEXP2RV7UZ01/AU6041qcfB1xmjFA5Y5Lf/vwkVCIyGSm9xU3v86x7fTQOx6ZCikrCrMyQjsr9
frBYnTLOfEx5oZbTPWZY7w/8yodRv0Mps1j32TmvaCz7/nEutrwVwTylZ30rr2Zpc1S8SSsJ6mck
XRtxvikaL5Q1nyFmCQvRGkTQys/ZsXVKkM0PFEC8L2eR66coNnuoJrbUzz36M/yqUk45uXnUTaN7
9mTzvpCPKYaz4cxzOlDeR3X7wX87naCpje0D2eowUw4NCaEn2naMe7r/s8ZB0qGOqo4Usgzla6H+
DfKzQYAWJwNBJnXusIgl7a8U+CEjMR4kOVUoe8E9AReig6yNpIDgFU8qKd5Mgz/cGDu29gSzf5XJ
/4pvsEks3ZK+lqOplb1XfGr/Qn5gMnakHNHpk/erRg2ex8LVuYDugCj1pczu06dHBGlrArswR4b+
4x+yLpbpNNihWiuHYX5+o1ta75InIKgtREhA3r/OCc1B8KhjjNZvrFDA0Eutdcz8shaBazPD/e9+
JoK0hfx8CMbZ8hQJOTXF54k/bZWv+ay7ceJ5mf+ull6LvDvAjuaDu7DzkJdKP6sYrtsUHfgieg23
wVr5EE8ELJ4Wwzcl2klonw/9XV3Mupdec5AMcR8fU+YczO2v5fJ0zzu8YMOeVpH0hDCQCvgVT9KJ
CO6k5EzTgWBAOTU0WLoJ1MqgU2QbGIq7X/CQRUM/nFor1xlECpU9D8Z4lPkCBdF6cNgWQtp5aL6V
2sDEamUwZ1C7WVKOZNHqCnkA9PWQIDcOqO5ql9Of2m/0knKvKUdvSk0s+IDMOfQZGIgfAV/PIMnM
I/vu0kL9W19+Ku6AxWaY7ubLWoBriYK6T9s/LLja0j9xYIowvgFXIOnTW+Y5tWzG6ySEnDrX8GPX
YB51IibBV2aOVnztg3YlhPK467rs66HnnQ/w37UrSNQg07ufTGHEHDkg44lYgNkI9xrA7LL+3dLd
+70PegWgCx9DVo0CmXRH+4iXYrQW1zv/wASFyWGEncCZubb1roK4K9o2UtM4huf9XkH9/UUe+NFh
AxacJmr4EpcuRJHseMbbqmqi7eQq/aG2dF2lF/AK3eSfIUuzvDfN2XWeH1n2oEoEakZJO9KQKE8I
AsWZjcNAoCOPAhnAcvZjo8BjXo23RXhBAP41e5QuNJOGUfoYIupYGAgaL79cqPZt0FpN0UzwXlsB
4k6I7Xjz3zlnVzGcQgxNqz5vO+y57WIbQV5/JfvaeIkfPwjAy2VoL/wrVvYgAtBbdvX49K2vFZIN
VjmP069SedEXD5+4ga5PJSiFBEiN5ZZ+3HwjIw89gFWi5Pvo2/QodZN77DjYSsChm3BigvxyNk1W
QfMlvfo4dTO9r3rQVtdwXlNRAVF8OwYEVsBbxIJ/iIu8OZTfBrvFfRlXKNj4SRgEa7WcK5ncfRF4
qlZ06gNS9QT8G34wzdp9e9kpWn86RiXeEZX2WlUn1X26GSBYKAC1C/wWAPCpwBH+V1eJY/QsNmrO
xTppj1D4GbJFUwXA37wp2EsH+LQ5S3PwufJIHxcCLTS2j3fmyPr0PNKDgTtnH9+lOCXcbNVg7wOW
SH+qP7BhGihiLIkvSsSD557dFf04VrFmUBrvWFOB7HHKRaYdjuIjWJA5jNn3oZyErgzE3+3ccWws
6d202NqBO5seHkJlohe+vTtFZdu5HZkOA4FUXomn3DXNDrAaiV0Yj3uFP+2h8X4V/qtixe7bonaJ
iVxbIhwaP/lsS1zrgEAJBh3tT3UH6nboRMtXoZgdCOhS1b/Ole+qNX/BsvK2wc0lbSGxIcQyvXIJ
pKXvjUW40C2nmu1FG1uw1MqTGJf6zMCrSea4M2Jw0BozoWpEompAvvBo3sT2hlhJig2urS+BzBDP
g0nJzN+OaleT7UKdlb5s7qpTcj9gUHH/6BRl3X2E7SDzNOh16W/z/PNtLQ5DaulD8YZHwopTPfag
vgBnNb+fWIPULgjAxeYULOHmPsF0Ch9M5d3bLnnB/wXeOEYluoB4KW/cMDxw750mO2IV7Kx2Db0n
cB3cWZ3MA/L1B+bzqlMt5mpj8MkDlai+TXPJo3hSSjgo/tmgCPm4foZfkX1sodGeDhxVeyx3evjH
XVsOVPshirr4cTlQeWPuABX8A9GCGvGtlMmiZGr2n/VL69K68L0n18oC73FHz20Y9QtT3HrUWtSK
ZyskB8xKnvmSo8gN5bOUwJuwz+7TxI8tUQBNa/fQ9E18DJVxztZXaujiBp41wh+Sg/eI5Y6rCuMA
vARnF6qG0rH3ggQe9n+PlZqoQrIfUYH/N7cnlJKuszHGMjfjFUXs7kmUmi1UQS7YXih6VG/H03Uf
ONVnGJHR9jTWD14NW2sDlfEgXPy6zALhdDO4vSduvlCBgsBsdIZO4pyzJ2enWNWQLCUvRs/0NLoj
5zTX90BFVUirFE0+xgxGR51Ko4WMmid0dwP37pRKpexEWRicPZMfqO2AMsKHS4CQeZy67efSrdpO
aC9h9r9gH38UnjQ9eahHz0sC67h2ErT7cr7Uhdny50KBMU1vxDoGeIgpirayvIGm8kVzvlDKpam5
AZ1+hiCyk9Z8WXiBQEeQfOIIqYvcyKGAgVFbFfrXs+5UxDjS977ckWW2S68SUsnpFSi0lNlCqu7h
CfEA04oLKyjluPMJZTs4IL8Cf2cAcJJ7sOid08Df0sywUqZn0cFnfiadldvUrFZ8UBRqTHbyhfBL
ZbGwztcXR+kPRrxiLqiP4lmkahUlHa5n9+SRlKPkrQXIB0vVt9tJXhAxSPfYZsr6pAEFPakk990N
QKaHym9b1X1HGf1UnBeep9VunDE8/vvMVf9atkpwpMvcMWLQpshp4srQWhWwEyc5R7ksEjMMtc2F
gVMhgIActsTCJia85SBEXpaIy9gHXcWaFRbR9Kf+7zHJSOY/yuLb/tucp9ap3Q6wdHhox2NWFjXX
Qy12ozrA9bwYMYPcerok2F9nWe8UIXiCbP3cm2qb0Mo/OXjJggGyfjLUCAzu4EsHZksk+2x/88zL
qyUe4HeHUpfpNhe8HWdvLEKh+GovQo49bDut04m+ZNqge5ayX7GBCz0MGFX/wwDxpueiilQZhaMZ
PWmqTQSyXhBa+3TxGL7zXWJh2P0WUeLQf4BG07WZqO0bt9AMU7tkcp/n6A4bXE6ch1cwucX+VwTG
GFHllm33yCfxwVUhcvjeXey3xxZZ1BE2HvEx/6cYmL/fnbOgxCF8k2qxIXRraDXUyEX6jwppIoVW
DrpYzpX7SY0skwWfaR8RmRUHCTEBKiqFdPcEuBShRr6E3/Z7BiEeCxOknraPDk4gXZS8KU723Bsn
HMCsHN2ZUtrC9ptQairdgkZ2CdOa8GaWrHt+pCh2BABrXsRQt9+zwd6p0sLknOAgbhsJokLJSt+z
kngU6+N5vkiO+zjNJCKfViOrtO1BdeUiYwkhstufC6tt0k+BfiofsHpHcoXQq8fTvEhzFCS39yJc
0B805mMV99ykhRqCn1T8mVRnCCe4eSVpoB4Ne9keAR2lKwrhV0YTfDapJUACMuNlV1M5KBP/bojX
6em58fL5ms05dmaHp8ATA7Sh8ikH9tf4EZN1oMie0gY/chV+GRwaWgK2oNhBjAf42Prk2SGVNOOE
L3e4KxbT47kOHo0Xxcip2zLbwZIVkFc0UcL2DkaCT7GvLkmVUr2NF5b51Jjdha0W3vjzaIh5/qDd
IEsMcfrR189X6WagdmSB1rdoN6UgoVKTO0FH1lOvgH+fRvb9jdKypLIinPdhZZvpb5br2OqIOa5N
GkXEw/xrHf1gYzn3nUmms45TxDG6wBeAh654LjlU4OY03meqEhU7ksMd5GRbUtiszGfJ6vsGenPd
CR9FBLcbyKel0JjMLRnhmmLCWeb33monDQOd1n0Q4afIOogYjKFXdIB9uACxhFQuobxmBQtm/tPW
CDlEzf/c1J0G5mwPPgtxVVUW04y+jxkSh/66d90KD+Oak5xbTdJ5eeaQp6Sb7fEThFof9O9N7YuM
y0WI1QpneLfQqTLG5/QaIBqJzm/J/STE83JNmG/4uQxrJbnxsqPNbCjlM86ZsUJhmU6uMTFpHANO
eK98XO8Ug1ww/TYoCSqxWFFn+dnY4g29ZYCVxqXC+Id8He5aNm2BzrCq2r6Spl86UCVMwC5dNSJr
oHhoX0L7FIIXw1BCjMAA0mrPaNPRtvu0XMo4e+Cz1fz0c/OQT690tfDDnWuDWJf/SR3lFole+A5g
nAqIZdBMkR4PHPh+SqrJX9QQGBhUCr8Rl9lsbv2f3iVRmnxv8DVxdzZ4kAak/qZBYbIlWIt/cfkH
KXzttkB11VXa0LIGHADVft/OPKsLftqeiTQsLdlwTrWftOhl0VhabLjQUo1cpLJ114x0++9Sx9DH
F1gheOIgGGnjEfpts8oaE6q6jiMXyKbhKAiyTotqPf18YnTSltqi/KB9dZdRsVD41bu0Mu/cEbDa
K/OPNp0BDjV9tV8C5hyDhUyc8JE2G36rHG0JISe68PCu6K5s+gcTsxmecV2mA3X8lBDl6ERMgijB
ziQ86EUhv7ko4jNL4+a7jcTpWllYEgvfJRLf+oy4dAYEDqKoRK3py67MRMoCGGw+Rxt1RfCUuHui
zatGW02HkV384n7nAdDX8DQ0IOUOccws59e437SI9MW9lYjnMOGRLMnpeBQFTvENbEVBdxzkCf9B
j78lZF2LMbN5Yqtl1ZLbHebdjii+MKuHSnkiTBH9R8q/D5LT//l5z5eKNXok3Oy1j5gbdYTaHNMU
xALG/rejUOeoBq/dFDUoBIfjnwTL07+eEbSOSIimD2FUNNkFn1vNVxeqPBWtknklnviChHH48dMA
JV/UljtWvXo3VFnc5YYEl3/Z9B8hXnE5Pi2gE654eX1hnuDH5m426dJ2qXiP1Mm++13LtRBS1WOl
72MJAHfFpU0hRRpQ0bhcJeLMzZG/c6nbS6hxejcsW9FcERzPJhgib5irHPWrZhThYPzjmUIqqqIb
TJh3dPhzBfdYI07zIhjWTGmOYswKWg3H0rH1YO/K7eQbEOWD04TGYP4s1TtHkxSpGPMwoBDtFLjh
Demvm29+gvxmL0uQGFEcSCmGy41Mo3A7KUoOhtC7nEJXdQnmuqEHgHkzxeoMI+q/Vu7LElRnYa59
LBxOhqau/i2G8/VpnmJ1BEMem9OvakDTAHvpgh6XzYZZpf2bazlWF/+0CHpPrYj3Rneg2eOkBq+D
xdoiNyPhFMU1/iu2YS6k5c5JOtpo+uGWvlPD3MxKmfe6R55SrdFeloLKzJPbRJuMtB2F7iBT6S6q
4h01ex5hHlBXyNcGb4J5S+whE21B2Y8nSCFYb4CDLRL34/UnqOObbbpUa5WHRufJO0prHYCZaIiZ
VkrUIWxagsZfSJ5VeJT7QV6EnS/9NiIC49rUlF2mqIv3ABeHTsNpkUyXa5PgCfwRXQ6RrcLQgghO
imhwIQNgWRFEdPytSkahCDWu4H9rnQxqUdxA0adAeHb1dRNY2X5+nKk4QR+/58oQv8dMKfwwUq+N
Y/J9wnmRvY6p/0d4y0LtQFFfPgJvOb9siTKgUBFj9JyqnNYNDhcmtZUrQtC+/aR7JxdQEfkZnpOk
PZ2nj/SjNR2uS9eTghjj+w13Xkjl6EgR9r0LmhYCC9w2h4+rZoEbdfct4mvcMy9s5+YcjGgLL2vp
F8wZnv6/rZ5q0HU7cuwWXmvjgjXnk0bQUlL+G8HzRDV0TdAH57I2yPsDMslBFdqqamRgoYK8g1V7
uC7mqtsKbkuaPsWLyJm6NfvPVSwca3gSqjkfE0+3n8z3zhwQ1A2c0kdhzN1pxBgyDC2UYr6fzUfz
lXEzeGMrGbYRDmJ2eXyEilYqD7tIrC7v9n/MnGwEKONdNF79pMNjZSi71hApQ2KRMKpBDmYTIS6m
JX3BOtBEuDF/aNfcBLZOKibqKW7vavpNHYFs3ijJjSvtSF/CJ9yUq/23rR5Qoy/D4c5+epM+t6/y
WD2OhgB7ak+bgMcwkjzH0SNPiX96c/PJgc6PkTmsj3byN21xFuF+GAch8+v5E0Ql8Ikte9E9i1Qm
oXnYM8CVTyOLrGi5KlHhac/oQsUVAlDtLh/8lUiZAPDFpOX8kLVW5fJ8WiapLqo6T06bQU9D2QFT
EoTD0pmcp5YilIF3UvrYdB9Tgpj7LJKRgQ+5JmS4vkK9M89W6F2ZPWq9AIoqlCu+RC2Txi8q138C
m1koEBiJSqsLmWCeKmSBhystxFPkTdeLbBfiXzlUvmrcBcM7ca29TWycsKccetB+0FDykX4Kh7+v
Z3tw4kSU54w+eKz4n0GawVBulAqUXXJn+KKVBXb0foXIleMNZ123LiaToJc5W7sPFtwheRGOaI1W
Cjec5SPM2rFQvIkIDKZQ4y5j2vlAeRJIQhpOPel8qDdTPeVR3C1WrCpvDpOvZ2sBSngyhI/mlKPK
62Yykg5nRkjDqLrCLXY7ZGh4JXgbJuOBMyvVRxBUIaP1Vdd1YwwD3YBrZ6+hV+6MTSHnmCHBBimq
e+XYUOXAbXRVp9DJp6S5r+SCtJSBE1lmpjnBEfRUHOM6sM9JNcXnHO9V0nMPFjtPvs+qCxHhRDDb
TQmiqheP25r8R3dNftfx4148C8RPhJqoDx2NGjsQMwsC+XpC5KAbb1F/JPFTNv/G7OBNiWcEhJEV
K787uzk64nd81XvpcBe/iDYoo4HHWQIRP5v+2jkNcIcsFdgk4RbaUD1YXXmNklQiLFju27jt3krm
nbHvwlmIlcefWmsTv7ppY6NXSZP9ctHRVXAYEL3sfpYk9UpS/w8p3wLx6PTbzCDJplot+avDjrGm
/huVZrA+zvegwJlXLX2JpSWmB0QVpy5tFlt9cAEBtnarOqd7ggFKdK7zoAbckp7chEkmsQR8TinS
NnNseqp8rdN8+lJVvi3GUQ8mxlTI9RCzAd74qSFaaTjUVMobXPP/MTjU7pYtw1UWImwm/Oqeyx5h
9oABY9TlxonMgNuQ3I7Yz302qmoBJcsfeEmH7/8Ht050IVQjRSalc6EuFgJb/uROPxcFQv32kf8D
LFH/ER/NIizdw+I4ueltkJCZ6btgRe3f4S2sNytOq3ARpr9l8JaeV2myDyUx5dqbrhLGaV9Cdxbx
sR284rGNeTdkL43F5v5w8WcI1pQR5ZHP2Fjk4QGcNle90i8p+OiVE51lK3+vLDBBWu4UHK3n60G2
3vHLn2cj2YfhPAUsEwig1AWNBkRubQav5YUrSeFCNPRFzgWz4hLjMVScCyfNbErlkfzCjOKCdYCR
Zx8lh2pQdVIYf9tH3Cc/s7mFhk5b+5my+wJ7RbjhaqDx2P3H70jAPSH46VIw0zoM8ujRXrM5jMzE
isyGkafFKJkn8hYAuaVk79FjwLZWplUwRnnltFesxUwX6tvUbIRPZATf3d3JoWMpuE0jecOhYseB
QoB6chmpnIiPh3h8/bGJN1i0v6Wqj1sggFW0rkJriuq/4TdUKJXhipmmg+YcgKW0QP7Ol8uZSri1
65k2GOazfqHOFGISabzWKDEFMYyBwhqtszaZ6Ii7dRgOMgAqupYdu6/9Cz3zXtuqnW7BckHgNoNa
5JZYd5Ysq3XLT805pPzbxVew3IiV8nlTYFzT35IkwKLXsLh+M4gUXz7CtpYm4s9ycA+xac3lsjql
d4uUGKOTa/QSbXf+Yt7NBuP+/sy+RGfhLr9WZ1/0mbKdUTqp+klzUgVqXl5T4YhczM1k7gPaKdUB
O6zFpOlNCz82xNK/c0Q/cFbmtTgP09nAYIHYRejl/AB2R+v+XD7OQ946AE1psmRR4YFREJlEG+yF
bthfvojkeeIXqc8kiHw+qMTt6d7vzD+XlRrI1n8Y6IaxvlMLB04ZgvGnxZVLd84drZFos4AfUY5I
SVgyL4JnOem0+0xE/iR6C+9Jx+U9pNNHrg6QTtS4RqOMETd1h7o/UAl1cea0KRaeobulWm/ZUwpz
7k3DfJHyjl0jryiOI0ImmX7t6Ik2CLOXF7eYRiAVOevV9ld+qnmQqGE2PlHiGvLdhKEGKYUUH+8j
ieHVxRaqeCp47zqz1myQ2gaXE7aJzF4OZomLQOilcPwhjtOlJ6l2PKZmW8Zm9MdUYRoeM6+YB5Di
M32TS/yYuLNjXgvenNap2u3EAs7xyxaM4LC8jpqwGDfN3v5dvk6r5VHLsb0sRe5CWxw78fSP75Ns
Z8IoW0cPps+GBaio1pzIsdqqLCMXblijGKl2nFCh/Io5aSscmdWeIlP5fDKLs7pEXpfvG6EZwCxB
WvrXJkm6bd9n3RNqtjgAFxqtp1/nflckevG8K1HE/NI8ACcsw4BBnSQNxz2TmgxUAwBsKrXZykNT
qdI2h95ht5HQ/mrodHYd/GXkDzcZtjwHLSys3l2HHYAAruam7kK1XimgxwBnZ04Y+oOhKKmizwi4
YS9isezGO9Fi0hto7OeHUnSRU/I2s+Awr79ZoMvGqK3agWZJmtqcFb3TFsckA/vX9y1RkvXnwtaR
upjUF8cMBRVM656/DesRVzXf1Bjkqhs9NjdrGD0s52l7mYOL/yBeuh6gJT/xTtE0Z25+lQkdakQz
P/8UQLihc2gy++xMr5GSqffmWBqGMKbJUz4QCXDhKjG+zPXb3dClqlY7k3TAVwQ8JGz6lk6fsEnI
r3WfcX8NDehCVqBCHD9MC2Eh/VJkZ5PzIn1zG7391xFyUKOS+aIT7HKYrDkME1+k1ItKcI01+vgV
5TRUDhTpuXQlMzZYH36Uaq4LFfcPmdEcOU81gtOAEjF8U7PebmFIjVGDmUrJYSIPcnPw9usHi19e
E9qERlZTw9/Kam1TxCPji8YR8WaA1DDyqXXt4rLUXQWld2DJI+Aq28Cp/edbAUONZzFsSapkmcrT
8Ia3+R/7umFFaDmkcYel6CpV6daL4XSgpWVHztzIcnIZOZdc9CV8QpiylfvNc6VZigWriS2DhEHv
Pe/8GroaOZs6nbQCvOso1QMNlQw1o8xhB45O7veJTNDUxrD6exMTZIQWOINB0n3G2W+iimadj2QZ
706TS2UamH2ws0wKQ35VqLry/g7XekL6Iij6SZyj9Op/EtmNjkpzFyCjecDRmt1eu5iBKB9fHcLb
3GOgGLbMYpBgOXnpPm1+KHCufDEr2dcVerMe+firlw8Q0Jac3IxCRQnboeH1RHcQSCGbdR0cqV2P
91AUAjVUoznxQOocRsRfARNiQupZthrWRqlYkDb+YaE4mjiUonlEr7ClR5H5aXh4qeXmETrKRv4K
Sf7BxRywdFydIuHdlk1FOAtM8H/hmarvvSsDEvlP2oKbcqdr/NU4GkIjCmnvYF/mjyl2VO3/og1r
qI3ExhstdIt6tbMcdF+J9qiW1lO/2rZ6h7DbGnmJMmm0XwwB8JtOTQ8Tu5m3/5KytFFbt+DieNoR
9bGGm6UqW+pX5x+lujiPoVG1p1V5tLHNrMZpG1gbLVu0QxRHd9wd7tY647JChUKwmrzEsLpG5VHR
+IVo9FTbSJV/XL4alLWbxMFoC+cZPBy01NC+txALRUMiv5dgbAELdighBbJfNL8hevR7b7h3befW
Z7rKRAL+2NI+aKRLpr3k7m/zCsSnhPmXs778Pyxg927OjX2ZBB7zQj/+KrNn10C8rOBXCvpGIgq4
zbDZsHtpHXrZmc9SeEe9PhOutkoffeUYLeEnCeMJUkwYRjbSa7gtR7H1GZGMMEx6yuwu1EnQ8+Zl
MNMh+HG0kOcBdZg6PZ6tAJEelM/UByekxc7nOcVcO8Q2wlMy/PvD+IkteOOVZWZY+DaxXaop3sT2
0wQXugfGq6v/XtsB1qjWvpkGBbG/vWBq/3OqWq5Kq44kq8X3V5Ph9riuWzsFRxquqBttzitAc+HW
3XMGV01MM9pXgZ8fa5INEbufeQbCTYiMAM2E6aPkAMyr5Js/vO384H+DRlbBsKBbCatIh3WYfXR2
bJ4I/1Gn/tmFrc1Knp2Sq1fWIfnTRc2ubAJAfZsCJCwlKa9BWCh5O9Wea5+OkurJVEuIUV9C2nYa
wB4WylzzYgkLftmXlkC/EuFo6G0zy+F0PYKo0YoUJpsUiu8B09a2QFejz6lpFn9xNNJG1JwXHcOO
z7LBPht7yo46QX+oGqxbea8BpFKZmSGD5CX7DpWobRK6/afERw02FeQbfPVq3nfwlIEL/n1ftMZP
K2PWNDvS10equvTIi68WPzJJmgGAIUbQSnBdxK1nxRQhZHs2nBe1ENK/crK4qfTR1qbLmnjLyKDT
kGh9rknl8bwCicPyyqDqe7/oGilafWFsa1xQIAtsnkmA7VD32143DVLiN/Ts8e/f7E/8MpFzXKhP
YdDXvloC0V/0N4tzpOXH64zjK8GEWmLC69iZx5WkPHJ6BJII4vgO544SvPIEsPICg9fac9ERcGOe
I+uNjmmWGBQ7UpMHjgYsxqFZ4WAE5RpUziOw3eVaQHR1Zne7NMEMbk5AOxA1nux9XXvWm0JZQejA
MKEK/QBkC7lVNwO/jd3jUUhw5i9jPMnaeSRNAAmx5uvcwOF+nY0XlLgCrIZPMQy7bACj3powbxkc
zsFh/8xkcYiCAlE0T5eSVGOn+EQ/i+hOHetOUiVAZ3P/WPSFq+YkIcf6TCVtD9YiW6MA4Y+grW4F
vPjC6aH1eM9ZwRgr17MGMFPjrnBwGxzTWerfGelpMsx4Y9J52W8RBnDmCPhRsQ3FzbwEfMvzajRO
fkWMSViL4f9D8obGT253EUdaRry4aNaFPy/8SgzzN54AyiVZdguFdNclA3kUbjgISEKOQtm5aEgz
+iwZ4yAvQlDkN9VitGLFXB9SDHPXV8YreooPv9zAJlr8ckgRhJP9FGVCf+QImGg8Eu8PdH197008
m9KM3ApmC2JVULAvkOfXBa3k1bylPtRBkKI74r4M6JpRFJ1vv96I36jPeNatANpWfTGnmnnwXmol
8AWc9TukPz5kFiofXTb8o0wSeQ6+itY8QdVO8H/KmlOHcka04hDGszDV+/IRbMMhpFSf55NmEYrf
ixu+GZroC1CpVaLS6XVxSFKCB4XbMOg8mOdMdUxgjGBznBQahn3cEF0lgrPPfHnO2AE3XyUF9Tuj
NYRTireCmW0ygSLyps4fFue6UVUhjTYQnnd9kckj9XkWhAbyzlfIa2vTxPexKU+eCzPxVAdO7yHF
Xqruzh+foPK1W2qSiF/sDeFOPEovDGZ+6uJZFM2RuEt7EDJa55lPXVaQXkXZcKmWXSHAKy0gCkVZ
ejACrCgWO+5Hwtl7kd0a4bmMakySPRGyZgk4bXghLsV1yHxwCGVp1LKJp6Fc3dbcl6sQsfk7uK+y
xrKZWQZotEC4XWH1qAhsrEuLAvqCitGrbG/4luoC0BwZEN5bkYJ1QuudHMNN6494B+NzYW0rJIHK
42t4iLd38UsGYZkMRUiNELvMCnnkJqFuzydv7LKqNwaAf7kderKoMPE8sbhrNYPzg3P1I0rPK0wo
ITaRF62sjKzMhBZ6iqgSA8VwlISDkXuoSDAvVi0JNvBZ2ZaqW5TRv+ExbBV4IIHwwRFECaSbsv5H
hIRmIdOwCBAQVQRPnlluN7Ax4eL3HjBRIdElwVk56HBbhEMlxeEKAgFquIa4BLZjTsGG272346oY
o5XjkuUn1h4wGMlh+uZBFc8c7VTcR6X9Etab7kD7J533YeXX4yNPcAEbzxwHMUL/xV0kMruAAkmu
UHfRYh84LuJndzLseVmpOyugpVVcdyfeLzFtNx9rz6D5vXJSHUu0kryxAGzD51Dg3kpHz+ZRRgKL
sAgJuAP6h6VcqKbXRepZWN6Z+CmQLQrLgLoTK5LsFZEss8w0Q720756u8Sp8ppmk4DV+i8sAeyjb
Ky6iG3AklKOg+WenjuNzFn7SElKrYceXZp2gmbT4rpF95RZMT0cgviFsnfWe4spPBhHTBWudw6ng
ylhhF1GRNeaBnoVKCa5kusYvPx4fmeRR52dKFbv19Gkmvz4LD5tEAP84wu0q+RkNo089PX/cVk1G
5b+Dq1f8DeVsNoVbynK7gtBBMpKwckIbx/ec/4gB7kdhEwSRG7/z1eF0E6JNEcV3b9zz7KMaTthr
uGI5YLuv+1Il9tyr9LIa79uHA0AYuKU230WOdHzOWe6e/dMN3UI/LHpsDIpEtGLjdJQr0rZU0bW0
dErPPOZ0yLwMON8j0b5jRdHOfFUR/iiQnKkkNSqS+wYtARv+tZuvGAAPg+6YZ+OaRXq7TTrqZrVM
6UBL8u24x+cZLx/y6zBRWwceLbAtBkcZFg2G6I9NNp/Z93aw/3L73A4M0S9MzL0ktUYGJL6FOxqM
nZYJsPKHjre3bzyeshESUWKlA9cD8p7L7Xuw6HzYvogIqVwefKcq3KR9yqgxx4CYhGWxQzYyLQPY
awRCtiTz38zwEGs0TDRP0ZJ3TZ9mI0hCHDu+90AF658EOny7WZd15vIMeQfiykV/lPj1l+Lfay7x
NJBfsZWL0HAqSsHbX1qXpGUBGfoOT1zigtmQCrfoqau0/8caNS3IJwWHk6Y12xrZlwNogQ0XMJAG
udmeOn9EYabdj1wMTtJlpYl9lMkHewQTzJcpe6jZpGL6uGBu1QUD+9hQ5RYtBLjKsfSCOXCW/ljD
2KWDjMxsKZdlkYjfQCAAnbkAPIq9MzxHaJyoOCZejwXWWXSu0m2vH66lAihxZ/xqrQu41c8z9Fe6
uo09/NrYyvbvH1+6uFI/KA1F0edwRCm1wS3QGtyGMnOsduZC7ILwK55oJ5Gqj2xAebS6dYRtrIBI
CQXTXUTu88rTl3+xbRt+wRVSLZpc3klOrjSNc4yX0ziDADtNxfZWDEHKIy9Sw0xR2jMtdxGCmVSx
Be0sWyC02NbgJTQ2rEj+0XrZm1lcZlDq1rbNxabsLoBgiazwgFdowOHfPdIFPnEo2KES0fr1LgOe
ETt+7wvlTqHxv3P1K+4M4B+17/X9aMLNwTPo7F5KjApZdPJcWGpbtAO7cFdUYlKUJwsD/szB/4GR
qVeF+NlRx/hv49l9WQ2JDGjlBoqmTdcHb5svXcTlXC/Vij2IKjXKvMgUXW0ZZv/9EFND+F7zF2u0
dgUZ6vMSR5ziC7ZmrHSc6inmF0zc7ZpgFTzVcDBsiPELH2SOLoAPLlv4HYrkjnUfojAKhuPBA91K
WrBkfZECo0TThvKW8dccfRs9LZsQZDcQpZOO6F5mbmsiYtZGP73cUtwPz2VEtelpY1C/8BkxqAJR
plrVFtbzB+b11OhqjDwZZnp+RbKJhrvsi4mD7y5au+7K9g10+ZD7vnB+E10H4UuO9UG4N39j0Jnu
Frslop1TIqObPZG2iPsXxypBfQ6/9Jzan1zE2OeSFsIDKdsJBKTdSgQhwBkSmXJHukK93i83UOij
53knz5AUIj5DlA36ekHv6oJa7hT5IsEalXbaCEz7h5ZA8AX8cbNehjDWrFPLe3uiRiFs3Kh9SukY
u3Qt0MnE1ydkkclKiLRc5nCEvd7l8rbt8vV+rb1HI2CmH0YyxJ2TEk3QEMzJd+FXE4D0UHJy0gsR
oWoJGW7AncBjP5ib9mcSw9dEIsMZa3gO2cMF9k503KOUTdu1SIlOvQdfLcpz8uk910sgEZ1UQ+m0
vD9Ga1aySFM93HQ+mwWvJ+elE39GWXcZ28avJkqGU0Joq1HFfSGRaxSLQjXdNcam9b1vO9Wotiv1
cINnYfVq1iIMhZAOP3aQAEACWH13sisR0kHKO1JkB1y2hjjAk6inDbizfGsTNPyisXSzgIc4L7Nr
Ik1hg8ISUX2x63bCs2X2ohXQmrfrFxafXzX/x2X0wVhILQ1dRbkiFlju6zwvvySOul23Otmz2mQ3
urRm1jQmzsRlkgaFrKGE1JPnSN3Fa23INP7jiNG6iXE9aB7lelJj0LCInKf+V7a4Rz8v8EoHkyeu
7n7+E2iOQTU15oe1SczTl9KmFZd2JRfGuA6YsYCX/X+pHegLrOG4zTMrqejwB7TWLBsUGfySv5qC
HwlTqbLg/7GPahnzqJsZeg4aBEsaaX3E9Mbb5pfMGg5zWo43oeJy7tUEyvxDKKjibOEQasD4HfUu
w/7hTk/18Uak1SsN8ZITMraJbG5LOML1HHFwn7wy/Vmtvx4KRkjcN+geXMv3cjzQW3tCWYGk4Xg/
3J/jwPwUojYPgABf/Y/RJDWkNddFiMQo8rn0aPznYCredD9UYbyyGAHZnKmTxuM/I+2GBu7ttORl
tbYCdbK1jfhdFWAybSndsbYOHs7Ef5IBQi7BYQYvrhk6NUevnaaN0ihRjgCZE5+ErjanI20ZiGyT
DYCN99/ufvjA4/YH9JF5MNpWPwU9V5WT34VgLDjrA/rJYrzCoIelhs5DXnaDXbk89KVlTvO70oJJ
C+3hiEFaa4yErplgDvvBJh+AQIyZTb1e+IbaAjRnZEiaTSDu0Rgf7Gqb8Y/gHzAoELdRnBYQA00p
7Kxm1JkTF7lfl1lRRgpfMEBcR1T5VtVctud2MUKDbZQYSBuQGm6dkPDAmG4Pln6zg+Pkrp8Z06jc
V1sDtxWUrGFPGoa/9lBurt1CWdHg9B5UoOmBtDcg6wVH88S9l4Qof6Oddt6HbCKYixEJ6ER8d/W/
9TXbTVOkaVZAtWkD1NBgCqX+Zje4fjA6hXA5kiJEYQ1n24SNiEF/1RzRD6DN0fcWJd/UJn4hcaoI
mdgG1YRjYSF4qROiOQuJAa7BfaOn9Ho+jj/Hd9jw5JE8FIAPU3g1Sq8hvLG/SnlY6KieBG4oFjc6
vrvH7RCpHO882LztuF9BkL7ZFeThqx4DIdgwCsdl8nbSuLsB1z+fIONaJMZfBd22vUmfnGBvA1dx
d6jqho2f9S47bcSCQxtISsiwlBbLXqZHydwC2KPAc70AE+6NuyLZ7NNep2g+7qazoB90NCZrj8V0
cuS1ZpPFj1sLChHIbzWiPaf7TJfQI74W5+1rX0hBMAk2aREnqWdp9jF14hlOUjY/U7JaOGC9y2oR
ycLR8yR1Vwxi6IBXUWz9KZweux39Pon4fJXLA4/aJNmzDdKJi4k7PJepk3OSKXLlJ/ZrFhnMBIAA
tuURsBLJElSqqv/nSn4FKw0cV648cwObxwht/zpTvtWPalruArkU44O2/le9Br1wwJD1tBepuJRt
MLu3kvXidLleVlf6I/wgFSJemmsWbkoqcPkrcFRWG7FPEu0g1+vN/xU5ZVf+iwNXoujUFH1N8A31
g9KASfUs/002y1Rb45NDKhuC+coP9ITJIgcbbwNgcbHTFTmlhJheDwQRZeXf78gmTSmYJizhBFlj
Vh5VTEHvoQuzZCA7r5U05JtbWgcFksEKZGXMBTCgtZHW1hZhBkNfoR9gzZAZuV17z90lhSBfgW4c
2gRxEU3OPg2v7HybW8dIluU071JA/fuNZRT0CL6MqcaoPZlUKPgxJ+WMOc/BE0CEwvG5ko0V5J7W
L0razvbVbg4rqJBgPHVjqE8+o+kYkLQfT4vaXZHTQE23POCDhysJ+8RjAelm39NKzCNX92Ugw/kE
ZKbjU3ZBfe8Uuee1v0W3lzxsyGAA93ti+OaJOOzv+3IvQdsFSy8bCizC6WbEFht08sm26UyREjhr
8YPDqu4DQrEH/5zcgwvAjvHZ1PyCTWBiUGubFqfu3YYNRtcPdacMWWSLssUyvZ7TRyc59JLVDfof
k5m2xr1aolK7HS7zSE1dxRNp/84FBMzJDCZUBez2d0jp8bKYRhiV1UpkGVyL4SRJtzgEiMcC+9GZ
PoFSqXyuzmlrPmKNuX6M+iYDpDsHp0Fvxoe/Rf06mhho3u+qkKJhaFUTUB6iVe0DqR4mWvMCXTPK
iJ3AX7r4FLsywG/v+YUWPZuk700Cq1e4zpUaK6b5LyzwWsp8wG6jhHCL4+4xDPtR2yv6Y2lzQ4Vr
NADXPKWe1D0GglM7qmwA87poYuvMyABNP/jLJBEBkgea0/Bq/3i9s/3FQVNyEE+hRG3EJxMrDmrD
CmEPkcYZx9qTpbnZS51wFArlAoyw7DsLfKlISCsSx0IHm5NMV3uTtxLVik03ayXu5SZDQ3usbnOl
7DeyinUwqLi7rRNqJAWALb+IUqULU0hKZB1Jbca3WTbEYt6Ssj9Eb6oArtFJabB81IQUURn+m1ZN
55Hbd6sJHUUo/TJi4QP5/QzdbL2lOfVZZufUQaWplLLsHGd9Di+W1XIlHBY5ErBqDDiRrcKdvCLj
5eSiw31AVwBIzJU2S6Ww+93EOftwXsnICBG5dPIzaRGlrG0YD+K6aXSQx/pgfUG0EZ8xmj/vkr7h
bAGdgfn3l7gvd5Qei9Ub/aZVe/xg6TN5GaIl0DP380iTZQH4PQ1hckC3WIQNociwUc5syMQuyb1z
xE+4GpwN4IBc2my1hylH4FH9UHgDqpYuKJQmZv4WARb8w8RpolECBjMJls9SEHD7RBKZaIfE5yW6
ARAVt8KecH3yr+9btn02wYfAiZhrLMd6B8ijqv17Cl42KpOI9P1zWE2GnXoBZ1yu3unGfu48+Jy0
UJ3agoltyJO/AObN6QQYgJ7evF5vte1aRISgYr5ZoDS8G2oo7Q+7dJEEdStsOtCHkA0/clQCpQmT
fXdJUJ+j1tgMEKE9fqasUprBxz4ev+AS9obC14Ls1LY8JeXC6xEskpl47UHA45ocdiWlV5R+Wt2S
3FnrstQW0WCOXG0a91c3cYx6+WPXt7nZIKEYoqy1dUUIDbWOwNabe6zeGcqSUtehUoZnuYITxFq6
y+904pwkVZ1LaDYkB++5JMvfTBp08CLPZ6NCoQqJqwnkPHuRtkw/H2WDGkkSGVc1c3D0g89Ivia2
5xFsVfhhGDgbhux+fTI2OtnONyCPIgG8q9RLADFGvoiKOhl4yszCFkGZ51WQwesIkp++2jJOeeU9
EExmbMFi0ltEMp3fyYwJrrcG5uvTFAG9Ai7wmHBqrXiY72LEbuFtwxUBDY+coLgMrXtlEdb3BOM+
JMdM34rZiiVy4CQqrsMfObrC6GLccejkaQjGOgXwp7CurDzTHLFwyUD3JAUzVLyb3CrXzibbwSdh
GAQkNY5RJyi+ksx2V9tbhRZ4j36xU+ZvmvlEQz3UXbRpYgH8IYwc0io6SZ4Hv/z9LofND8g9xBi9
FVlChfvavQDlVcPWJRLXkS/wEPvDI9lQfHe30OX+C9IkZg5X2vLoBNkYBhyWSTfxEGh4LuCZqPkm
SRrW8M3BGiERn6uj3oOtDVz0DU0amrr32KkQK38vAkoG94Y6fbHGIQKYvGFpsw8ZsuXRb/aVwx5O
PvP77Nfl1YPEkINXYwUSuIOl40r04i0oj/pKriuFwZix1MeqnkCHF6NjwzNZ+c0kkfCFDrSVkkVi
VNqH4PCe7b7nWot9ykE1VO4qNErSC0u7Xd5kXS0GIHDFuudK9cfN5yG+zqiX9tLs/TlSC/PzG8rO
Tz+xpeHaNPCz+rmaRrqhk6N2pa17TzkdYpYC4FpUGew8XMNuzF3kxzS3kv8MOOOAkTUxpCik5har
4o6dbx0F/fI6SynXmdGy2FQhD2NAnZaxzMZjjKrOtEOFzU21FUtimgdHcvFAn5XiVugE6Me5H1re
yZ3jB2fxaInDFTVhYizvErzZFzL5/+0s52AB/OMatmwOqgi3Uqd45HcmdhQYF/FQcI7W8v+/id3O
tsayFP2I5VsjOztXp2RV2czjg3gyQe0taLtKKVshwzEN5IDGX7rYIELIj1BnCXEGS0q6mdXNPAbG
iJBTwwrORLjPc6/UXAb7vJVmOk75QxR320Lw6YyzaNztVn55wX3EXdxDXk6Vxl7g1c49MrEhkI8Q
rCC8Q6j7wbuNqXxWj3oo/+4ez20+ETOj1CG2TtqEtVWMywr8enTDYNdPdb5WiPOWZT+qu90CIf6f
5huoQnsduHbG6oieAb2YtcclofFgBFxDFb2sHiBZJNeorMFmj6Ccv7vCsFD8mfJAMF1fTOKFWzSj
plJO07BLFihLMjfMrdGBnJ2dQoAOMKti0DA6LhZhXCge0ZOVhFuWS56bJfYMagRD/ijFUYfliEgS
JPJvrh8sIDVvZoS6brpF58iWrHdyQHyPs+Dc/QCwCIA3W9k43Zq4imnU7nc2+fVSCF4QGAVMORzN
X+TFhZi5eRRHZd/JyOikQ9ts6gnZwYcWzkWFAV1XVG2PwqJVEs7IVyYuR3DyR5x8iMGQmC0OBsYw
97k7Na4sjOHNTLp3fAWKHnIIP9UrurA9ciCRzWWa/P7JNFga/lUNborvo9Z4+MA8bJ+gvWhWRVNP
nTY6yw1iLNEIf5pjFV4sA/BIfUPYgMYs6Xj4wlx6F6g/vDfGl3d6OLzbH20sPKmOGNEJq+kkzbkF
e5+6Ll88E1YOitohPuYZp2MbDM8LrocvXAbottylbQsF35qDekY8fd/+f6CQEp3jiHNmspItAE3t
cViIHi49XfTS+l/ZVx3zTOBhqFCwQ21O5CqXAMnm1kOeyt1emPsxlHZi7n9FjCeueP/NyHR0HOi9
jAd5XN1ojjgC+3rB41C+xUmIyRz47Ovl6WAF/wAc0U/nBhv5SUBNsV369Ru5NmBW9uEdwnJVXsk2
eTmv9R+jXrReypxP4FS498OLGYYdTOjs3ktwCRlpjasM/ye7VBvbizCxO430FN7uaukpQnj2oevE
59yDyeLCtIKGAFE3FRh+LTqW/4rr0X2y91UQgWZxZhrLKQa81fqYNj9E4aVNvfCyAR24SdLzeNkO
Nb+O2N38mHrinl6sDYR6qy+nJ0EZM1DXuO1Gox7G/C9mVM+WawCuyF57GH/8gDtOitlk4p2Ku2kT
/wSNAKE3Jsr5zNAqt0m60Xeo5iyRJqhnQcbeVXRYgUHapuuTwcNGlNTeAQouoiVW3Kttr2Y9hirk
GhGHWtMjsvELa4wkJ/d7Qav/0UmGrsPEHX5ci0kuFsRSpkfE5eAgOAobQ7eGeqMh5MHXq+feESOa
jpqQXgDw/0FRl2VlghzHzj8SPsFcb2jdjJxn/6E91fnZtZKIU+cNT8ySuseCTS3fNpyQMGH4nh0z
zEyU/iW7fZZkcINOgZFpPvcZO3hicuZCtkpk9pJv79DhsW7axBhpAC9PFOS4IC2JpP4+jpNfFcxJ
q7TUlfGeoRxzAFxzoCSsm9D9T6jxK1jgbeJ57kZM5CMeFo2tuKqk7epcj6eOP1ibtbQQ0w2+Qmyi
bOQdCelQQTe2DucTbQrtoAVCgh/9Dv+feG7u13jg6sEXsXda40DcplN1OsmrymGaCZaPgaCshTrL
BkELWcRr2RNZKBF+yjVjNgc4UWHDvyU6j77v0idoVJFeG1s+H0Zy5ZS9qokUL1WHkhSMWaG8d5kd
qHrYP7IziQjxppQRf/Oxy7lbW70mNzJJ34VSeTuW3ChFpUVfP0EA0/uW1iyZm3+sqqPbL6Lg1LoD
I+Q3+CDGMZZGTB+KWlqqGYS4xjvfcCDj5Qsl1KDkvZyIiKfS4UAzuOL8Mg0CLrMz1FLjQ9XIHpT/
OedmNWZ0CaWMx0YLChv+3y7prUeoe2rAHreWhVWHTanod1LGpAyJxZi5a890y8Cit/yDYiF9o/kI
BOpSWSnFQ0PCrg8ngnujGbHm+1suXkyytKJm8gqYxEC/dANeFzvkZiQ81OVubZxRZ4NmybJNQWPU
SlTkLd2p1vcVHB3bYvaL0tXMi2ducOKI4M34Nn/lOvQRgA9FdLgFXqrxBBDnyvNT+3S7VVDsJAry
URkpw80+dJNEzii3DFWqhCURNaNYkUfgtBhX9vMmv/7tyYNQ9fklz8a9QRdrC5NzGU8MJLM2U02p
ouoWET68SfksF0hvlSEnHvtqKW/X8uGESr57s77SwV4mNeVpdUxVRGlCbtog5bZBg4xOcmtHAIJ3
LFinGTeByZQ6ZIRyedRsglmhVF/NmbFAHgLw6cEsRMyWN168UflzPd+AH56lCLHLV/mGwqYHRX7N
Oqq/uA+QxUCeugeMM2m5yBeKyyVdDBB/EJvgk8PU00BqPgLMaFXP4VxgC1u87qHuuNMJa8IPF2Gr
BpoDhejX05tMQ6yqT/H/LMiqQ+KPaYcemQhpUPtVa+jA6eHSXXMqkicHwdKIi2PZ+ywKuSv/tObw
Ur7pgqPvfNVpZpLsA2y5uR7rbF+YKIwQFoCqXn//hhK4DjRBHFXNEwsIG7fCwQngpqgGdV0a8Mpe
yTSUhW/S4/u4KgFUz5NpcYOfZrV9IMcfDMHI096kF5P3UYtjKTfqbgTwnz+dU2UJ+GSNju5pbIMF
McWWXUiLkAAkJ4pWHrYiC3SuOk840d+qEZZJJ/9sRJSkALLJUdO6+HFLHCz0XV/aW2jDEViCFPTP
pWbKhqL+7tcsEfulj52Yttdz5FbWxt22Dcn2XBBJLQ/1dDF+Ncoew+hiLdU1bc4/XTMG4GBGXdum
EKFhYa6CK9pbfmQMvFFtxI9eHSwfmPRqBBYvbjulnji3ZkHkiAo9AOFCXJCbfHVspEyIuMQclWEG
drEFc28z4J5mw/VxBbOI3nNOimtgEgrmIvSes0GTLFFA5tdfdlyLkiw/ooyG2Apoa+XaUW7zk3I2
HbZKpZy83XgN1tR5f3G4NqSVw4uLnQi87EbU6eyQeIPNiJ5tO2Wt54rWgk6KfOEaNJGwwgSDKO/X
a4S4dNF0BoS8gz7jxNUNV+NzRRo+rN2VA53NlEWEfvTzvbrLLvpgU/gQ7nkGhDIq/grs5z08RHJU
skTYyOsL1NvS9YhDoe09x7jJmDL4QP7BJI6BxwokMsSFmUPzXvLzyETysmOW20WfUnp6XGdaZ5mV
m+7TRToUcdMZKldvBwzfWPsTITpheiif8mjl8GD9NKVPh5XbJzo1VADYWr3wRb6rVD6XtK6Fgwwl
vNhkw/2linSlC6wok+FUibdA/DSs59tLzJWG8ikKnAd4kd5jfaMmO5J2Che31sy9ARuxhns5PF6a
rcXTv7P+xGGNLpS7sgmVCG3aD6qp5rQVjWlKLih1IOZY6trWSczKm2QLWlrY6L8afB9hz0kYtkAn
oA9q+RJWnA0YZ53w1FHYbmUSLX5fK1yrGdXBjBL0SkFijdoF8avM1lGyCZI3gYsDS1DbZVM9/aMc
4OZ7iZbRgMFt75gtpZvrQUSWSgAp6XUrR4aGgBrzUppgB/gH8BNvImD2kSWJvxm+7wf6xGRxyTHc
z3eZFzatDa6vtPfmmSy+fX3zU/Qgn0z0Z9RDcJGlrFWSNUE6kX40AekQUvJO4nW7AUG4dFXGPbld
AkroWBDLP9H/t2w9uoFDyK7clb6mHWmoDett42NMQXybNwDww0seCzP6rpDBtxldCXkgDTv0oyZf
zOxaEgNzq+uiG+zSdbZz9Iw8HKcdL15kv4DLqy6gRkSkuWv5Z51ZJExy7IHxrBDG+bK/NPolMRj4
G4StVzUBcYTcR11JZseNl67UrZtJGd3iSnWiLer/QnIFv8OPKpmQR4FAfLH6tuw2jpNmdkzZEwio
bcHsyBCLLfagBuiQsG5m5W7EwEGImC5gyOowy7aH3L5f+lvXE1jpNriNDmZv/HDuLooL2C1Bs3Em
aJ14VXze6UfsLab7IFpWXYzNO70hrrZUsgxjP5m+WQ67RZEpvYvkm7SmzpqB3ftycEh7NEKGF6ut
28g/ysmecoQMHijIh6SrZEnUZdOfKebt8GLnpiapjazE6fHuNM1cPzEwVxz0HY1K5TC/46bx+tiL
xkuBq8R0xnGGVWSW9b7CKF6zd3jmadF3t/BRJJ0NOdCTwE/qNSTooMGoAJXySwkqNfAHko52h+EF
qEU/RvR7bRAYIRLpEe/Tbs3xTJ6qLM+CHLGO8O98sRB6vDmXkTCnrZxqauMOQTpnZv24mLZtPRde
ZS3VcdqbMtkEvTcDyX48VAPJrImMxRxtnsmdzAx9AlwZ3v6YJAE1jPaA6I8rVXAp+IP7zt3JkEds
gPcwPIr/Yg6B5D+IrWzuNFCJrSVmXJQXZb/ouyC/LcxyuiDKMDV4ASaovjJ2NekvxgQsS3xbi///
Cx00Cr7tjn+wwco0jvSk4s1lG1R+ilf+AOGjJ9Or9TCUrx6QDXGdZKqi7XWazaG4zdENXECschru
kBalt1z0EQ2kFPhX7026EeA2A9QiSaZ1KzK6in1UTRSCIj1Mwv8EYO45NnD9d9/yVmifLDDYFIN7
yLBWIkDvqk2BYFKwql8g6Qm3NMJq2abuJpTGk6f+OmJghO3m1MTcNi88yX0PRgpi87mz7fDUtxQP
0J9bseeQAs5nNgsWJHxakh6U6yMoI4BDr9Ory+hZzhnqAaoJDCB0GuA3HPRi4wKXw9TpzZbq3js5
tonjQtYAFeJbkJ0m1/8iEo3Bn19l1ukOd2naysj/Cvp33+4t3lzKAIJPU/PwAoWme4l9NHeiMb2m
ctN6sU0/eA1c4QFi4vbZykF9NpkaFjExLOWIWAPdhmsJSk9QzaABMdqEMp3r0thl5DLmJTKh5S43
0mHas+UV20+IhKmtVeNxCepD7QyqPOzmfp4uFtUkarch2Wps+QRiW5ikXMqJ0BMc2UrZv7EJcrvP
ukUGAeWdp/RuHgD5wcQHw1d7W6mo3zpjQC2OSRzq17PAtn9nI0vXyEZw0j+gaFCXPUUu7TOvbgRb
zO9mu0weWgc0K2tGTB8En1yute3eHBVqMVCuPkWb/WTIoueKpQVxAKA4te0XnccEpelyh6vSPgtj
NDBHWtlulPMIP7Q2us6XsgzqwfA2ci6Dh8Gpokb9Xvdo0HU6SqQfxYr79lsaMrUc4RNFYyRvJMAw
D2Q0gAr/jKXMdUXkbeqC8BTCXUSdatJ4fG/MY3YBMECLV0f3nT7/tGWibwMWXeokuLR4t11HcufN
MZfTFtY2QjqD/mj6HM2yWI5xKCJv3hfSAnlYSumVmoQVeL2rFcL3VBoziRoIvFtGDQNI8yMMdlSI
BN2KG8l39tODdugag/+fUgFeQu9YdteDmnv+yDCqr++Cet6FifljBd8oztk1s3sJWYIlgY7uDYQn
U9pxgXbX6B2Foq3OXFnfopAULiMnssdwye5JDawiBgj0lVUvJE62WapZ6V+1sFc1FBECP1FAYxj9
AtOzDHttELfMQ2fZn3bdC6+nnfeZ/pg8J4nHTiJTnAg9nfxzs7kFqhj8E9rnrHJFvT+SjLoo16t2
iufPs1aWF9sKnjxjHOHIbjDIapxJK/L+HimMrLCLAKOg0RyQXN6WgQNtKVJ0HzZNhjF6gi26RbmL
oTgLtndpizsIwlqtdzGNv5XXDjNwPUataAmfptOVR4pBdKkXfR7xvy0VxMMVcdPfq2Ug7ss6IWN3
NWcBIp9H+Ig+Qub2SPd5RxWSQrcjSJUEV+SrsOLdzCkSwPtHZplHx7YisXjb55z00Hr/nMYMug+i
aMEHkozodf1t/5ThYzKi6TM6U0/d5jtsQ+38dzR/bitWamI+8+BLTIJFg6eyNNhnyTi9uHxGvGFq
KdO/R8AR4SQeXw6StOEmsj71aNDPwjecqoSlR6pPe7mFas/L/A9E7VLxxuIJig3Ny8Rodnce7Fkj
yLnLoJSg3Ba07N/+LYx2R6+gBdFv0oMXwMyMyA09KS431opkcupJPdngrXsGTWPT0QuYWT2KzjKy
6BwewF/O6PlcwnY1zNtvUMlrqWGiWde69Tl7vdGdkM1312aCdKgAEyxdAHSMyqFZHuMF1ov20INj
ltlM4e3OQuFyDL7kX7exrXeL/UkAUbvQK1ngA6osndLBBuEO4nl4SK/2qeUyxq06hyYawR48s9y5
ihVWnGTbH5dCp0M7QR4dnBouiMpnetoJxK11JuyToN+wdNK7L84nW21RvGmzP+U5ofwho8VenBaC
wegrAC69+eVOe61NcsRmGvoYnD4xyTKYd+Tt4LxwqXrehNokWWgs8penPxkgWBlU/H7OMZjT8eev
yFo3UTghQKDdLGjCYMiLfv8iRBo5TQFwiezZfujZPNEVAwEFRbfIo6z2iZ4mUXuo8MMbo/QbRDtw
P5jUjf1JaXCdq+OkE0qI7ZRcu0p/WEwn4mSfQYYRurmJqB/dJkMpFLkmVv6ZzmqR9muTC2HR+Ct9
0MEgyP5gmty6JuVq9yqcbToJEUH9qDVLb89tYAnfIZ945CHfU26E6FZj/lUIiVi0iNuxJVEV5qpK
gAy5peDYnHRpmJsEbCWrNvpPKVyx7/vjRfLWTnv5Rui3C0ygGgq6OuV5bJINUUqg9W6GQttPonBN
eg5O2+mOZFz5NpFJ4ucVv/XoOTTbFY3fvLTYftdigqD4BHy4otalg0ljJDR0JwJ+UAb1vdHHSxrA
zsDzQa+aHIYzMFRKlj3c2QyTZB+L2pwpTlc/0VRTY9M0v1/ASmIbyr/9leNgke7B3L7fTTqIiMbY
j92vUNMo2btwRS5VrsNtnukPpbkOMlKv0D8FVDIrd1tCb+80nEoM5JO7HXm+woROtgN7ff27FKoA
dwn/sJsAQXEy3CrLZb9jT6Plfv9wWbIF/eJNMQOvgWe+a9unrgFcmhSMV8bDfeWg057wU7tBMOvL
lQ0hxZUO2mqwvsJ/W0tz09E+smhnljIBkOd57jMVlyHJYyaBsXaPS7J8IVzLjsVjXzY7BKtE7a7y
fm4Xu2zL0nlYFTyi+LdpLdFuizmK59dhMJWMaM55Wgt0DA5sFcxXfesps6KI+DgdhHogSZn7Hymn
Ti5ijTwLL3uCvhxAn5g6OSpawW5SBpnRBYriYcSPuCACAV8s9IIyrZ592mgVaUvW77sUFTPx/CJH
aHLKxHF4O+fRVfKxvzyfdrqwSZ4HUXLAiBYfdLY9fOrI1n/zP2jcxkk/da5k2y3jrUx3ahgP07wf
8P/yBydk4wLPdJuzbXy1HC1dnmTY0b/6BUM1GGFgalh67M6zuPp9ZNKPlwf9F9HaXfIcR64wRfNx
yexhWG+0383oDbIDC2GPTnfpOTENseNGu7UoJpT5Ab7S/8Re739YIoZHel+GMSjIah+rdcCuPs+m
MmUo2f22eqy2kxcq4ft7452QDlvJSnGDfYfuqmyBXg4/7YqnyyyO8xhTHKSFlG4bfYT6k2fB+ajA
FCKxtnB1TnscCdrn8M1VI7ytgVhCsLFKpzt6Ttv9V3g4KHPwd9ZMPveRUuV/5EJhRS6jXxsf4ZXt
kLcndsj5SPdIZETZzOktVrnZsuxl4dspox2vjzcDU4KZUkUNkSBm4fn3SQg0xkZ6njHmlpg/X5ce
2CQEImhK6B6RMj8fEyVfjZGMI1EszTBAJhs3XlGc822U22XxoM7m6h/P0ZoapbXALXLAuGk46drV
CpxorXddc0Sdmio0JWmH2mzvE0D+DnLd3HwVYdO331i3fEPfyrK0bcgRO7kkPy2ss8/ju/JcOH+l
LQY99fAynL1o8D/IfWM5tjZF9EaYfWNsQVQvQ3oTTX1cuY+jS+fO/vCjTXpuIT3HZKO5M6HwV7pw
tMqVhOEa8ZtzOb+V1sQHat3NSjc9AgdMDqhzmiaIejLujOwlCVT5uV6wJ+VjembmmY0KhqkuFQk8
p4/CH+W8CGFsL5gmUkEhVvUblX1SD/gbF2egiIcFynWqwVTckmbedCY7Pcm0NRLp2AWLCnB4Bksc
biJRQFODdo2sAVAqHoH7Sj/qy6tey/VL5OUO6P8ZLBKoAO70mI/1+Azo1OaT8683+xkXtvukBs5s
BP/qVpVEyliYt21gLlwoGmNYNUNQow6JbzdzbCnZwbvQKNPYLK1CuEyMqZ3rsSdM/oF0sIPKVya+
HmnYkOJPr/X23HZHWt8Ia7DGGU1AyMKOj25laOPkrL0lX82SEb0c7ouOxKrvu3L1wJw+MbL0uTqd
7BeKWTcvBw24LuSNzoWYXkE+Fx92tDic7vtJqBhhc55n0V8uPs1/fHTSRLNgLKCd25TWcil6+2fL
DP1P5qtcD+78aC6ENzMhg2Hoe2CX1hrf8UGAKuIa3csQeTaGAfyILdusmg7Nej39+NxvOsXwJfHO
pOonewmqbylEOK3+Q1re1LdTIFg9JaoR6Nf+RK04y01rt7NhO7nHtRJM2v3omHuhXYw97xJZ8AvF
L4VgGohwvvfKEMEFe1UYYWIDA+U31K/blwdUSPf2YEy8b24mi6P8nQeYAjzY7dRwKnOmFhiqHZCA
CxBpJJ6YZzGJ7/CLnGazm2ajvWCFU0uZp490N4dn9+IeVNNGIvfe6e63xJQEQBubnPZwpBbV6Qsb
PAnH3suJ7T7k6VD93qfVKoNe+eSIN716LhoGd1TANxay+Qg1qt6aUGpaCi472id7T6NIYe91Pu8q
52f1MjXZQDqL38gGtBLVndrtaZaiOkcQEb0cPoIttArblopYhuCKGhlbWaKsE61VeVKHJkGooYuQ
1meYwaTATt5D9YXU8Giuzep0ecj9TKRfAMuRg66aMO5UYQTslQd6L2lEX+sHQYxz16Rdyixcu+js
llYyuiteiNDiXdEID+CCRpHmcIdXJX1Y2gKUWPXMNfxjjzivCHW8EfNDAlIkx+BC78tFyJhy8wfF
dZNduumQc2J/sFMYwoxq0pnRBUbp6ktLmVlBHAK9O09eN37dAadsOz4xt9PONj79XNlOzBhdGrSz
J4n3S4GiTutIFtRS/gORChc8dWFQoi4USvcs95/xze0bbl5y6RcOlh2fzs4+NZyo37aYG3glot8X
tllf4NKo8gRSKZWsLQBuhde1iDbI88YM+utSJ9vAzbq2OKDngIruN/Ibg/4+jEGDYc+xe6q6bFgg
n6rNrKO/ZGjXjRZTDKy7C0rTbTZWmbYodwiINtvmxa5i0VgZxfhakFOS+phRWBtAHAMytJ0JW/mR
Og3wjfW/6x6rmijgNQvGTt//4hGDPTSKsnTCQNyxMTmZUVMlxm82HDpHf7C3btWqsndjriq79wT6
K3JFQ6wFwOd3hR8mDVzb9xCy9X82MWj1b33xjrs3snShMLWL1oPakrgalYbXMnYdLtrAV/+nTrum
hUdHHPgC9ZaYlK32zchYRSspmBz2lchTJDbwgkteThCgzwndRc9TkilE7m4F67QAnbRycuCFZupD
YhTiIS9eX38TCyeAEOoPQsPOFJf8Edgk1x0XE2sMJmJIb7oMnmK8eX2e8Cnuz0gPEbHZ6gnbQhKL
ShFv+r6/mmOh4S31WL2qqOSmtKZxS3BQI33kwyXvGQCDgKGXAlhYBBGWuZNcYwq2eqqhJuAkNsWE
snVpBqSpgiAIqHD9oZiM/pQVq+PMw2n+KAHwEjmk0kT7Znm9+85iEJ+hRTGIflRFKd3zumu53E/+
vvf7k19xSGY1XNh+iTe1nAej7wXdcciuqn+EQT0gF3am415iSNL3LWMy+Nh0tN7I+8LlxJ61v+sb
TKkDMKghVELOIsUj8tOFQGfc3J29AX0soE0PnOI+Nx6mmmzOVHa1ij3W7SbwoHlbPofv/mzTMagH
mLmkXc5FtSVCFhhh9qHlS1K0BMArU3H4Mg9NV1ucVRru9dBDAhi+SZGhgb98ja3W/TCbjYKYUb9s
txWSQyXKD55f57vHR0gDdAlE7SucVPKAPPmn3F5IrOsgAhqWdJoMLnPizLKj5ootRUVH7MYxFdzc
78duQOBQMO9PZfOB/+vfRcvlt++6OXMx9wJ92vPAtw3bHEhH7dFYF1j5BB5dRpzNPbZXb0DW1PV7
acZAvuoxf7V9BP8A23oj2QGeyBtkc/sXFftEhwucvE56ZX3/oMzhV/7fTTfNQJHkatiFf9Uhgi9Q
JwsL/rujVSnPn12BqJoeEEPc08FNKA5DXzaZ9Z6IIyhH0vHJ86MlTy07CadM3TXHNIIIppr0xCNk
60entGEZ1m2zNK7sxMM0DMcYTFC3Ve0t1H3DGuxCf8ZMeGMROl1bEdw/8nLlRSNiTnmHBbqPZ/YP
lIUXZ8DzzjcRnRd3BFXDlU/Q6Bz9FzAlctJI74SdtmJVh7uPFPSO6gslecHdYDLmRlyft1RxUavT
66D5ckcCxW08SJ1FboZnrYuj+nwVJSfE8YHzKXeeKb4a8QcRopJ4oIl7MAs1HRYLXfNx1MIuPVV/
Vdizz5qMIqrZk1lIok9/gM1pZwZOYqSalsqLME88KwDAuwc7C/CfAn4XbrecEIlCOBTcZYWXZIM9
qhjzbocxckahc/z3s0ua2wgotbwGduYaVuUm+8vhlNNLNxqJcVpykOqbB3Dw9tXi1qmk4bU08Jqv
cGWPLRzdDYVESfy9IEXiH1uykPoW8e7ZZH9HWcvnJNOKjGuI17kKiSDjAw9FFKAo+jKPVehtszJB
l3Y4kU3Qr0qEmtZDII93CAfnU/p3aH3vgtGVHuaoP+j+SDxbFCr1M3SL/WtxnHenRqvDncYo9uy6
vPtHJ/7sXuxzKp1Sgll7NaYzyO71+YHKQiOYzo01FiIN+1UZiuAZXOGUZRog1neGQFLMydFCI7Li
rar71ztoUDvfAxnCw7zSkpZjhkcWHepOoXbsOPLPQvhpbo3fnAAh+pYz33VTKlr1JepbBtwerzTy
0/ouC8ol3YrEdPYfZN/kWee8ty21CUIXuWlHcHc1ypcj4/XbrZMk3pwQv07DdV/BROsqMA5i822H
uBbxxAu/PAAVHzfWRwCWhvRj4sWRjmiSY0ygmK6sQz0qf2AdC0ZnPDKX5NyWUVW9MbJka7dlLSZv
zB0ZYJqpjXC3S2k+MDqR7XbCou3S98eJ0AuGe4MU0w3Jl11QnGmNtmCq/jyzU8XT4a6PH9+6tmot
8znn55dnq137u7LPOfxQmh+QSjxCT4jTfVg4iMP/9MmM8ndQ7X/9a8RGBAXKaztuJvH+labRrFkI
GIipw7/pE5KMwpm5tDYmj+J/3ob3P7rYmMPnL2UyRMiF1tL967F0NGioCKWH/I62ZtUNtUVR3/2u
XPDCIEqnzmw1GLM2OVgnYlTJKoRTP1VoF1LdbrPpr5jRYnlvXW9/Kg2HlYJCjLce4Yx0Li9MrkM8
qxr8u5QhbaTzknMIOq28FJb0f2gsxPJWrrK6zRfLoSfpxz0PFOBuqqtqrSxRGi7pwKuZ4M6r/uhF
7tvvH7w7CQEuvk3viE7UTM+vKWDC9sXTGgWiu2BtLi4g6SNvkf9njZqPVWtOHZHEyRlP522mDLRp
RjkAD78sLyMmddtgA5NNTF3c9+tCyRS9yZ7gzrzuUap2+O0tqk53hUER4IqaDjX++3Ygi3ViTgY4
N/HlGjuudwVyR52MSqoq/VBppZhnk94LtePLM2AFS6yWe98dJQJpJNRVrtNWCFynz1V1o2o6Cu+K
SZx1ZTr9PSN7oVHjEJjCtWSgrXlE+OHC7OR4uKMIJAw/SxsTV6li3KZ6+aCUhmDvYHZMjS+FxHqX
8FbZAgKyLuf50pfl/kJgO3t6QHPz8K2lX2HL2GnLSNkkpm/czY9Wt/4Z1MYOvCetWlVeuIUnRmxs
o6Cu8xXjK4NqxM9YfCnfhk1I+kLRe4P/dNfhj/RtSRpwqwfr606GHPt51+qlH2NkoLkOrBlHEav9
3YO4ZZUWX72Sfbp0B+p7BKmvbQq6UaQ5b5O450VUNPC4nVc+GLuBomfKInA9MNyZb218mYDfGsl8
wb2Ra+25DI3znN7IGpA3DdSzk/14Pfh91xwI9qvf8r2RODBlxCuzGl6rfbSwPd6tFqg4Nw5XstVC
oeWMYXjcIMt9Ca4n7iKTiWFE73TLFMX2oh30gIm5jpbZgVu6jI3SVm+op+WL1Y+55RMJX4sW02Zp
dWvg1ok61OcG9BFB41RgKdy2j0IyH2DWlrTKQN+NwsWCaecsHg9rGOx5L3hJ0Y9+VxMrNUIp1bo4
Vt0oxdg5M/NA8Kr6UHkR2oT5i5xhpx4AvbObYxGWPNW+WKZmdjPKSkxlDH98UBvGqXX9ZZ7CKzzn
yVuUB2fU4q1pylL5NxFvcbFbQSp558s6jYK8vLM23iRXJ6a1mnDsNVTi8jTp7NkW2fkavL5EfqWC
xZKkXtM3sLHkdiDvUSMjvFCsCLTtUAxraMUuo1ekD1FvSTrIHTGPAkUsqnsD8vGm8LtezRVgSGti
Vfo/mbLNHbdxRjT/dN31qH/FejbvLLoPwIJIItnX50NUQYzE50G6Ae8VrbELRC4Hc+okBUNix18E
ouNrt5hiA+vkJXlpgONtafbUUvK30DPHN+E2Z5mwCD52UE0pXwmbpQUqUaGYO/iDauf3og6Uc8V0
uZBsEvocEQf3dqNyf9vhxt8vH8XLF0WFw9XaYYb5qc7e7VXUaZtgPJNWkBBDk3+iF8AGkW8UQKny
gRM30nnoZf6sChT27BOL0LA5Kzm3uW7DYiBvb6j/ClIuD0hgtOTa28TxSWnSy4exRZxes9NUJdCc
LvfgVR8wYqo3wNSEr0DG7abX5owvxqAT1ArlSXtSrz3H6cBMwIn234PNK8KYDd5xj0tHEKmEMETu
xEP5TETJlSDsvl4DIClB4HffRNJxPaVtZr6uQWB5pyXOVWcxXjX+3IfDndmXU/eB0n/nMxbo34vD
cAsiBOOhTYkgpvfSDa+oJLYIqeHhkTdMwdcEcUID4veJBIvclnopTfZSfQ0ksJkR8/pslIEDAPqg
nR9q3DLvhOeV2aeGMqdbJGCDnYcLDsOWx2g6UBsQJMcs6/Z2IblccbGHXJdHFRMf+w4JmfIrvLJL
sdLzm18npKdcdvf2ewJUVK8ESs0ttzL+i8IksRa8950Juy3fiy5oGUCuXFKt25Job5cfdrW+WJLt
sRCT0LZgZN4IGEXovbYDFwu/K2VypqbPi8z11TjL7+1n9qO4xoJoEWrBoLoRn7fvXQfygjMeM49E
e+3ua3ykHrDbMYobC5UPhwg1jvhgSBb2TWmmRWo9IeSIkX6Dn+GyNOOHanFcmQp4b/Io6rz5lCdu
DN2KpH59aQ3kPtu9ts5MbfS4sdmZu1bLyuUghdP8OUlIPMAmtIYwfR3gS8QwCFqCbEpmR3tPTSK7
FISfvijvSTTxF/8bexrKLnQdj9rwjatpVEVg/gxjBr2Oy7khcwVhVSNEzqJap7obCtCb/7UtPkqe
G1ECizPcC2rLl/2LjnwVb1T+y7C7xt+EOXydNTxuHILgk+o7gvMlCs6lTkOKSASf6eZxvvxrvkih
aA3iSdoYk9iqUjcLSLbZadlztkvUzfChKZfQpnqVjlvYXV4rem5NCGUtq51QEsFOefFH6QZq2f1i
QLYKMGDSypMvCOQGZOlAQOFORqVg2UzpEmxF6WebxUjz0xHX7saj1U4thvk2Cjj6tXlKwcj4aviD
q9T7uLwFaNF5eqh8rMSfxHNYiDsKiYO3wEmda+jIlqAWT9TuNPfkcXY7L2qbg+bpruA5HptaReJR
gXhKaLjX+5IQQMSTSIamnqfYQfyh5KNGQFNBd40+UGzNwb0doeZl5lQcwMuMxPaNMqhqpkXDnzhy
ETgIS/P+CqsU8k/GqrK8i+tGMmDgLaqKv1AABvbDNuX1jvdGOnM9FkuDUs+o8YLZDNN56chX9FcX
ZTO9KRMMXLmGXKnhE5B6Km+R4RR/ZONcyo7e0T5sy8RD4iEcx2n5N1QR3tmkEbVeXnxmesiyq1ta
+PpAWnZKn8i6Qd8pxpkLjVHbSt98o2VmgU81LEqDovOihynyffXe58aGgd5Ei01tCIk6Nw2WMSYL
p6KoLRXOzZ2eEJ2GYOuT1huCE2Dbu6hiScCxkrba67pYKYlIAqYKrHcgomxt6/BL5qnyvlLhj8Ko
/bcHwzrwEOrseSHitgr/3ycK/o3ONNey/tErVS/x04IrXSPNvVNRf76pJm/iCtqgiiKl4fkKHZ81
tWWJIN5HCooInhBWBzKe3ACgtk3XperKF4/PxTYNieeFhi01fv8pJYkWtGofDvyHk060X+/M5wJp
Oq5pt7OmL/9yrYaZnjuu85vFqqwI63bE1HsJOGfH8PP4+tkr3urWfrD4uxoS5t7cdLw7Z+jq+/I5
Id6D8hHzcBrfwO7EXBMG5W5suSJ6WfOMBMkJlHTV5UNH7Ntnku2rqiwrJdwHdSyneWl1V25sHMoq
4FNWHuiEeGo5crO6Rw85tTpW6KP2bZcM4n4M/GOKhXP7i+jm9kCsSvtqLCG8HY49F2T/xnKAOo5D
+ZpKMmChQuptXjOVKG2/u3FL0Km4+0ExV2uWePe7T4A3ipX3413qIaJUX5khW+18DD3eoh+4Mal4
9mr6EwViPszLCFUItaf+JWMyrSNUCxbgykiAhutflbXEprqmsvOPKZDVvSYXWW8tNgeR1Ewnig+X
HrFmRI6T/MqpJ0G+UVAPdmczUW57OKdaxc/DlKONF+uPHBV3pAeNGFBXyHexLDx2GmRRUFVWjdr/
hMWie5PW6wceG3u09nuo4WuCPW0mGnNMP49a1YtGVpqwcaGY8HOH1CNRS/fbShpcrBbogHQvF4yF
pghqlVUi3cvJ+iHNYOi5cLdz16V0RD3w7amiR14LG8l+8xnYCCgGeFs/H9X2ZfCeS2/aFfJ09CbY
Mkeic8QoSgVAsIzJ2UWj5BOke6XDN35vjhSSmSo3YchEJnpMPytA/RdAFHofGxG86cI5S4ktFAzw
rsUw9Xf/hJOxFF3WSEUJNXanVA1vK1TPAnLQijIUjXYB2hcxXTIo41eOVsvtErAeaVateWxWAQX2
Q6vBQnOKnEgu5xn37lcn75pk0U9rC1BtaJSbVCvBiCFL7itBi6TxKI7mk+G1s4LxD1J9oB4MqNvk
g+n8LB0TzVzWaI5Pn6U3JBvxT3fwpKqE2V1QhdyO7J3Xg/VLzFmdndrbK01iVcKk68Pwgxv2aQft
ZgkPU8jdJ6Q7IFTYcrMquNgOjFQaAm8vDHOD3HJvVT2nmdzgPZcbdBYAuEx+lebx9CUwQkPSwxOi
E8wKIAPW6RHQpYYdI1ReXZMNeeeOCTPLK4KySHC3RnZjv0izWS1h9Y8tKWRlKwdh661PG/lMZxdZ
IvJPZkJgf5SMZP2qK2RvFzVEp6Z33hG6fdm2Zq89mRPaau9IsyXfq2VBhrATPnR9FEDPW/JjXf/G
lT+BPa3w3wyPuGbpzMEt+A+jAHMToirVq/aL9r9nip8LyjSggvg09KJEwLcW9eKs6jWjPAJIJ7o7
uyF0gi2fwgK6fsNxIdgJfCXj4noVOeZSjVK9PK/nvrlMrmm+clkgeP0kTegjrNB68X8rYmdglzCA
tkTwYDp5abDAVMbqeUypzHKuVk/yhS8T1WspJ1bwhM69DP+ya/5dC07ZSKCxWwal3JijByoPedTp
qnC8C/2XXMphBbAdIRc0/bqF7y48v7PK0xo+dOaqK0JfHXkFR600aCWGIADzVU07iL9lx+W2Q/Ou
18cc7+d4ZrqaMd/9ADQiz4fEBiG795fe38X/FAljeJabsG9YyMNl4mWJ0AmFMa1zDZmGUVJBROfs
0enFWX0nYBQnjJOmMbUT7feVKd9VRwv1Irjltlz8QRnLy9Io1+YiQs0XD2fmqtrmlvUFBSMOUn7e
Bzi8SBE/z3FJXXz/ba/6069x33xmTG9bOpSsx3ydpGFWvEV+yGMAmMVJG7IOEb+W4Ywgk+v37T0I
b2/VtL1+CEzQbuYVrVBZhgvmdED2ZvMfErdIoqY1lShPCdha2d4FHkf9FBEFKPfa5N6hXBN5qg2r
/PjXTbnU/+OGJQZv80KTy7900GuSkt9Y3HU9Rbas1ucM2CN/9fOlGkW+7WUqHaVFm8CSk5+ivxPL
XatCr7givAK6ZrMU8/E+2dnuoLWO0Ox3wi+ZXlSxYBqtilt4fw6ZTBBiYL3NqooDVCBeWOKO4KRv
fcDzuEorIHK7MrMRt6wpOYhZnEuilW07znExmPlbmtvqgwPDvtuYym8Z81ikiazOv2mu0goCOjqo
yvCNeruA6mDhUIcrwU0hK8BpCBgxD8IqSW6yQCOHB0S+nVBJ2Lk8QRZ8Brn/FlQbkwXxua2iHmwg
E5xF1WPJSItLQzkzJl+DaG+FR4GBsAlOxPoOgnQdWrDg8cfdlG1Qm4HG66wVuszxvraYjDFlxJSE
2GTmK4s9kikxFCROqozzOGcpI6dkY28Nmg7JpS3NXhI6WUSxWr287oPEL3HgVqnE2NZgZNpjUPc+
j1oWwQNd3GkR2oqLgLQbfs03D7O/Dfnc4+i8Qmbp3499Bp0HG18ONlk+PCaZeUXgqouL2oVa2DDU
hXhtiOsAYLRrREP9dT0cZ4Sy4yDp+1BT6CPmVSJ6pXuelz4icmN2AjK46S18qeljxj+D7IJt8jsJ
lpanqQZtbojwBjjgUsH4No9BCsipveP6iTVH0kzAtkhG8a7fOKcTBZ2U9K60A1YwsiOkDt3ofAkZ
DD6kGnv8pLX8GfV1UARyzFlEs9L2K3sMIg0N7cZr59gB+h9Hd9bLGQ9iJZhaSZNVbGPgGCiAj9+M
IrgfrhskNxqiP9JPECx6rqw2YSOeXKf9zxHhH4YsCJNszhXudd8kR6LuBEfeB16uf3IJJa58Pzwl
6Y4f4poATMsucFz79GVb5uYONCO8zasJ4eEzdy73b0V0FSGihAi5fJujSHcVRzWpQ/6NVaAkGY2+
4Mov1Wtnc6FDirUoZMgXm2wh8rsAn/9zamqY6iVWnUniNYuubMf2wf0fmVCyBRCQ31bmGc8CjdJH
P8j9wOKDnSh+UWTGUdG5ooxfXfWuCGgnj5Gvv0RjXTKHOqmQbqSeKZ5hKPnFIKcfF1se06GEvNsm
PZTVlpKE22J4CYU8QPbXOrJ9D0YGHoTznWP1np2ViWm1pCS1O8ynKyYqxc5wZWshoauWa05GhbW8
tmnzR8HQvXnBfe5Ej69VSW7sj6z/stde/HgdlJWfylDyPCwr7QG2iKxqK+cEkhdpuKeB10zxMbtO
33MX6S+N8H+yuRm43A8v1pxxERg0M+ph+j2ZHAjaYdZcT9J34RxkdZNj/Ng9dEFYVxtLB4C0llly
VojIXBc53XuLdsp8mkG7IY9+LeJebw8w9Bwdu6F70yN5HRci1ngINLCofdB+s6v9/yr80dv2CuhI
O/tdL03wkWGuJNbdO1tomoGL91Zu7eqT00p5MGs2Pf4yvCXhqNcVxIrlm9oS+7ZZLW2GtDF4UqFx
VhStJpuBZ6IrOyrir26Y51dnZVayTTWD0Dy0LHuf3Dzd1LYgps78mLYzEj+BXJhPBi801gQk88k4
0q3e8LkKQR389o/l8ZjkOkDm/P04VHCVxzPKfSPB+0/nvql8WECMPinVUMDDBf/7mlp0ivCcqbw/
rw6cTvCYPpGfomiWD9JDSWnRtPCS6wjh9D+M1RqX8skeaKFpKchdq5Acn38WKSoE+0nXr/5QldaT
dSdYDKo+8TLRW+2mPxIR1lP7SnTB6HE41DD+MZ1SoinlvdVgS3XrNciCdUKMQA5GzSRxS3sukdl5
A18PeaKyUNqOVNc2AoNJNUn4WBWKzuo/d3oMxIup4wObhYpbsvsWfkeZ1+aXefr0nd0NCKBXg91w
5zWsvQ6jpLCL8ReanKR4M/oT1tvCJ8wO8PzoEt0mzb2dBWCEbtLG7NUjySI5UzsPP0W2ZHOay006
c3EknbpjhPhlq2h9kJ/u46by7NEeGqLLDI2nS5i0IcXWCD6H+rhEtkETt1PBOX9gxi+p5fl3/tXn
jKG66ClglqHWfouEK6zpQXvRwmoiAA2WWEa2cauvBZem/448RYRqfX5wpiKiX6brtZuwZL3yPQGn
eKiuBvaMcyaIeFy3WQe+wXBcb1fZ4AQ5SmKqcquzTBW2PpfW12xny1sxJxGNvXUX78GE1uIe0/Eb
uzGkcMCV+wLe5nczbCopR1Zvn1dvHPfTo1pwuPoWe2I7tsEi1/W4WsNdDwllLA1Xy63p6wOmidzJ
1up6wCEhumRQampKmJtHSOUDLcH3pld5w9C//FrwqiKMEeTtUbLj422EUU8FezOtXHT3Nlyxfub+
Ct+NDQSHgo6x73oPiKMldbMY1gaiHvvzo6uGjWfhFZRWveLH8qPZNmd/k++JHHJCv45V3LrqXhoY
YdrWsZECW86hMQSZoEhh/uz+PfpRxQ21bgwghAENBdO9hXFV1U3TldGH/GJXzoA4J3q4IqUZsZPV
E83nfNxvu8nOxjbvkGg8hi+4meEPWsUybOx84HQeRGG/md49GBheoeJi/0rPlh2TOz333Og7SxhG
xEkGRwYrw136UJrhLPijLVsZKzz49o2pCQS9kM9cxaDeNIo6DZqsBlfGBshhUOv0RlCmIzekDkrS
4tJYxnSBIJAdPpCXQYyoEXFlZFW2fRf88I1jfszVY+ZodL/KuEOwZm7+QPc/m3h7gOVTg8774iJB
h6Zd29JqlJdvwEp97d1z8VMJ9pi6TGvyZtgf5TRraml0TtVq5awEnAkt5JInmOFjeQNNlFh5WK8u
Bwg1W/RcuXVIS7byZ6nUA1QHF2KDotToUlKavZGT0OUQvsgZVxIjZ+XfHxf54guL03LZH9t8WfGD
/yBd0t0HqEc7duUXK5ws75y+NxECu6RKZgJnbbBvQwvbNmRZV1MzzITu6KBo1SLsRfVjmT4v4PI/
C8D7gsvcazthxHnFs7uf1mEucyQEWCkoZNPAnaKVTNKXPcOa+3bWY6KMfefc7G4eLr74npqvvuEQ
vSpkxYkkTkDmIPnZxkOBiMp2HfwoMRMmPVioBFLtCiVaT66HLV43zsJ/rHCJsWDicuZkS871PiWc
+KTqZB3CO5aVMA+EEDycIW1BJjyN1AbZHonzL+84lNBk6WtUbgREcy3FS9Ee5OzCoeg4kHjq2Ikw
/vWcrsGrjT/x6k9nDj9vqRnfbfiisB6g0IxLTC7ErFM9cKetaw/9hKCViGSxyjJz+EX8Mj/Y/grX
F6ihKNAaF6zMyjKMfdl6gi64BoVSrX8FgvhWBOYc6cFHU/OJT1ZTAKIZYPoACyQOKtX3jY40UEPl
ci1PBUmwCpuAnhadUVIpeuSphCqgRiCyH5U5O+AmORg/Q4PLRMavsT5RSgxJxaNlFaqDohAyY1JM
Q+M752W9tcqaVuO4Ab5ezsZi4fBmF/M0S2xAAKmofsGwBjClKzBdjrkhX+nh/rYB7mY6GPmzMR9o
NyjLMIjf115HXfuVy8C22RVNqPBKLHZP6JTahTFx8+6jLuRX0R9ZHtH9XOjQjFNiaFnQcbVaLup4
Bub50DNKKpK6xnVo2Q0DO+FlKxxdgZpdMCDD5t/3mopDogSO0u2An6hadcwZHHmGzgFbUy/iOxoe
n3/cpVk5+0/HNGTZiPbPdTiZ71SGV9a91X+eFc4mnylrmGysZLvnAKk/pidq43DVgYlbS3Sl02ca
kdHhS3PDqhiiNyKXli/zU4kVukvgMv9hf2Ny7feP2FqGGt28CztRAU2hx9v5iCPNBrM8v8pYN8Jg
mQo2GrhdtRZFbA1u8531Pyz9VMkTwz4NsV75alhFHlt3n0UxD+ndl7LBkO2l4J79LRIc6Wf7hclH
0Xnayb6/lwTwZK66lpPxvCp1ZEeeRqzYSCELwJiDZMjg7cujk2KPBMDXleDGchBMMUoGahbson2D
JJfZlVYHtPY2VGX4NiJbqhUXji1fH84vQmBl07WXq4FQralWM9lJx/j0xxeHWgYcUPK7f67zE7sw
BzWrarFFO66gUxQ/ZhG6NcOcVGAlP0ubTRC3RSXpQPliWL0ObT98G6XJ8c+/FtgEx1dla/vwViW6
/cM3FSD0Ge0se69gw9aWOemrang7kTUX0sdeDYezolRa2TYdSo88O/sa0xiHGAXVfTIj6kt1sqPa
nQ2ixXgK5muRAiia0b7UAenVqC46wBvp9U6XkHlmUvncmfC541OZwL2j9FrscOkgCaSg/OPpv4r8
T69/+DLREkzpggZpgoq7eiYS7dvj8Qf9B5cIntRWCX8o5wrpWMYejkZiFQ+kBWRMpkDqmb1xqeS7
mDuWKQBrwVt+VeqyTqwd8WV6eqOlt+910FaaJrsJSvwnYdUjEDggfR/hCQFwTylgSDzVXJ/AB73d
UhEhvfhmTJabsjley6Xbqo1Hh91hX1idankEDX+Lj7oj9G6uBjMTN2RkYhhVZSHaa2EfLiVVntnn
OT0m9HfQKPKdYVST+MMCC5W0718obxw8PE9kiPGbUUrC0wQjE0DT5H0ZnGdOU71sBSjvCgeOFIJ4
de2MlXuV3X8iH2sTKNLza8imtrid3cDM0NyDTgOpxkmGnhGmZyGQkd+1bOFzjfKqGgFfcU75S8SL
UHb2KYhlQLpkonR3NLW8gcaaGJXtIYluDFA/ocvX1fLsy0i5RYwN1ldjXUbzSYiF90FPPSMOYgkc
ES5NqE6c47DM6Rj5QHBsqQSnmFKTbaTzaygK5vPVBJ0omkqYm7tyWF9YDgHqllC5XLLhwTF5UezS
3N7O17ab3/qUOmfTi+4wVJLBBqNfiMWf6G7tpS84NngctPM0EvcfjMNdWGvZDzVeqmfUiuhlq9II
XEoNEDa0BMczPCmQQWQC43vgYveMVvsXO9LIN4ca5xlZvAREA5i0pvmoyGKIkekzu4U2DjfRfK7G
zx5q+QhzyvLZQpqNl4xrnOR7uw4yTE7KlM1NBP5y55MkYsrjFBqc6cRBMMIlD6VEN8EVA5ePIQLV
NNpbkxd9gPbmBvHyHIhf4x2ClE5XtKKRfbDFdHu8DtHVuwixh6yLdUeob03DSvokcwBRlchXCWEU
cnSN2ot1+eHSxSrYgy2ffPzgRzgcqeDQdOAJFEKqzk+77+RHEiA3pzJ9GY7KKXIiSi0OuvFsvMzc
gF4DBtg+jPqZM/pW6lZDI2oq3GHGpPQ1s/aUTBC2liMvKfbS+OL8OT1yWug5JN/S1u5N0Y9pdDGy
2BF0oUq0PLDJytKiMjmpNOlFyNJnVl07ab96JNL1usuXvOS//iIE1mkSIxH44vg0pRuP5xYI4zaB
MUbQTGLrErRqBOiv7CAP1Qf8uFWY9uvKhvmb1megVQSnPA9xWexvAKAKZSPrlpn9xYlAPXx8/13h
OT+TUh1ul1VryUIKO3nrHynG/capgOFrYJOt7b0eM505WFbDsVIVN7lIlXp7SrH3yfFyHAZYPzGt
oX5ql+TMGOndNfKXSkv+J/YzF55OabsMxXpa7wq+fY+L/Ju4r70BhZybgCEUOaE9eINkCFYRsBiE
vHtbAx+1ps2MAb/FPRDQ4b7qIsXNx6SqEv96EEbZZuxUWGxSMRIcU7Fy4hIL1SpZ27dspQxI9cFc
E9U0BXrVSukrSd+eBsxU1Lv+gFRXmMVHYJhB6r7gjBJMwhXCE0j6Pl8+/R3MxFiq4V3QpiZ17V8r
hHEybtXywWCyIIcrBdFbs65SdleIB+GbHVd7cwrK3UUu/LxSH+pFQv3aYBJhox62GysnszDKVJdh
0Hc0wyLv1A0LV4Vg8Ngim6EBhciVFW5a0tUpOzTUkowNDHaxSt6y7MEB+qrpR/n8+4KLH9Lzqh6l
ISoqZDhHa5RROewhijwwFTwBkYOd//sctTI11Sb085ur9j3uekcaPqmSoLExkeAKf4spdmcvyUWA
2LD7QVHAL8lBl23fA6YHt8ZdonDwVxZq8TeT5axW5SBWx5kKfzKw/+qOJVDssSiJ8sYyFshA6L4e
r3ZBIo4Xwy5pb/Ub+20vcKMElpI5EWtxcmf+LmwaiDaOXOlW393Z/PhVSzhURMwdJj0zxafZmv0K
OZggVe3SwA3eOR0rG73fsj3aEvM0n+hnI2Ib434LqGzUysHv76FXaj1bVGJI7El0jun8tyncUtxH
VZPmNw/WxNxW2q04TY5r4+z/QQCmtk/rZa219sZsRbAVsd2O0krmYKcOOK5VQAG7+Miae+CLM5uo
HB1frEGAkkG+GsogMLdIxxl3iDhFDGjSzX46eMOdhcrRNmLIf3KCh5JOI55Ab0De/vqPfEeFbO84
mhFUvoeX1HqNsJ3kiDMai3e8+921Em653H+5TNZ/PxuMnXYTdbL8G0zW1KSr75I0Mj/Wq7uuV+6+
936j3LeVk2FZq2WQOuvxcRbuHLUl0l3fpt7D5OyEa3ifC4aChTTMnUGPVdNOgpCvRHJMYDFYT/QT
y9s+BBcxPi8tfzscerSgsQZFgpGnmqPDbX0Rfv44T7LqolFj5Mqc/rjdMJBiSmz3t5g0TMP2sSki
HWS6zr16otCKSGYH6W2KEkwXzUdcIJjM9j7sVVK1BI/n6N51WWNILcYDDhTkBejZACKkMgsXlNPz
o6TxHYWnHo54jzXPxvCTqJmDjluvz/ev7b0YZEvovkbDhGJ3FrI253kp4+xN8UAK2I9pFHUkSS3S
3RFnVakvcafA+idytgbM2EtyPM2TJjA5vmGrMPG6pQeNUyVCBebqARGPfVbWod7OrnJz58iAINtR
hxJZIiY/5yHyJE+yCak7U7ADcoCBWIk+49WYlNGLtR45IoYgXlE9fVdDELfDpCONkpU17hs0H6bQ
dv7+Sk1NnmFU8k50bImIpgGjeWN+p+si+LdlN0HOfJrPbLgvBq4BO8aKxtzNKKryWyJeaVR3GZj5
otmqRci3GsFcPwav9NznGHj4059dcAhY6wT/glCovUDzt3WE3RHh4PzIYQYpSVWVmymO9S9BI61c
gZQjmgnIS1cgVfN9kvUyKrtA/rCGzJgqpGCgT7vJifEpGgr76lxuwmpOeFbM+f/3Eq6aDV4GFrHg
D/LbK+N0Qt+HCnOFrCxGWDRosFDTySkiU4Q9h4SgUi0BcLrat7p0t0N+/AHAlDY/l/vsad8jcKQD
PgzUHRSGQGKHKWYU/atrOTJF5h8KPC7kNGSAXIQTtxzfo9jquUVOENQ95tf5lGcBSUqS0qr0Q4tT
pCcLWMyK9AMnaY1jJhv+UAQjDki28Yhk+Ej61FrIzTQLiWdOdG2mi0+YUHdmWfZXtwEcW8OZ63x6
itI4AiihJa6/3VqO7dBdigthCLng9j5J2tBxRKkGVXLgDsnU7tll5UuSP+d6QDLLcHuypI1Nm2ei
B6eH+GVyrkyAKxEJzmOuxLoGrgR8J1swzaYqodU9mzc3ntJ32gZ/cyZhnVqdlU+JTu5D1uf7zGW/
7hZ8bjgJk1T6+Z9AiTtKZAZkIXogpy8MI8n0uZLpvcWe3SHI1Kv+FqKPU7zE5DPkOEfp/TTEhOpG
V7Dl3Y256TRPzRgjj4Zwzg7EIPAKEGsLi6Eb/C+Y0O6y3gl5c+JFa7CyPH6ctOkO6zDQ6HuON6JJ
UqAA9jqUKAlhN9rtDKNpS+3c3Zt9QvoXXllQZO1bv/tZWnf4s0TDOAEjiwURjgTVo8bd4FsX+FdX
GdZd1f9Riuz8HRPGkVP3TJP8Vl/ZSMRIW2adfUw0vh5G4/F5Hw6dAPrxYCs3vlzPOfu0nfard0nG
m8Yol8hqJTgKif3zEiPZ2/B79xFVHWQuE5E7g6wj9pUGpqilMcepH+A/cjwj19KMc/clE5Y8M1JO
7XLfCp+2OAUVhxxkZxMrC9rcvd/oidJZqlhrWVIn7WPGkwTc70/qgXYgC6m5e5iVOZ+ZctcSA2jh
lUY4R9SxfKH31/l49jFBSYj9M6lrej0QUsTzL85smzuld1ouQJdxmAgz0W5kB2YZZjcD7KYoikJV
Q+w59PxD1AeXsDdmKfrAI4WxIgb9Xh0SqPnVZ4hbJCZcgYofI7evWn/UqYm/0UaF32Ih/saWwVeD
BJPea0gqpPs1gGAvmMx7nrUwrvmPgWbaSAqikPiXizudG6HfdVJ5TT7vtgNplWGGdF4VLs7CbVF/
cPkvT65NdfYqCkkgcJbxL7NDb7wfOiKMqpj2YKYSsm0LQPounVi+SqfBk9BP3S8w7dx9/lEZKuYu
j4yN3gusdDFdpCDYAxo3MUcXfaExji+ZZnLWirZK9TgJ8Nm6DNODfDfJEEC8VpkOID2tnWUPr7Ar
K9/HBThbSl78inhtxcSFbAU6iTDa8Bva/Q8YlX40rcBXXwsnDbxuRFGWqFkLbsp8kXnbwsBXiuDR
erRDVRxiuHDqUMgZwji8MDWj/DzEQzSle3ournwgfvxSqRG7BLege+/wXqGLjvNOS8/8YxdXAq6X
/4QXWMraM/iom6B8s481VUaPnczWSrV568rg/0gH2XwKG6rlT5wvn2fP+wk8c+gx5JPVHQPnsVxf
HGL2q8Aq0FwsEIlEqRNrPYCQsFuvN3uN+276FFXbkWzq2mivb2eHJZh0/QHB4P4GFtrOf98mtJZi
hxbnHBBf1yIfQIwAh/4y9qgsvKutgUyjpikGYoiQO33xBPG4FW0o5wnZWvVOI9kI6Vsd4/sx/+KK
Wgj/HO5K6I9aX6n5SXr3qfbbK2wxj+HJowePwoS9WcFRcmkQfiu3iA+1ykUJkAjYvpTK/k3caD4J
bPsArJGS7QIYYqXUWyPwFhMBXgbnUNEsqJgRAgWTzDM5EnJwHsk0wOkRHxTjZPRpwbWVYo4BwznH
b64WnODxwO3ZdBckeWKxVyTF1ELWMOLMRhMIBhqSN99DJxO8S0M+ZTwTxhYQuHCThAyi18JGaUdQ
tVUIT2TeCMUWtaDgvHOh/iKLlpzcn/v9ZJkQPCfWlkDk75YqFojYTol9iHiUZhLu9rY6bzmAdgCb
X4MXt2x+w6i/YK+8nCycg0RWAv1aV9ecM00aDxbgNBCBzeb8WKvRYZ9b7cBuuf0me+cpKtnT8hU7
5Xho9uiGtw0Uw7sHtqI4BiJ7HZSqn9sJX1YNBSnKpCx63MUifpmMw60ODPlCftTS2JEesxDo5MIc
yNnLcg3PLY3rHsd02bpaOc8uYXfuw/nuvk2wIt7Rs5sk7lZU/XGKBqjEWzJoOQExT3nh0lYZmg+y
tb04y8ZJ1cG2bM08VIOPVSvBKOV/Mt8LZHasndJu1QXmrRR3QgxBZ2YCzuKq3ugQu1z5PVJMiRA0
7VEC7B63dPbGk/zpmsGEqgVouM1/Qh3gFVJKfUxGClk7esphyg/02F9KeQdXt8jQd0NFWZEHXRD1
M9ZQO7kxvhP/syeWbZK7Qlv9XepVxfDCr3RzflAc+tT9s1hIWGBe1uxlqvw7QWjSfl1JDyN9Q8xM
zQNFmM7qcAq8KiNTFt5OrHbKzn4hrhfoQ0zBceMNFXdYbbDr/e+L08FU9vFdHJnusixKpDqw+vb9
cQhZ+V83KaYIZINZsy7XQ9RfdT7u0ybgTaOAul+CdhhbRz6kIzWdn0cnSjrvotfynUY5s0Kd0/Av
Ob+5/eLpORQT0kI/xxfPbgvWRe9wojll7y8bGkyPV/WcqXVe6pbIZeayEFiG1r+SS1mdBIhvd1Zu
3FhCLriy+3RVHQOCkr3GmRVf943eReqqldCn6cGSbVowRLgFnBpKbQ9DrCPYWj8Pdp/+rev+fmt+
1CyVyTmDzcJ6M3ybj9c0y0uYmMgUQzp19+7/6zrLjgql+cyYIWXMumLU5YBqhbbosKb5dN4+X/7g
MZ1VuAXMSpVdrsEG6T7eUXfvkBcvWnMUWTMbCnh/D5udIEEAZfqPPRbhhyFpnsb8t+nv6mFgNgdP
xjI1dhp3S3h99UT2TjWp1G2qp2bszAIHjV9R3PZgsAKdKratELOOi3PO4F45x6D3AJ3/Dv2RD0hC
bMQptuiRLiWiqoUQfsLSHWRIpCxQ6kJQe5L1/KpQ6zaEnSxU6wWDmsYLQY7Hj/s9evAJfNX3gy/r
d8Wd/xxIIa/0DjkhUmjAUDWZxqmcWLDVNIZjR5Wt0TjyeWTx4E5C/zMdBvQxW22mxIedJhCBGWea
uzwozF7lZ22B2pAbGkjCZRYWEroKbCV6MDyJNaqBAhn2EoH0g2d1Ls88L5O3WGtvHo1uJtvkwVgH
9da1XpIqB5PT4xqxY4ZZ/7i93AepYt82NYlN+/zqhSnOIKL5HZe1Am5X6TdqVA4XaZ/Vu3BfLkCh
c0VrF1ZByIG9Op17s3U0o0zMiQ3GOeeilhlcpz6Y8qjk5g1HOvUsNcwMmaX0uB3ut1qZCgXrF+dX
/hRBhx8iRW0VeIV4/qa2S1gJyPxybe8Y8nrrX0vlBJ9TailOr7/Y0aDvzjkUxdcN61gbkOxUrSa9
ZwwgOb5t6nizyQdoH9KGaP0wJRSAK4Oo0IWYT3c2EppHix1oR/yRXVboXPPQRx7s7M3laUEc1tSi
hcthnuMrwOmUi0yesCKgMH6RV4+Msvxw7mcm4TwDYIu/dYDQtMUMvaTr3xH8Lnp6Q9POhF+jcCdP
RE1EkQm43UyR0OuZfdaADg9F5QMJPQdtcK+C7I+Ky/MqGxar1OztY1mhEtLAfV4EeSz0nv3RKV2A
Ypc545sQFs8F7dwBdQsIeLVPwS8XXr0KPEE4sLfMswrXPx4kxBHJsRvalXJw6WyI8jPgjmT2utQ2
BDGOlqJKX5mf52504CCmpHK7lYLRPGce4xOY77cb3bZu/1DblHcQy/DkBsJUNfU7tuAMz3igG6Xw
XZMSrqepW9cgsjlddKRgA+Xr+F5jKJNZ9Sl/CT5w7uaOmDgiXQnoAWczyRFRqAeTo1W+OSCGzRIc
iwgSA7RwuUQqgtWO50rEQJT6gu0weN/F/5n+r7NborjUYsizOTuWV4CJ7MS/l0Pnz4pZ6juzxmWN
Nq+HxjJlVoq+tTTL7nJ7Bfca1O1vfsD3UPlDBT59FGMNA2qFNuyptEXtAmyYP2R3iG9wzj9cSHgx
z8S8TKqeqzx75poh4j5oVnhyfHwGpnsxT5sXnQLnoD2Afh2bCPg6rGlsfIaWfpLZ80fpu5C1MG12
ksZxt8J5feL8agO/lGSVrV0wPdcqynUYOSU92PH1UNY0lMhgjeCP2REATimQVdKSCf0IC7giGkqH
h+LVs5FV5phn7fFyUIIOQQtgBZuEHYCJab+OPRAWnz1R4sL4FNt6a7ltrifpiRtO1mKdrqAzol47
tV63SEzPqnzejXQFrcLK0Q4qQEIw80PS1IUaFiq2USP/ItEYxyCXs+1WZ/0V+UvXs/RyVomf+Lo3
9o4yLZ7XXKO5/+kEQz+awMCkEulvqj/up6wLMT1GkimSfGCh9gxBA1SrRdWAnTQ8/Uvy4lwDMimK
FhvfUYyQCBpABPzyiWI1uTheUy83ht4zTQhUjGLh7HgTZh2tsqTLi7fZ6Nhz1a+lz/G+b4AmspGx
bm+2nAxZfreogB+Lw9nffIBwzbq9ZvQ9slH/xRas+stxFlhs7oXd5sVpcTWgLKYXo8GKFCnisLB9
xfoO8kzcqz7yKCyLi0GEJ6J22ENE646r7QGbYmrsHcWYTITU09S16I680xxvO2jCArHSpjIHP9VM
tElr++SlHRI7cjCexUTsujAVj7KImAa1jtjdN+RxRq5lfUv2Z/2R/AEUNgcyDgI9P/c/a1fJ2HID
FCPi7q891Ru1TQaHgQ47jZKTN7WJkF6RgAaP+YmB4w8T/9VQ3wFusrgqDm6uuMS7tqlRrzJoadLt
awkpazC6uWrOCdN1JxaL8MsrGMLyHJJWn4RkpqsxxDdZO5SCZ3UrvYShCGsCS0p0OPBGwr/NpVKt
Z3WmjSZ0oV4qAJ13HPiBybiMV09nKryMg8GNEh/v2UCT4P1WFioxMnXSLxzRIMB7XKWHYqXbxe7x
WpJEah0x1TtlPNL7zyGETYng0PW/3ttFJDSZM5T1CkuvL5Ov+3TsxfvzSa8NQv1liCa+SxMSqO/r
Tciba6n7Kvp0AL2bQ9erA8fFzmpTYnQkJMDsycMC4k+VDLC23SChDJ7sjyMaWjNeLO8+lB6khu/7
FikGWebOn5q2xOHos8AWD2nH/wwwbFHnbi6y1SNhjpS120OIeEbc6NKGSUmV5dVPfiaGIsicCxrW
JZj5bsacc6d5/xj0dUNEbvcn3wYZsNl68Q95bdDIv8jY4Z8pyPkCi/+DofYQ6pnxEbslKPRNlN+m
NLxB1XKn8zCfzxGTCmFVqFUam+/UVD1/yCk+tbPp5SJkUlphb0CF84uME4AFR9hJqRPMAUj/gA4e
0utDoHUgR1vZy6PO2DDP/nsULtP7UA4WX/2+xh4l8tXPoJ6nwQqN/SteocqAFsEnQqQKRc76PRq+
jbRtFyyEyU/oxEGA3Pan9Hb7HmX17qTGE0Nzbr8kzGONJQnsjKAq6bGlElxvNaTGMrUhwjWYGwZL
y7xkQn0kysKtAwyati2iyONrvoIcehbZT+UznHgC01inayW8gRJgEANv8Yfb0jIiDwo4r3kEC20w
eDlbk7ySynXNypr8umNsbB4I3/ZQvjRSKSjfOddL3+i9fm3ej28fqDPFLfo0vW9mjXI1GMXMDkoS
EwjLwblk2YRlif8tYe+laK/Rvyqw6scs1ukdmGH5NDSXhJyncgqB+bF41mujdl0nRey+BsuBOgIP
HfFnzvApl8qshhahlR/4ZmMGPjuNmBY8vYU/ibdrW0HjHbgYgU8S9XWQWvDjNkmhIsfk17GmOF+9
cl2vHWXU+cg88u3N5YkE1J/DWwcOkcr5VIaH+ofpO+JCCwHpB/VMEu919k4+cK3M2DzYWt/6YM36
hx2lwPuvdbemXoPbqlvsoxmipFiDkjnyjcSb7JL6TQgk6cEiet1Kf2pJx0n4MDKwkmZMo09LwkUE
m/c2lHlbz4PZWTqK9aFEj3RYmbQ2016xJ8+2TyRM4QQPG/tovJBbfSA+cdcFdoOIg/ODI0hNm1UG
16iK4xnyxJpXeaL/hKjvEVJwMiwVtPRgu2o3gNcL8m1dRfzWN9ffzoX8DZp+ikTWXukvU04Y9rjs
KULaBiaJCMIM1AQ7+h15ylcbjPjiwkEaIEQY7wnfjRbHwiIg36McfqBvy7tg1ya3Scq09Kz7+Pq8
3YzUUyUrS6UVL5TsSNYDCzwB9nxJMYyiqJ4izigqFG50wk2d6T/A7rcM/uO2wWA3Myre8vqU5LTw
jn8lkTjkmFTkhhA2wJC4Jwhhpc4HLFmmu3sBS6OhLl/J5VvBQO+52QgXJCOgJ3csn2AHgMMvmIvL
pm7eLN7YNeK/oOQiPH50Xx1Lc1OocDueMQ2nBJiS650XGIdg4OIQ4pDl0L8xbhKw9HvoLZgHp3Jp
Oc0+u08DANr3SSm4rkpLs/Q2+eIS+h5WgIFc4od8cRoCYZcpXSzXpl8qE/7CWdGxA4pnK1sLk5tP
MuVUVHHm8QIAUmQWWV5Fr5+KbzOHApNYek/iq1IjGo2vlJ2Aw82aYVs3LEYmtwp1PW46I+v3lXmp
RyxEUXZR69QQchaonLUnKo9X3i+6BgesEE1zz6BKUP6w6eyW4MZDptEhI39QHyOO21XSTLeu5YQN
+QsQgR7SeOq1uYgDmyaWNKptQHZdO8vgG6cGtywbKOGaAm8t9JzGEQrU/dZAL+bTWNmbsH+6IYfI
5xrMxYHrS0b4GrRrt9giWwGcdHLTEoa7sOxT625ntXwQSRX+jdFyAmpLFrqZOPRTpgWiV3lEtRQl
ELJbdzXq3x6JKge+cUZJhF1kTgLZLwY02xnxQrb2mc3BUIrxUa7ZwCo5I3F9vEOUtQI/WxHaUEcS
YV+ixAkSW2AJ1PisXhypLv/wgsujHAeMi6eEKfz6pNxvxzmZWhpyaLaM8frBIdVmkwB51cvCTH6z
yZZvdwAtiVzDePNt26dHaAL32WyZUI7YsfxvbQ8mrVgS3a532wqa9ta8hYW9r8svCscoFD/8xrMv
AL6qQm6Wby1UHHUXhRFjRvdVxD55p0ZYPSZB4WKIJVP23IOdd58sGT4jef1I3v70X0Tv5mfbRpXR
UtXwO9KQ6M7VydJNgbPPC4xuX00FJLCsrdeaLd7OckIdI60uDmb3dW8e7HFzatnSu0vSlNZoIyzz
WBFGygJVX5/GHUXcsLbTDU6TqKc9A+qZKcFlKK+JVuWT7YT+CTiko2zBv+4LuqyoEw9IvhzEPLC/
KDk3n4OjroywvlxZtghaDemu9gVw30jbdzFr7LZYCYOsOblp1NLpo0ZOT5i2UaBFwboaCYxKcTlq
ecRylli0UozFOQIFVIX/c6J55RQt6mXn8cyCh5Jdvu2XCceHBv07bub1WfOOfRX3RGUPpDK4vJIf
tuaCSL5zIGs3YDivKoNuyBeJcHUXN4jNNEM1FevkvR7K8fL+pzpTxK9VMZSSIyWIWiyRQwffO3eQ
on2cNbtpPAkVwjpK/iIohYLHIrE8Ms4JCdYMlJwLacucQqgoXTAZhXjLAJ4a7C+lpdub/WPOZajz
k6lBrNzbkG8gH4j+qK4KzCVD5ckjEiMyiGmuwNNnxVgqK/4m+683JG7E6XtEY7z2ZeHJWuo4Ar/6
xJzykpw1pa3biGrUfCdl/GwKbY1FLCsQHeWhV5ybnbQIcUW5t8hmFLWV3/oRh01PLpz/GPt3qdWx
svR+9pXQnWVzs+Acmc7AvQatAki4cwy0C9/4XBM9MX8Z/LWsLNiiEznbbZW+U17qJbrW1fmih3e9
+MHvQSMM3e18byGEHyw27ZTpvjscHCku0A2ZGTwuPViGFGhttH/Wh9TgFVrNOGLocGlJeD89nLv+
kUBm1nS87pWylHJBCazE8485SJ++mRt8bJ2Mb6IKpILsOV8QsQHaUNGEBWtVJm/20MNFbqCVXfWk
yypXXLC1KdsBSYsEZ9SVvb+wMJ2LuAfO5V+2nP+nRMgblwgPIvxkezt5K8YHUFyfjj9ZNMFraJq5
mz3FeJXXts0rNfUjJl2o7+Ldfgb/aLh/xt8l6Zgh/TgzY2cDEti+24lzNBizZOG5mFGDoyiDTgnZ
PxEQ/8J4Y3yWoTfkfDSZZOge3941TUE7y+aiUGPKnKoUdlwwW8WA0xxWUhAuhjUgCO6zuVm3Yy4w
NgXoIzar4d4gzFEO3rIMEOwMLF0UaFyW0KnloX53bzU+ciQTUjCy5+5xQHwkOkA4aHgPUYSdTOkA
FNS9POweDgTMzFuOUpRygIruAHQHsgtB4UeqEs7CWJ1nlF/2dksjjXhGc8nnJ8zvofrzkAwJvxg7
1HpceX7Bm6nY73kOby3OEGWK0FNcoCcHKHcqeGWr8OResIOSNk8ms1a2elqki3sVr7iSOg+7LIK0
zYcuWGolb+NhqIdurWhhshqiMa5wlzJXjToTfWUDANWDgx5uUMEK2N/seo1UF37osUGmT/Uep1Ez
G8DJ8usK6HJ/g50E05QNlloYiEjfXQNLVfwtfUeYs4vfalCgflrjYsmEmnm8bqiYXaz2ZhuqoJuX
yNdPNnq+rTSsOneZ87z/X6wmvd4ITiinaFMuw+3rkGChveuhpwHHoOdGFkwVfzl5w44VWFk9qaQS
15GC7TpHEqVikTkjx8O5rUV1aMaWaHCwcGys/yYCWrkBthFoha19Pbs8YC/wheq+l2Di8gVzSbkZ
f78jTlB64oKFezWJdOxfIMLp8jWVbiPsMA9w58rFT7+cfGIznLkoSz0kav2aEBBTQhAhC83jjDEt
8YbfI3nFwkaKJuTj8pZEbGlXj5ZBeRTXzz8J7XiGS4k7HvacYdIsj5CGw94QzMh3/fNSyzI16MFA
IA8IJ7gpflQOjpDFQFUU4jSN9T+W1kZ8mHRaXrzjw+rkaL6LjU2qlSVeK9IvLwtZZHdkg63sbxtu
HHUFtRFqBr62pw02GrrHZyIpBzQ/7pgQRPxT66inkel03WUBZBucHd6U7L/YcEdyEIr/s+lj5RKb
9wQObvbOFdkQMJiZp023vbUveGOmYqnPhBk6kQgE1nojILVvk6DYH1ijy9dNjIRDWcYGs6MWHYfF
s7SJjstvQLZOSjSTNi2GU7Tmd+EuU2rBFSsJvzEZrXTkWA+IZt4bWNqRddaIUc3llyNlUGZaneqf
A1PJujT5kF/yjf/Q61sQCzfY0FC/eHM7eErNDqUe7sav56NlIsluqcDVAry6GNDmc0vJMys/0Ajv
UIG6pm3tbbJjtgrU8iWzh9jZ+JAJ6S7bPe4KvZg0Kdp/vHD3CzHr2A3LY9VHsZiDm54bZJXudGN0
D0N9/9Ix5etSgn7Ugj0IhN8Blf5XUMmyrpDHDJv4jJ8faCLz21m1M39bUrf6h+PHLd4xHwHvMKjb
dE3IZC3aYlmmpBNdCIe1ySeHCASi/XeSrBz9Ru/+Xp2hgKB+b+beR5tYtB6khYBBqhU36NLlHooC
8xxou833eklKLrRb2yMeNqt0fwlv4acApWpxhNKtz5ouXqcshU+JFyteATZaAsASIAmEUUDgIUAq
XZZ8pVrt1umtdxtikB58yIytiDUV9WzHDHvhBD0pvfFolC+CRxTwKGKir4yIGCnHWWBPhHWNp118
M4Sth6Lk5N6VQPidQGQ/UsEeXbaPKzqH5Wje073HXcOpKW6HVfnrpWXkLk5CKApDr+jxfM/1ISCR
3IxAqM5i8VxLSEPqruuSpC7UI34f67wEd+IovhXh/QWgTXuI6X8Hlbm7L2s+iGh1O3RdcW4fTeuY
eDVLZR7U+SURClK41EC9QWXdC+xMDKVZZumKTxf6yrB9Vq6JdKnZ3SvskPhVSuUAgbx9Dub4+b9g
Jm78mHR4vxrA04i4gjxYbV8SFMr7CxiZ9+igb8edjx6tPpl1pVqfjx6wdmSHWgXRrQnje3HrU38d
NezTAeHGQe1MMd5JVdFSL2h3fcWFOY0yGOr0aKsEPyz9t/2i9NkLqHCFt0r084sXXKugZY5BgJ8R
tpvqNSB/8IdzDlyzlXZBGZDZj5h9/hZE01FFrO6sQIxXq7SAVITz1l2th8t939lqmY1uLhU1xH5+
EMqcHuL6hCJlDxt86T76D5R06REvCPsaF1WnKRqkRXxeJH2vCcy4wUk/bfqhGD/F+6FKDAqWQWtY
+lz4nPXiXzUh0UPMtEZLrpesdCj2Ff1Aaf+capzXbd+GUOpcvWSCvxM5jUj666ULd03tpztdjK2h
eBOPm1fZ6uSDdtHIw2U/Tq4j9LbjZTunPpQJZbc+/wCwRyvp1+6omLayZgH62XWmnG9TZSe6uG7E
78Qfe+Uokctki9NK0D+jGhx2DxEOvo+zsfsUSALdNbn7cmf8sRCaSW0UvflHkKX6q9UmFRZOzKGp
Y8ytHUqXBfOa/wHT6Z08fdVtAeBfZ3ysSU4cmwkbJAIBSturxWgN6hYaxbu6g7N2rWd1wbhHfSgx
bCl3pm+b3u/gpRHejjsjeI36Gk121bvQFL2aOR1b2Nt91JxT3knUZs8oJ6srJpT73IcNbUDw0fKI
NwXybWn9u2ZM/ctXONqz/llicony1UvqMG56pEsTb1arpYw/oNAPRLg1VPzWE1dSIwCqiEMMUPVo
kDaUVUehU0L/EMYrXJvQY3/C2IUhcQ6QDdLsrK/FVfo4PjnFjO6E099xEJDKGNDqiUPV52rvmBhS
PqjStQYasLS57+PwdYgSa/gaKdsWqtL+hZbO1Y5Yxi+exMkYZkr5DNq0PCJx1SVEEud0PRsga0qe
oZ1rZZBouopiR8xJqK4O118FR92UBnW4mOLryEycuwL0RPhUO7xNtCDq8vgG9bcV4LZEHeRssAYn
nQmp18cNXlOpswcBT3gLSC5SJhbKCRsQ4oqeVqCNiT2nJcKEDEEfUysa/IJ/eJjKB/IcaTrGSRa0
i3ouivVZE2GxY+kfJRPqXDldcccdVEudtKGbrpoM7EJq5mpq3jCOHVvwPcQWQH5FISI0GiWT6Vty
/2qUZbUIo/ilU+eXzRWFfQfRiBeglcBDUHDezhcIeikyLJkCmboogkUcndZ1j6faeTWoaT0Y+j27
3gaNZJETp8Xf44qgp4uVXhXgocaSFwWeXM9UGaM7Uhafw20YSjcHlUfalD8R4Gjw2+d8QbAAbAik
pjC0LXCk+uWDovjBYknDB466WOtWvyrnISIJdtisqR4DcZ1LK7QP4xa5Q/gkRVWL4XtQydTJlkRd
zNRQtO+MrKClpAnLGlyiXt6BKgqeGL6slb5ikq9knCK+WVTxdjg9TKrvZL85thej1Vtzp7/hnHDj
fmYauth5fasfzm7cW3YUyPvhY0v30rkR3Xp/y3FfXVOFlr3aThxqhSVT4jzDjaM4IHy+VfRfdjkj
Q9B7+Tho+zqhGBKP/W29fhgONexgEnfr/6Y82iKKp/9I15h0KiKyU8TuyaW/MpYnJmXmMc7uI8fj
YiEsyxmFF7iNLw68/5xPxvvd+rCLvYW6lD7BfRgYmgJt1o8TPr5kH4yq9NWQTJOzhOORqMNIS4I6
7KCw0RXkt0c7IIYtPTGNq8hsqd5VjJ588p51ZPYv/eBJkJnhmMA6hFyZZg2HeW462DA/r0vCsE/8
K0z7Z43UU+tf+eI+fQW3WsJO8Lmtelnl/gUbSecUqLKRF4DfEh84dsCyzXM3XpZ79W2uhMmjwQEg
tf1NFLTFWoVMRXJHOY1NNbEJEEB0wG0wjq5xvsSex2TfWhIK6iyUxcrrZIK+SsjXQO63afwg0zU1
neWy1RalIGu9OvTbASLAmwBCvoZLhLJa8tdRlWswJKFa3XQXpaZvuYUdAb9IzAiWbNUASzV4FVnn
THoZkYKvrY8XQYihRuQeiV2GIP1TxzfhamxxlulO92nwu5CnTBCqSYUbycpU8RrPxscHqBrio+Jx
Kkf6k3yqfK069ijzZW4mjymLe8Li0GVy7JwmLGE+LYdyoF9XZSflv8wg4qqb3e7JiJzjH1ljLiic
rwzGcuHNC4t1eZYdPvZFU106hWuErefkehrdLuD4H+Oq6wB9juTMHfNyaHJdJwW/AUG+JL4bZbJ+
0Ro0p4A5wOqHGk5jf8uLh7UnY5lUxkPvAz0X72bIEuDf0HCK3v/x+WX4iAQN/HBqkD76UJC/+Qds
dz1vkVhqih3qnOQxUCpyNSlrr7iegfiymazYX9tANU2hHNI5nYXxVTwy8YVJKWsvcWGbRoEo0O+w
FtjnS2HP7EdxsYwsklOmylPQWo3VEpHpY8zkn1JQiSPwZyMqcmAUpwVIPkSAGN1hUBjIf8JpAExS
nNKiXEz78tCTcVgjDm5Wuhi1+wTyJlUrcyBbWO1IzgX/2e+SXs+zbpA1kZue6IcXrf/B8C25hFgN
/lKjYRuHyXu8etVmq0rIflVTPlU62dy+DtCMxzuYo/jCHLRtry/z51QL5JaQxgmas2riZHIuWeWu
pOqoO+nATzFpT732R6KsTwB//hbK6GeYQhHo01VqbQqJVS+1LIBNBzfuqARc5MkPlieJYA2em3sk
aScPi0CivgWTFj1VX0IBiwC9KbCoPvtINwakkLHa8CES3KzKkKgYs7Dlk3VZTbdutbI4a51xbaRG
gFhVWhGF/XfVtQXYUAjOBZgJ8GbHZTrFnXSDAcAtx2fvXjkt7IFQEXOPneuyLFFhJJ8WaXrwgm4d
2ln3IBPVguJQN3+db2wsOLqWRVWcY5cwXbrDTKkWzT4/gp0wOEPLFk3Gu/ySFJB/ffA7rPy5f6Os
8DXy8OVNOaAWtb67nsDESrP2sav5e0vRJamQI90YUOxhcJ2yUrxmV0g+F27gOp2CPc1q+ZBp2qW+
6tBdYTb+5dCRJhC82Zprl186QZ1eTGwH350tckQEZYyqt4WGzGH2bBio4infoDL3IszrCtL7qGrv
2S0iq2zLgzCOsYFDwe6O8EqGbNtZ0gVsinJgZ/R8GyC3uk1jKLtWt3g8jioNn/W71PTUijm6olrg
lxVkmhUzqE77Fd33xaWVRe4e0/C96sPBZaflsiCHp7tGS5UOx3rM1tIWCQMvYGXdoVkQ1tRi6ZfW
+yho9aEzPhaP0erSf9WSOA+Xzc4GR3yuaXLIzqFdXswReqNJJky6Z0/N2LvL2S3Pq08xpHHaW+cT
pSE/FhFQSazEqHUCTlrl9t1+HFps0Ga2gMe6k3bPNGV4Y1smbd4t+JoHNxftv6cn/f5bezRvr99g
DbBAYRtpeQ44Qg1+Ux1GkDyWpxkGBh121hgdtcbx5JyFEj37saUcjMJM/fK2F24PlhVP+eY1629Q
6oitHP0zEbdwgt4uMe3FbmJ/Xi8dTEKEJQsBsTC1UoRFroqhKuHcVpIZPTPzL6kjjNvWWmzwKTTt
karQ1huA2tmA9cm/TjCo1JSaKF6O8DshUJKP5m1CK2SUPRvIod+FVzJEOJlKejdypqdA6mqe41Gd
76HkTJjQWf6zsgdAYHElidU+hpmbPAtqu3RJjQHXPU5r0vVLyi76FtwDxEw1cbRT7cxWtHPYdD2o
m6+zg2rQCSpUFa6c9g+SWuXikpi101ugDNlDmlFU1/HR84ZA1FG/aallK7tuxQgEMRELQxp0WyUk
exupnD9vzU0OrRfgDi7G6DkbkHe80wIVLTjZc93aCI8POMEYCyC7sIy7/al4vQn8FYvYbtggSYW7
Qzdyg2ZXJZwYNKLjtoSv2VLwzyecTM0L6drAWoonu8gQDXMJnK4CdJBjfVErzfxpIpv/ufv7Rfif
Ua3oLmq10MpBelT5ZhkDM/e5KS3VWiSQ6Gjfig5fjFeFvcM7XJISH4ungjt97Yv3w9/AUKZjZ/tS
P6jFqbfUgF3RNauOEIP3n/4RYJHxoBWffPZ22Qvf58pf3koERvywDYes7VcWXM8tKtxwqh2cM4Xq
745AtBa+iAZRQ6F+3e4AMjHMx3K55mjtkq+3VBFgt0EuZeC2/kQebw4HragIju23EowYBTWyPPYC
EACZxQWdSBw4e4rulmESaIpRBd2/Gt37Cud+NV8KCgW/sIep4H7k/2sMD6OKgMpbuk/Y6Zrxz4Wl
YZGrgMmbylS0IfMTW/QP7oAssoBIBuhXYc9Y0rLB2skAXFOXyhZAPFh8KBdyu4Z4rrRwZeZBATtE
Lm8VJwL8gDwV8aAK/90aGHKYI9vlLnHBsotfm2kCGBRpnnLBfHF0/McKimDEXA3Shi9DmVkFc8en
ggP7EhBqGeFwlu3PAnIO4psqlbl2aLCTev1J2XkIXtMX2zcinTYLYVn/KSoo8VSLAEDUG6nHYhyn
NLE71NcxtIlI+DiK7TEBFw8ycC42PYgK+xkDaKrf+WsFaQERQeE8uTayU90E23NcEsZpGnq5Quxu
A+MWsnUe2/zW8T+iZgNmuppVq0FbOcVbA7J3Axyt9Pw2JzW+1N1Pks5yPZq27pBHqLp3uoQ7ttYG
Hu5t4byrB1cNfmQVXU1IpuOyp/9XDO31jQb61JBgws+oN9bqggkYY6/ztOmChE3Y0zxtsJx4eA/5
SkHdu/msP4Grmtiwu6RrUXc8Vi5jKLBdVz4pxN5G+1SszlCSZnuGeJzxpdQiU0/VP+Nk2z+ZpcZF
3u5nbCwmv5bhoZUjypTZz4KHQL9hVAnwTRjRdIGLWbBXJp+z5VTrRtCBJc5W339jdOoHhXt+TicO
Xy/JutZJmgxsRWtcVtMlWmaCCMw67h1WHuhhIKtyxFR2kZgrH76CVUlv6asjFjG4krIvWDxLzfYU
1voxb8n14iJCHTWj/Cyn8T0wLcIPaTpGLp/YLlX8djXT0ff4gaKZaM37miIO2GWjcjslzjh4OtZx
SYYXoPwawuJIv/7pYG1rXMZZAZoXB6Z26ylunGFplAJWC5C3kLrnoNc48SZ0C3KNnc8GhiuosrT6
DZDDBTytTHcT1LIM4dv25n7TIOmkPR/+mwy66n/PM+d01ILd/ysBj59qm1T9DFowkKbEmWOkmL2Q
M0DEzDiVWNMIxuD2BTGZAN7Od0j4aJTRNLcrdacZZkqhhtERQsBgzqT4nx73Fxb69swuDPwJOmOk
yhNSWQlmwpwiB2liemuvUSC7Kbxmr9qg90eVtl6sjeZIzGGa/ofht2usBpu1plVtvBUqckuVYXLE
dEhOc0GMAP7M79Q9gwuEfJTUV9tiO4zdcNlG3yhBhxyTFmc5kda48S+MxY4PfZWYRNDeY4Q8Bugg
kQ7GE0nmkORVmy7verQAQavmrDlOr2E+xdJDZc6WzaWK1RWYUxaX4zoa5H0LeaJatnTgrnI+W841
c6j0Wi22/o/FhrDIyiHiL/AAUJpwRnMwWEC1l1LJbD3CZFcGkhLspjXWhzJKAv2SjtWobbMPtvMY
G+ddCa2V/Ca2DduKUBV/4slYY+w341wfK0wnO2/VNhf6lrD6pCfuxlFefcFw4a6j9NPoghU5hhRN
CP86h5r2ap1Eda+HIR1frLB5UaJmJ2s5+0TWgLFDL1tz/ycPKtSDU1bIlUMzxaGQORN+dlt/x0tA
cGDRNna+07NdoFdU2cqMwFae2Lmyo5RCxAh8dEmuQtPd7QOSfl0nq4PwIng4kobGY6iFg+cKc01Z
wrgB770zS0o4/2xVXpl2OhPfhQeFtrReOYPlZ8XTr4TtwqUzmkHJn3M6iTCkiuiYvhZxwq8lE3QN
BLHzjAIfHPxb+BXZjSRLtH6H8nJuJqmtsfMGYF8jDAi5GaZb0mwVGRPbPCCFNewQhEBTAm2PoJol
dMVumxcZuFGKWsI0rYvuPqg398p91saTlW76XAMnPgn9l64QEUn0byQlDqZfDd2U062qiAAstsMh
t/cziuZgRqzzpFUS0wO3cjfj5EcM88NOpmIK8kZXFIuQ2TmEyRiQh4WD0mneA3NXalwD8pJdxv0M
XGzc8C6ADT0Yl3czPcTtW227YR4yH/mlzEnh/T4F245PJHHnrB5CIVXlvctVNVFBMjMsNl0MqV1P
ciOOW3ImAAE8V0O4BQGqZOJkSi5+vDCKhBams+A6NnMaOd9vVTxLlXfrFxjSVwvWd48cRV8uZXx0
o9hK1YWrvP9M9KFOC0jWpji47MH2SmOmntZcYFFXNikTIlt7/sE2E6i5HT5j9zjjQv5KAUkD4ikH
R7Uc+WZdZRHjsj8akoQ9oURmTeB7m25en2B6rdpxAotuTdW337PIZrNyLWlQlyNviaCtDp2KzlOb
42iO9+ApfPHZexFXhBsMsYGZbJFHusxiNZ7/31qapj3Yr3s/mhbvm+VPvsMlC1uz1oCxdIPMKtZQ
efwzp+BgPPN6cn3/Ijl5j9HwGludVNP3oZr0/KjStBrtfxpkBcACCrjlM4VdVr7Ep6is/GPqmj4S
U+4UYkrKwyAaIBfnIC8zrDBw+MxDY5nXLdFdoDYXdMkkzifvIBBhPsTKCXoj1LzitKYyIb0Y/JxO
VHGe035Ut1iElSx6Mqmd6mDJKpx2x/jWp7kxFvFCw3ZVEji576gPRPYHfYs79BHN/yhOd/OGFYq1
bGarwApKpQMFkVI8nwX6rhAV+RxByUPjz8yqDcSqMn7Uu1FeeU7cH+qPQzgMEe9yEpzdnX5CEaVU
rKma+e2v4U6uq9w98vl00Gv+jSyRbguliHpkw+TfYCOmO+6IzlGAWTHHCatNgzx0oM17AmwVecFp
YZ3oHQA8sFZ3uJk+4V8Qqi+tHXuVHZFlXkdf8yMf9wfedK7uiTgg34DXSEYtk07So4qRr3Y/Hfhk
0TgouyXADcKr8rsn4FS+gSjWX99lKKJYd5ZOKop74jNzFrYTMGkOxAk+5KuWkRi29TawUKf91VYh
Vig+CzJR0ts9HtQJtxtg8c72efPMvkl1tDPXy0ia5iodudZQXP0Xo4Zvm7Zagq6eM77cTavmZaSL
KOhc4q/aqhRGtUozUVNSv272lTnQSttqz+0pTaDTJP7VryluITi60SM6ELPKo2fqc03p4TOj1sRg
VVR7XcZTLxfYkY33j64R9row5xfSlLVQrp/0ICpstp0xRZVY/g2RdF2f+S4r/AXRkOY/p+lx7BW7
dZQTXABkbIl4Y+inioUwnnZ99z8ip7SlNUnBIdGgTgfImbw5M+g/U4EOYLzKWbWh+O8EriIgtBbl
SRaTxrk5i4gg21wZfgEHeoZxObJLT39jXj5hpYjtVDt4woQfz1KFSd2x341sR5LurMRqEP2lKLnd
kppmOcEx6Vh8nHHz+AiW65k03sU9X71gVdV9sq/U9++DGk0L4uW27fjKiur3uE1ftIjT4TJn4J9k
I08qidxMHjBB1p4qrtvx4F3H5uUngo5kKhJjn8qHMjrKZvhYHuqZvkME6gNpd4hlsckxLvjvY9um
8a5uY3keNCEfDGIhA/N6flmk8ftRA/IPEU1OILLJVDs+eMDRFz28lNjQeZttEnZtBh7Z4ajImoUd
1NFdsbnEj6wMPkiaCndePI9AqTiMpH5/Bt8rg5EXYWO+k6U0jvGiSkF9XRRrJRNXZBgvr2OZZiUg
t7e44vBOKHd3J8XncMkDc577pcLVM5qV6QfxbLLPrQGjn3rTDGwPeR29FP6rgGowZIm2TeaPYrs6
fgXigdHTpcQXOOYeFxbc2sMXKjJlWvOmZj9IB7r2GSvs1ZfMCbAQ97pjtPrkMxEf2az0h2YvYeJl
gbIr95hVpQJv/GWYPHZodNX0dmyc0HvBiiRy7s0ZzTc+oObefibBPBKF+XPJk/cnIThwEeoltIM3
ZAHzexG6s8OsUMFuQ6aTMip12v1vJBBHDkog4sN05ULPzdBLeU83I2vRhLCKEBm5yFlki5ZU+VQ6
Y7dQDyfeWUSNiK0ZDpFzzK5KNk5giXfd9c1B17WuPLKSuxgMPJYXUJQZS6pAh6c2AIo75F5KAvR8
JIURI+oNaxbmp901kDds3idJo9etX5dYJSomA2n1o3aJ8HrqQxfwlFmhJjN+aY5nuxf4+nGjWKyu
jL7e58qRrb/XEDoDBxURiFUB6px1BQhniVZgYiA7ch9xBA2ud+F78BhICwwwnE0N+PUa7Khump/1
OlV14SB15pYsKVFE+mgf5zgKqdAxndEiEA+c/6jvw+eqHzEuH4MTFjH/wWP0CsLZTiM9lA47JuaH
QpCpShYh0UUzYuDKjouhFuvygk5cGaaRvhAqeJVONuutnuTB8kpBJUJV6hStlJKn5DWmqPigiEls
ZaYNPnFlnlCtvl2Ne+51AWGNi19U/4hFGgY0kY1Qi75a4DsCEU6JxXqitkAe4ClgHQsdiPZnO5mE
Tq/jnAqwar+a5Hw9RlcYq3TV2vD8QFi4DY2cjvkbi9nrlOM5830YBA7gkTw2LmsOnTrrgjJEIST3
o4LrBrRRlayhEdVfTxH2t+QMxY3BtKsjhD82g3xO/JB+7rGpFB0Q9ruA9tzYOOvb+ZvbA0iS1Tby
QhAGjxUQ0ozCURQM0PHZZbbvV0iuXjOM1l5virwcs0dYj4AbvLyycCQmg64MW43bbdAuVwT18ko5
OYfpY8kfDcRaDNz36nwOG8fYdVMr76IRpVM8hq3iYpn7iWwfG/2Crr2+0EoerEhxdxBieqMqi62D
mtHdrrJVx0rd7YwxvjxucI1keW59K078GWXfJ4KRj84PTin0aofD2SdSt17Aup95JyDyY0VFRGj4
alK0MRUIYaJ9stRtz1P0JJbOkDKwNcdcHSHPAcRwi75InMqj4hnNRnq34CSpwRDaUinWkECTQqRX
nMzA2FKSVsZIMoMN5uaxrdWhnE4WnPoJiT9XeNwCppPXM8GGFtnBzXGyoQJRCFSPb6Sit6nAnsKJ
/RFSwmSkuXCk3q7lmBNhEJ8mhxjecCrlEd2Fy47dH9LdcYkCrLjWDYHGseABqc0NIxv9MI6r3OJH
WajRvLBFUS2NTnY0BOVA/9hoHH3nVdS6vgAROpFhmzTS3Hfx7mmogED0t8iWpk59mdtT++NJhEPy
FvDL2kINY6uk/HUQKEGcbpLJcHQhjI+9sm3ZQQnPi35NQh0ozRzEPQA1tu9yYWJ/oWgrFIdPTwu/
xD5bbzwMovOIjh2a6QF+riTDHSBXt0vdW3wdDRTDshPbV85mcqRkpXJ1LXbtiIXnYQ+//3ua+hyr
BvMjE5gkTxLQWrTLchcSUaZ6GuZvTVe07wKO9dmSSzXlwhi5RmMUKSO5oMujRaUE9WnjdEZlBnN7
aoGok7hWb9PSUGCyimF/PwjEl2U2+r9n41tN1gogb/uO74/tv4Z1O3Pf8KiP4ioqZaBLC59WZ951
QGvginIG9SkrXWVRCWk41HfDZwj0tySvJ3ezq45/G9a2s8IXXT9lXNB5bcNIP4hYQxJpp7iJRiOY
svqOBNK8Q1G0JH6fOJaINj9TPz3UtWp6ND5XzUJp5PgXNdUf/P2+j5wvE92ORcFU3fsmL/jtnsKX
fYUUjgp3A/y9IOnyPSdagJgJhkf+PcG7kAtSvV6qWPAAceCEYJb/dKP0WaL43LUQoR3DomG7GnKp
iMdPrtQGPiN12KKZjscScE5oJE8XGGJQJNnVYKj3Wof6lV2JXZN6mX0MX5Z3mH16+niSCNh5jydD
/iOTdGBtkpaFbrjqQpX1sS/n/Ks/nh/gv8c/PmaA1OxOg4AoZdLVbgeblAUreJ4KKUNRUX0KnWSL
3CMNk+NOY1vYAPL9JDCvMAMDfji3lz7nQ1nzIDFopFyiBw+kWnmqwhabpArt53fUriklv2RThVas
iSVUgJqut/jNGerDKjXEvMG9MDL5cPaReRsqFn27tPaYBblvPY4MUxmz5fO+LyuWj7qb4TFRy1+b
jMK9+zKOociBqDfHPT95REGMkVq2F0NMcsA/mMYRDQGNhTz+B8UqFw/RqyrmtXyqtTYaNH6qVT4+
hHg/xP6n21/bjZ1c2FVcaqR/Iolf39sEH1fNZEDFBfATzfSHTcbU70XG9omGWXbod5GpSCadWQXl
F02DZTcsPVAFNGcPfRG+puK4y7NxxamwvJu2lp343uh/hkQJst947rOJDtRbGQDZFladY/Ae9tDw
bsJSxMXX4nmw+dLr/7rXZtjBs6Qhi6hzgprzCfkTwErIH7QP7tatzbGBm95witjRlQuOIQNqjVw/
TViBLPXYIyix6b4vbMIDTr/raJ06S/bhgXWlM593JKw57+I3B+igUJIyyGI0ndcBgeWkpN6qQ61I
keZWb5dkD/Z/VD8a8NE8YHbnBJ9VELxIjUnoOAJe4LVSMRjMaO5GDEVPLp716Rs83OOJywa2t7B0
lrHx4TR+tobZg8mos+vEjbSXlUpv9IoNNDgJBY/FEnZqhs8e7MDuH9rP6Zt6+4iz4w8HHck+Vzr8
boLNx2eItmaU3xVUWqgrlonj9ODykk2yAyQU31MDFZfGwHBy1SUDyN0QNKQWRWJQxb73Ku+lB2FC
N/86UcZbpk9+/tAmpHOysnD8P36kZa7+MAF1wZ/MfR3SymwYdYmO7KF5ps/4Dcmc4ol7+cVl7EBu
jkTy7ZWgvldmK+GV43+OZ5OxsaQfBjPO34caFG7uBpVunt7sIZKeB7eTeCd9zSqnNkN9BYkNZm7w
w5DcHlWi8W7+WTUP5cdu0KGqa4cSx5Oyiy2+N5mKTRhilaaYjq6Mh9djg9QxN8oqv8bay//8AF88
eoZNxAaZkSlHymEPB046btDGmmipzXSH5XOwIPoc1YFH/uj+oEF9dGjks4yYGjvgiLRhCXkA3RZQ
6mHVDTKJOpnM6DRyHmini/7Jhi2D+tX/wdpCFsf3ceyMw5W93ps+QMzDCu+/k2KddK79OPGyYFer
gObUkbOC+IuPZM72CUsCvV5cYA4rMw+ymaMGIREVzT2Tz7WreedYKponGAdQtQEIY0y42VTRqt2f
MorYGSchtsGJexSK1xQnZA1d9pPJgX+OJf1GMtWO8Qr+gUg2tyBOYP3lekwiRWkNQGILW4ZlI+kv
Ozo4a0RHWD0FO0PD2tehp+tlU5guz7ZO7h8pQuqi9pLCKSnpQtnyCQCYTqcTsT5NNXJ6wAlwqb6k
+k0oshsBf2JMJ5SNvpHOC1H91JdubAqjAXDStCmjnCXm0DHJwSBPa99ILUZmTt4daJIMyk7VCbfr
0Gy/10unuCpotu5N14saJ+vHbXfwRG9g+TNEs6af+0Dj2MTwjrrjkV3BrVMs1OSSNi4PsGs5tRAv
+vAI0I5n9uDAZ/Ro4I0kPyCwAXHdiyEnyuLjAG5tnoiXVRMochRSFncufxBkWHV5qcf6AhIXNlfg
19Xfke8G49wzMfiJUx6b5Nkigsj5dEPD1oTH9fhS6+sJWidRm32sBx5+7SKg0u5RlrM9/pVgASoc
L+K1RfzOo68lXVmD1jfXEcNcfdzgUao1hAI/WphowYVy81Vh+pF7N4F6RjaXYxkxFwGCWdRxE4j3
ggtiSqmKHbSUq2utVJ8GzfmH4Cyj4+pwcoq6ngZwAKZ7VgDlqXSOZwnkCdV4aFMp1ncW1Ktcp/XS
0wquDWIaG2r32YoxAW7jKu9QSDr8A59B5QEC+pi623yTROyL+cDPVo0RT23zZx7kW3+UmUDJ1j9D
eLAyd3RJZ3psmpZYxV+lhY66i9k/b2uLnzfvZMSmSJDLJBB2PfFEeVDlciSclep9/9sjirNmu3Bq
CWKQlmYL8AH+D6jRIp8Gz8adRnIJyAqaV0SwBPt8+vAA9hE2bVZDQz7Sw6pZh9jlD+vuxzHcVvSR
w2bNEJ+53XFgqdEUYc95/nS2bfUIyjZRdjjygpmPUEHJl2el9sWcY7BUbDQ0K8Ix9/YJ8laKf6bk
dE8HLral9HgkeW4x05xH6hUKX1oQ9Atz7Zg8UWvqR12F0Kf16bt0zemS09xuWdHcFufua3YzdYVf
9ubdhWqTJh0Qk3psL7yQw6/MKRu/IIXuaHC1kOBjdsvSXtdntSQ1Fid9wvUle/ozHSbd7zH8C94q
hKs7+3X6eBNYT2e09LFOoWjjqKrUo7GStde8GsWzTmk1tecYP7Ks7MaAk2fXlcI7LMVT6rDrpnuL
7pHLv5HGAbz42aPkOISEyg3k/owxzJJimENZf7fLzaBdx7Dhp2po9drGTY2dkcsh1gDuINUSkhMV
YHGZPRyo0+T0xVAyUVoLWwnjZbVeOjCLATaZPnHpVwFtWRz8dHG/A6tU9T2ymBFQDp0Uxn2au9RK
+YVgd0mqXYzK4hq0GyLDrlTdcRovXckfeMPD65EYpVaDlKpph8Tr5Cs6LAS6OCufNK2SdjPeKNLT
PWS5TF1YduAXEKpxrYwxcSdk6W87M6Jzi4P4ilp70dZzVHy3nnOjSxyKZQkRFvePagldTwhSpKa7
W1tqrLAMQ6Fqiop7SWk9T08JyYftGq+jBJIYy4ZImjRB81sQ5OjkYB9KtkblVUttfmW4+hhkVnsa
jFZ2KgY9HZbwSpW1uLNErCCfY/vnHxwJ8JJEIamJKrMoqSLocrvYy5jaTG2fyLggHqzPrsBXVLug
Yw9BfKadxIuilRcdcXFqYzMLzd0vVpK8/yByrUS3qkH+RDzGcddNCA5Hgm72TR5BO19uBeTGXZNu
yhJ62V6oCGziiQ1Isi2gYt8IpUqUXlOgWOeD2Omj0vSomDsNS5D5QYNW5aki4o2LhLBu1NJCdSUF
xWKaftqi9feUSQ+TnFFnph9yaIQoedhajsjwg86WQzDQWKCwz9bYDCHMMYFDFFfqpnxfKd8u78xa
ovc8z2W4p6f1YaEUT9mjNEIBAtmeog9ez9g9ZOsYJwJWuPR6qehg/nsB3m27vB9wwfYZ9gGC7hCQ
q9XUCX/+Zw8igWCP9XBkwCVgwyk1zCu2kggbKQbojfOOlK8bmls3ZcelyIyQiZm7ReZxvvoN3jvs
i6QyMCyMJuHiBuAx1COE8/x0XlP8yoEWzcZbXvV5A2SJTfqo3V/bEs8RKpUFOrMbhUQy3PApNmN/
QgjOuZ44UAV79xbhzD/taupqmkhVevm1P1sJ/6mkqG/wTxzhCB27WRTbr1pdOvYeratjhwZiOrwg
g4wc3ZvJ5Sg3h1DaFq4tG+bWX8D6goP6N8peATHwKorlnIT2TsIgx8riDNbWfqcmBFob3+yOBrjo
JSGbbnTx1+MsJBLsKS8JTPDS3/u6F9Sn/x4gqsllMlOBOzIau3j2vq0M/w69GbV6axhQ+4eCNSeS
Qg5l693ZjSvaiFllypHQTO3A/HmB1KTemd3FsVVdUPLLJxRM8AXuvkZwYw4fV5lGjURwn+tXjYkb
HkGmn0635IWOna8/1puhtJcUUjYcHQEOw98bi5rFMcJRPYeveEtZEWdinYJmJUdQYp59T+pQLLrg
+mrc1+DBFnlO1SwH2TToEQTc+SMkT3Byzzmb5EgastNZ8GjEvufO5BrqvhFnlu1XoGMs8H8m8YJm
SfKoMhAqXmeUEUc7EDNKYIk1FAQ8mcbc15MohOY1aiYqriXpZ5HSSgotsZ11RQgoqcEhMyEdm7fr
CUcYhsSj6dLFf92PUD+nIgwwAzlDUZiyQnDgjVq7kzZke1jksiMkhXjiPVeF+Upg2aJkBlXaeskR
OG+zDtOkaM+ZAg9v5gy7Ad5PpkAZZKWBWJxl0ljUbyXoo7pvazDZpXxkBOjj4IDF7hqjRu8fADyR
wpKEAwpXrn+MmXG7e7N58g7SwlQTiXraNHOrA4xh/eS/vK+6RDukgYkg/wCGJ1A2ckGnzV0PFt1F
8ctJc9+HdxqrPxAAScxCulCMO8y9V2flQSIwTbzFPZN1iMyLc6pMw9K6dih7P2L/2zt0c+WqDnTT
IDEuSZ40/L8b53w3NlmSryLs9q5SDGrKQKSxgN8obBWvrwhiN1XMckzjQtFCNiylSCgdmAK+2ETV
Rq+4gM0DOaAuVDWXRqHsOqHUQwMsTeSVNnKnV+3gUpqbJweTKqIyuJ5lYGfRWy30kU7mW3tXx/7M
Pd+qWZ+oTswkxO0t63OrwBJM7c4SWI57MmOxJ8jg+7jtohFwhmTLxltas9vqwoeAr/FmVj772riV
xrXOESrf5uqeK3k+I8GX46iaV2Yxf9t0lnRatjv8SEqoIUapfzfotAS0WzT9qoK83JiswrFEPQlz
8nojlQ1sHKaQSzbm0yGYCia+VNdS5EMH3V4LoL0aeZOrKM1m10teiucopjpadTeEKabmbFqa1GF4
v87zQq8Rtne9GdVnP3iDmkioYvcZPzOVV18A+ZvMHFEdsE474U4oP3P/DLNDeKTI6qV4D895xjxy
m8FY3rCJWZwTu8GbMRx3Miyrjp0rC2ylpcK9mF+p2AR2yI9OVEzdqMMLbu4j0EekES3oiZem3vk0
V2eApmC+ZAvmxWocK8ljxO5p3BI1YSkQVPPir2wqXr02D2fThBBZkKDgyg8Wr31/ko/WBA46mzaM
k3MU39uVMyrx4/Epw9TKQju7+bVSxofjm9Pkc5MNm9igCY1uEL9xrOLGdLycpbwTR0Fvr7faBoFp
kZO5luTzOHIrzrhVcfZSZyUIJ6tuAtqN7S7gpDwVdqG2AFL7Ngjp4Sz6/ph/U2eoMadWjWXwSYiT
wUHyKZiCOHow5xLaGA1whK20xdL8EZwJxQNyXrzX3wWAdmdZ2Vbkg3bCit9juVvXx8qLp7Y2SZeI
/2YZRavPllR2yKq9mA8o85s8Hbgb7pxr4602aizGkwvS1EG+PUD8XF0F1ULsD7+4WVSOwLyF6JDT
3h+AvqOFnSCyt9nLLBybyJdJdGZ6BTxMafvH51VHU1upb0JFI7CxWWEq/YFnp0wMYoNK8Rhvr4Zg
6r+58nR0oM+Zd3Kt7eO/fUgXVGQZ4hXnnG4ne3TyLy0mCIttq6TQTLxgtMa5TtPM/t5kthr6FG1s
X+Fn9zIGrMAcf2GZ4Cx4HOPobCzAwQ9l5fa9NzHU6BPvkvUm9pRmzMYi9xtDb5ix1j5FebdvS+wS
U1m6p77dPscBfsw5tGxe4o1L8xxNZQ03DZAvAVogiLAG86QE1Cw26ngzzksLg4MoW34c/a6H3asJ
mrEn+9Mrs9Zpll0n47o4BY/ThoVPeHt2x3moOJlFQjnySSgHIbZPhCIk6UPrbk55CX/ootoMD2fk
c7cJ8OiW4tl9QPnQJQYca5/SK4uz1W9e4QPuFhYQwC52dK9gwIgNU1NaZizeobYhKTkJQm+ozhH1
1vO1F848LOM09FA+XZMdPJbw0yGFmmFE0uDKYvQol5ArsR5cp175MHEYowj/CDkSCQ209gR/wUGS
T8Qs0kxNwSjbV/AXFIECUhetc4V4TrQCQZXPguvgcWnUN+6EKgT+1J7w3d5MnaZN58WXTFtxSlT3
vyDVJExTnyaaHWh5xIo/qVZxS3r5Wnlzl4v5jC/5DR5DMQrHEKC7K1YYr+g5y8SbddOI8F/Vu8m7
sgxH1enxjLAF8V83vJ1PYDqO4KgucW5Xqn161SiFD+QjXm2iu9UQQH/uCcBgaP37dpou30xp3lAU
06npVeeuQtkIU9p/IPp2aVvFRAxfOF9Nl2r30AO25GkN0BFZwi/fz9x2rInWPfMlq+A352hz88st
bayBjfU2o8gAb8OCmiZd57UsZz++Eko2Or11NpVwgJhuLe/0TWFDueEbSxw2bM/y1Xfp3QHI3pWu
bHciKDPWIAi6mj/i9wISemPCFe8Tin3QazO6f/YNwOEHDBxzY4eVpkEjdHiVGV6/TvmzZCX3/ERQ
H2/im0SmFiNQWubWWBfbyQs0lLJMNhrNPHX14TGTelFTepezzcuu2hjuRuz0Ypy5xrGmWhWHSQFQ
sI+Rhu/eCTshBQO8k6CaqxU03JOSVBWBWwbGnAow+0olVAE6i9drgvwmbtuja0Jr57qgvkwRiECF
F4l5rUrA960HufQBkUk+cdPZb45Ep0JlAahZ5nZmdqW8o7oPN40dHB2QQJ4Q9JYSJvW5725sCc+T
rDt7vYEyCdAmyAaSo86ZeDliYryd7g8wxRi4quyyTFq9GC0dm5GOCK/XPuMM4FQ4Mqu2+GvmRI78
pHx5Lmb1+ZPuzm+NlMhftBr5lown7TsxOfR4/H++4dyXR2lT8579Y13jouhyVXS2JotswJ/dUMAo
o521u0yJi0wIdqWLGubFwOhUdcMYGjKTi9LqmaeS5aF+XsSUBNN+MASmhltjeHZmthCQZ1n2fyy1
kVr0bU3poN/RcDxCXASdL3I/xSH++yHcjPODYoezYjU24vMRBjK+LGL1c/ql5zpNfZ3vBJlkr1cs
7f65q8ii3I2PwAUX2VHaT3JePX/3s0doKfoy1mqjMHQQ/I691LRA3mkgWtKwi6/XGpuVyVA3e8F9
HjeQ95kbJPuWU3nCNzThT2/tG6uGbj2EhAE0GCYA8dKn9aVovtwKUjMICfPYa1TjcElOjzfNGSWw
ozcrzkI3fNpRLA+brE3b4Fp/Yclu+qSmHg5CSlUpHBi0zT8/lvU/DF1CBeI5R9WO2N/YlrJZOEKu
e7ifyJjtKuFLu0IkxiXosUEDJ5GtSdtS1IX+9Hxm/EIDUe/YOVPxlZC/FFX2waGFAeZHzNMlsT/4
7NLu5DoZkQaOOrqoLco1cf9Gn7KFuPYa297zOxd0KBXW5gM0GgUPEM5XfNuGI773kGOtRwLkaYDD
os+/k8+DpmFRCn8okfh7kMc7QlXriKZIfr9GO+l8OziBZWL+au1bcT4cS8ciVk/5kpd1encLA2w3
gZFx1Loc3Gi/xjBZOSNHtUSMj721R/vK9RGLGbr3TYEU0U0xAI1WYhuRyXAgRNR8OLhxSs+BeStJ
4mbbYHdfzzSnSQIhVkB0O1+BBI2rq0P09se0mymoOIHaPMj90AmqJRvCk5vU8qhWH42ow7/Nw1+F
uM5h8PQ8xfgmfl1KcP78SEKIYoGKvABbQ9gxQLe3CP1rMH+w4LtiTzX0gEAEyqNlVb8GvJbVS6C1
xa2t69vUYIILe2rpchl4hAg4/N2stKxsGdWA0InJOA/ZjHehBki1vzKpT49J4Rs0B0WOY01rwQFD
suJgmi06PsXtmPMrcyD1OHbY4XlcxYOgReMjiopxPJXcE/rPdiZMAtiaCmMt1c+aOyKq5LZm/eDQ
TRpWkMDGoMxPSFglms4IBHMFHw1D83fwatpV4i2zFwLZxcDo//tdv8n+lt7lMc+D84IN1EFOai1v
JSLJVAN4R4U9gAr28i57s/vXgrpWC+XiZEAs7KQummgsSt0sx9DvTgkBn/oRs0+IYpK7ZfxWAJgl
Q8fbt/Q9RrcHDUt44YnzSO44zSHJdQO+4A74FbcFTCPiQEvN4eWXxPhXR2xGt9/JTG+n6ibHtbSH
D3pWZkoYhB+iLthafrptw2Tg7pgM+4Vn+e1LRK0sJ5uhabHy6s/mBPfVdmX1FrUm6O4LAH7y+L7z
9fIrCwlUjgld7+X7WHo7ApizZgJdIa6L268/NjJMRNViGmZpu/x/sPA8Pm1S1oPeOnkjkSEdkOIR
3jkZlDaeklk994DudTHRiYAgm87YNKBdwXTRZONHuAiVpG2U50iJySoEbeOnVstiY4mPEPrmWDhc
vRSX4rROJ+SdEUx3N0y7MLf6ybKEpMT5pwy9yJHP+q6hVlP29NwiS3OAbSwFW109RRXVkZ2lFcWI
saIsmZ/9OWhib4EVpFJlhGto2Kzh9hyXHF7uJYZgpjOcyRtR87+RKkLENatafZ8lcKDy+DcTcWxW
gCHsrRCf/xPnm4LcAlJ15WR3AlA6KXyVXYkBx4f7+09SurB9oxWcWV7gBhmr93rZ0DvharS7wCiR
MTFX/9FPf5OWvdOLdG0MtuGr5yJocF4UzLg65DhuzEHSfXRbU8GJy7yKcz0+dMappsk4/rijjvk1
CYnSsKrvLLCYBLg/o3xwRc7A7K8IUBlsLIbGQFBvXt/fGIUEMT5A7LUOcKfnCZZDKRAQH8gmt9Qy
Dwmzfi1qSaXRmOpoFQQTJq2VyWDXurlGM1Nym4ur4PhJclJY9+tw+VmM35NekGJImlp9M6QNQVnI
zGMGoOtv1KSsZk5OxZEFtCiCoFmdXJajl0d0XJkt5pJe0S5KXB4E0Sj8sTigdzwF+9P0apHhiTAK
WUZA2yOxQ8wY2/+bkBxokJId9fn9t3/9uwgfWmA22iBqEhezmnnvctWKqlNrbVtzODylVyK3dm9d
qnO+AiveqwOwzyVOMdSS8Uhn+t/7ohQuCrIFDShtl8dbAxpaprpDYLgqp/0c5OpyOysPfdTuOh05
FH9fmNwN9HvII6qkR1KuBG0LwVCOh17u9VheP8yRBKe91pOq9I3IDYvqQIPbABGqksbtNWzElyNf
nLReBtMRkC+1lcRzZ/BMPq+3x+eX/T0ut2JBQ958mllvY0QfP2R+tebQhiLT5ijivZjEI1TCGfgc
xLZE8ClRVs3fOA5b79aStrXeppe5oyBeTdBR0+tm90JfrVDUoddd9nmGJxH8k7ZxZHEY0S9BSYHa
hlWJLLznblLEw2VLRr9wgEFdg+Zvb0zQpX6wCEe8V/6qZTqeT8uJyzPXKpFXbIOcIWrZE//uPeWf
3+ck7rPfaSidqlz4FYhb3nNIEwtOlfcnxfnAg7CkIOQDM5zGRZHoFNGOZmi9a+oq7JjPqpV5H2E1
wIqjYgsC2PQWUb3Kv1RwHN2lwVVjxeTuw7xm67ijEPY/TXaoWNZp/Datyx+5aqU2YUiYYpayzRxC
zzMttVq24xwqDNJ2LrMUMTjlkiJBqOdIZoV0Dph2MwCfTorKPpACSbGY1Zi1aYt5KvIplAZ7ft0j
aCsezdKwJf7r8bdC10OKgQOaLpD7CG5QMIdCMyBjU67K/UI6sLSK7FA4TMtPxGVT7zCftCkxf3W9
aHB0/oQsNcP/mM5WW6ypbe1h9ugD9iPygDob2UCeU8r17PFLpSjCm25oVrG9pspXsuUqKg4cbcq4
39o0vXXP661go/tMhGVcgOQzPkfuTDyDRswkdUwajN1FgJc1iAPFDn39otdFMVpp3cMN9LzHUB6q
dgdlqPxK7iguIVpiJUx6BuHlR6w1+yiWw00ZB23ZyKVvxuTZHuj71ZBEyiXGT7iq2YAxLSC3wFkV
s7/40MwVC6i8H2jsu9khoJ642CvHWGxGFaJ9tiTaNWnb8Td8eBc/RZGPBT4k212LD7DA7KgkopMi
VsGXcxjs9kklkKgSaOKN2GM1Ngdkqk6piZZgHNWNkStk8OrqgZDGy49wtOFlVMPyNs9nw2Jk+jJe
BaFJIUvCqCVWdskYS7E55s4gqaShfP5eZ9I1wvzo9E7wa4ZCX5BU9+YAKgneAUUhc4rcWTTXRANw
cuzFI9vQm29AFIvzJ9BgAu+iqKaXlICzPiQv2OGjXkVM8uza5qODByJH29+FTRV8n1oyBo5VyRFG
Uph6X1Xw1idHt48ZkmU3BOvoSELkxB+RYFASCEYNWercH6mTFkxZRTmIb7xGIwhTycE2k8sUEbcO
IR9kuUuIRGjzeEGUHaJcjWLxLut0PFmYLNHCdBg200jExG3KwXRRjJ5z7ZcxA24rWXK6/TIHc0MS
nnCt/ZgOz9ap9bNePdaXWCMA8IbRoeDAQFO5rGXY05pd/ss7A+IsXFNSzR6xVQkvPdPIjNm2wH0g
TfTFAWngLeh+qfz9lQWrm/InJ9+kGQdXju//++XFFDNwhHbi5KtxOaHZuzEDQXfgh6riSJ+L8Cxr
HvBpitHu+A0UF7dGw+rwlf6ApH1lvDnuu1GX4kT8qHIu8YRd/PceuXMfxTtYlql5hi5n08vq4f99
akvu9Zl1wBrsFjzPKhvJgU4WM7suLSLKa7fIZFJYyeEEKcXVQbo8j/ceslH6gVm3OWnUPWjm8RYH
2ft/8g0qGDZJEp66WQ1t4uxtaA+yATYBU4RIBzJ7k8AQH3Mxcsagvy0Hy7CWgLl0L+CStNZOhqMG
ZmbQIczBx/I/gmIIF2yviUlSMdd7iRlqwv0cQqDojCo92GH2dlT+VZG8gWQhuMuQ/HptQLzqdawj
jCpKEHXai1Pzd02JTYfjkryq0V0n71rVAGOMn7GjY8/mv7NVxtRtcnxIjupoHXCHQjOCphDCz1eK
8TH9av/JJ7mSpaNBbjD512mqAsSOj+ArKsNE7qigIWpUHC4pVtOzGaKLTXc0lTMoGA4tMEQqPy+4
qBJkcNZPCm7pVGjp1Hhmjfx1fIMwmsz5SOGZusHxjjw/5lu8ZYysL6Qt6USkkoMhU01uZFjkBP31
AXx0TJ8PqCpTf1D6eD5qdFNWo2OEWrjWqJNpIoBs7snfFVn9Lhc583TAxfoweiOxLrcOGw9xL11F
Rs6wOka3srimIHEINXtNZHWYAIrxum3aqHukmVCPM8Dl5Aorum/x46zb/UKTl/hNVjFOw1RaBIbY
HE8y6OPGvoeKYK907B8C6mEsZtgM+Zu1HkltqrjeqRoUzApvB1Ujg5dCeN91pPsC5pKV957PnYUH
lE3sHTcoH08fbJKTbiV1Z06v2Tt3qkiQSZQyc61HX6Pt45+K0sA5iK0sIV+MRjBR1z2thJYsxxGe
niu9ntPABehl6dVo3qHNMSLtGanBEw+urrvTHJHJmXm7/U8Z+/YD8ciIGCWsGxKcKRH0ELlntm/w
krkCo1+fSjJKRSDT7ac+3puTeGNRXO7JTbFyJzmJsZfsrpEW5mBYHOhIQj2BuzILFi5y+PUQvSWc
Hjaazs8KgbevGsF1U1molzfnfcyfjmAaz+0nM9/I207/uBtLA1Kto4vdjkgqTTTUBr6NSYwM7yfO
OU1KLGlm8nglim4oMWAyUnGBegDH7ho2C4SmnsT/0nILT/7kK76DTgMkY3iVL3g/zh9LGmHFYhXr
yacE4w5mzQM0I9zRKhwsFhQQkjCi90ZEn09RLgYIYaZXrihWgZsR+U74Xmfy6M7bwPhJwY8utRzR
AC1wSH3NS2OJX+z8HvnHvLbegMODSTeKzZq3MYk7j03H63IqjxwqkwN4JDYc3lR8t/ne+qNNIgQp
KxLvtiA+tVeAwieINzteJAeodpXcJm3ZJDhJrvEptpFIFw2YvxnG6j3F0LebLiklOQPTBTcvF8NB
ayn+sLdtRacciUVoDi1ASAvobpDn3layIONTOGSmNYWdEvjwR9eKLU5Ow/B2itBgAwQsgovo9ay2
moiVyX5FUd3OJzeFr5rmyz61wmnZbjEK/PlYxvy3FwFJv81WBWv36WqOdWZ5opNQ8t6oS5KzFQMC
MSvviH0lMcDiA2XZ9++yZsTNTC3Sd/daZpW1t1zJC9HlF9qrZyXQDloWFn8mRz1dU1ZVgMZ+xJAi
NAbM9TRAbwbIzhaNKrJSaELmeIAb61hi8irLO/QtxNyaj88mvJScdxiZ6vI8eSqIqf8ntWjqBrFl
iwvTt+r5jXFtssEc968WhCD0xmCk7h1GjjIcYP/Kod//DSNQBF33E9lGt+ILYJyY5Vx0osLfWPM2
m+Se+jhH8nsiaoqld9Bo8hb2Ndq6ZLZCNji0ZqbWYaC1roMlsXCkV4WEvRR1nREr6CXwOzPsSzhB
P0kd06+o/KUkGiNaelYZsKySCS8b3aYi4YCujF8VXLnQfF3asXarO7SvQbBl52H+IFDivZ6SU9Qx
Mrh/X6t3O+ME2utuBH+d8/pgMyiWZD7sbO6//akUKfKZKtepf7RjDLu6c9w632CT0ZLTYid8bvyd
Y+Zqb+WRowfpFtbnphpy85+Irz0oMipjG+uJBOPUtHYi9GOfViOC8Jxf1ENzSw5WewZbhaoHMZIa
xyz9xPqL4bB+rmz+3z+TbdybiGtCfvO3sQBtIr7S7SEbhKR9LGj70JmDcolmMbSlUrD02aFAM4Ue
mX5c+Kn6DwmtaZNn7E4Yv8rnoHcHlMF20TcM8gkSoTz0izA5Y1W5Z3XZxIQSmqm2T1GU1DAq4K9h
CIywSrOuVBDF29JbAN5AfzXYyDq2iL9UJb3u1w1/ML1zHfDtCIcCE/k4WrOHMsl+/3EZwJvQtwRy
PpQtKaRbnltqQiV5I2jwTga6OnWTH4/QpnKcJpQVMijPnMEjxtyhnW6b7vLP6I9RdHQcGcsCzBou
Ic1ujLTRycPZ7wwISIzOYmAAaVb/xaW+rm5HUUwhh+TLWdt81nM8STSbafE7jmFXLZngBtZs+57t
/HwSfF4CkiezWwedjKSuuxoLKHih3TU1AZGaR5Bua2q5b7kX81tu4hBed914u2XYm+neVowe/mCg
K0099LW2UyFO1Fmz6nKuzuN6UHSikyIIS6tsf9Px4qhQ9X/CbcU9kovAdcS2byyb6s0r8XHg+Ry+
BnFuDeKIToxKxChGbIM37OKL2QKdFKeqTvGQYIWsYH5wvcPWyIgpzvGd9f00cXO/Z+FVlLJSuwQG
ZP9EAIsLcLHWfIasyltTnKx9p67OhkngvYgIG6dL1GBPxXG7xaq0cm76FNCV52m+9KJVvWhV5Zmc
EMk2TYBbBJDuMgSJ5KzW9MzebGAW4F37bo+gUC6zdjrkWLMua5RM4urJVg8kC9Agk/ylUETRNpqF
KJAqxg5L8pzMDRwlaJ3D96Z2R3pqovWVZH5vrNMl3zP8u2AINHIiCy0FgakZ/ejGKLy8MUdSMdVq
us9x4jHtpJCynFlSaiRRKojEOjVTDpfngJ3rDQ9LJMjNgb2+pUC2voUCibqJXy2Z6tZio/dvAErb
N2cMEgzpVSne/GCe0J93vDssczt63CV4fUMNSZIvXHdpMY4QEz/W5fwd4XT+/MvJLLArF1O5tOlk
gJJnR8YKSDFINiMcohXSIYd8ijG+GHhYGrRDpcY+hpbKkiedsDev218PIkBHziEs0agUax6c9Aaw
eecIP+pxb1HniQlHP/fpHjkWXACUFQs/el5T0FSjjlp261obOuploSyB4nFUdrYsUhYKY+lfxgGF
yWiV6R7P08N6gKnJ2Er20D6NB/LD/cDvZSU5z0KypS04fXWQDeygQHAXaep1lmPJEjrpTCaFJ7MD
XVfMtl1qiAlUGY/BYsiRAZzGOTjIxzM3VyUmcPeITB/MQrc3F+cw5JrcWNhdkm06UcwejEv1jRK3
5Jfc5kOstV9RIQX8ILKVI7Jg63Vfv/SMFv+Z5iMK5mblYphqfziqz+MXWgbLRMgFhEPwI1akWZcF
gPH1uocUIXANpIONnIzqVTIqfyhxKnb8tkv8ZSMGhlwRZbwu9rVLxFd1qCu9Q3GEwmWJ9idHrVce
NbcTEDg7whAf2s1wXS5cFHLARPvrpj0VabBSzt9a1a97NQv3Bglpi+00J3Ehk4Zz+YZUWmRh0i+c
1fjRuoa+KoZV3gu4x7b1pjnYefX0yLn+Ikv9Hy15/N6wTKDA7OCSCRh7XYmDisi0L9VcRluuEUeY
HyV3Vz3jmoHcHfbjRxydu4edYBjsLVdFEP1fe5NKtncYQCxIbF9NZ7kOmbQHKxo0YpTjVykrotGA
HXfkP923ZiERbNgMg1LbVwAUi0kHaNHK/8Da6rwr4GuzFmA0q9rBFkiBsdVDsZQkdb1sOfSGwtPa
lwj4h6Jr6LL++16n2BokZqfRhbpD+Wrto/A+mCSuZVLEnmQ1e07y+nK4MZ/RoFpG5eOW5Yq37u0L
CTLGvSBwCPo8eeub3lVh+i8M3piVVUuCfTk6ymN1f1hHkn0FKqq51SS/o8pNjonoZyX1Adc9c0sr
lER8lg6e6jiyu+cDcRKt5Fox1JxaOM2bk6xP5xUad5ojN9Y2lrUuzo8ex2/KEceBMkosz4TcRjrP
dhI0XUGPeZ9rbIZgmLbhaW0QymJkjBrpGbRJfiEo2dxwD14GqZ6vQsTtNQw5xwInR3ckcpZlpmeH
A6KL8xDpJjBNoYpZ7UuqmnIHZ9t6sYcVjbsGTsWVcOoGY2YmKS2DA0jsPlH5CtpKcJpwHfwZR+gB
JbbQCHnA+YLJ6O2Zi1aGfySK3kUv+OB9BiKP4oMssqtWWmkfy3QF74PeW7X8urRX0cSa6weX7kCk
qMMiJemRThMs3gaQcHRXtmaUx0sTIPMPm/8LdtQt5gTuW91kYgCBuM59jTqfUftNUwaA/qLfL/Pf
zHBK7U6KxtsEGEpL0j49OWEydFylGXMQOuD9poq7/3X7aYrnx5VpSifhXQkH0+RaOUYjsiNRGRio
zYwv8IuXYLJo3Nn6/LBg104jOn6t2E+bhLTvlE+0CBuL86W+HhsXmwCtJACpQLR7GiZmwb7NVa7n
sZleMIPoWgkaoxLVhksaXa7xLsRa4B4IH07O86i/8MNuqcLGxwFACNWgXPuplNvheJSPYvsB1Wud
LaWurNf6gKo64JTSPklF3I0x0QysHo3qeGQpzVGc/Ji6TGclNLcUPn4pFlxFjUZr6pFBZCtOObGf
Z5Phpl0zSZ8A8Plb7rePYtXhOtpoalgEAONPQaAJ4tXDXB/hCufNUgtTlD1G6Z6ZBNkhdScW758v
owpQQ8uBjtYcJrZ3jUUtslxNgTcTj+gl98ccq9wwh1oMdHgI6WAQjHXAEkD5bk/bFBE8RrT5F33O
F7t+EtJOGege7oFTGWn7JsqynbTw/w10YXVugq8TKNs/2rrqCRSb94D08iB16XLw6jvEc63t7EnN
VCBjGA0LcxYYOjrDWz2Gq/Nhz/Dw7YRQeP2oPqp4hd8F9weP8LmvCeB2jEDD1W3FbCma+JJbSgod
byDzhMLesbxetNqaa620ZwgnB3E3k9AFYYttlXborwctw7jSZYT4/Hne0o/TpQsyE6DIJml5OCpL
FJybl5HII4MC25kDtFW7HULpK4CNwpFZjClkjkaN1cB9W7SPxwd9yGh/sJ9Mkri15Hsyuo/SL61b
ARX1N1mI0tlZDPc62EBi+HyeQt5QgqteIojAfjmiVcAEa7e5ibARelSDq2S3I9XFw9muPxmWxL0j
l2tMcNr2auitd2SaH6CLbzDbgQ469Io6B5RGVa1rI/uTxzTXlK2dqyhlaQg5Glk3xYWeyf/iU33Z
KiQY3Dwjny8u3jm7JRdX0ADWsKGAahbn7PaU10R+wQJLBdZ/dfAsR8VuaHbcHcG/4qO3a8SJ9f6a
PZYLTzraa9HUES8Gi62VBhQC8UYBiPzeTciVqjuOs2P9x/hol7NsOdojYUNaooTOzI/9cOC6CDJz
I3XaWzkHLs7tvz2OLACGHkIhuDNEdLq9TGzcGCFaKFoPcrMhKGWMn2eUMXTMzCTk5FUHDlwNK1ac
vbUzg9dDlG+ehC5N8UdTCTXM+Tz6YFmZDjXPlr7nMJ8HQUGNq1MR/3fUsLyY+KyLvCPkp//Jyu68
Sbv0RhZBBo7Wt0SYwdp6TrSQDJqFaQrVaoUFwHuzs+7jlhxsGIyLeGavxXsr+cSF5TFTAy2WhJJN
5bMThjxzeMYU+VSp1fY46Mvh0B2dPXMwJUjYZAEk97j60rG8FnatIBVraQciKEU/fbb7Bq3k9R2U
smciUKzcDChsoPJxNREwazuxY31i6g/YRMFOR3kBwAw2BBMLRP7ZGCVD/EaYEiG+ho/35L3GH61h
vwrKZyr/BQTie+zX0rye1huF+026HyKoatJdP6bj4XPLvQ3USKhDGg83slIjnhHO2NxppMZFtG2h
sN9TlwRPLNAr4yzPxYtdYXs16eWFf1DcVzQMXgUt1fNp7HuysASrsm6baZubZ8yE3DDJrRkV62AU
HRZupR9iMuVcCLCt6wJueyxRKr0HlNyzGaEstJLHiI+F5jmd0Cf1YhpPpt6q02IQ5BWu4JV+m1kn
oxHoqQdyxJ+aoPi1uwyQhygzxRq4/UVaaNTQWzfoo0wa6TtT+3MhGQVyers4u0uJ1pNJzZ5BGGBV
fWHHemx0diVdkecV45ukA33/JsLeRkLvtcMC079a0zsiQKSEET+ZRo1HqFpIXaJPzWj6lhfHKFRn
bJwS7F+oMpy/Xx+dDFuEB2YYIsQIaOIwnbW/tyZWt6vl94eX1HqkJ3I/K8BnYb80EgR/oCRHbYh+
6VOizOd1tSAL2XOf6NIBNt/m5fLkIOhN91Y5KJm/4beYZBhoXe1rH1X1o0VxEu9F8jzqFe99XdDY
NasGWDcCfobL6Et5oQUJiPB8IEvcOpcYCfv02eF2wc6qoTzVzHjSiUnV6VeKA8QgAd22706O5igp
AEGD59h1LNSmO9HkZuJt5q+4CNQ5pQjk7Q0iapEwcEE6Wtv9OTYz6HoOWxSJVUFo3/5xoBC9rWI9
djzlQfi6drLpyWf35qbwWtVRpT1g8VCGfk+cX2TiFZvNnJ8Y4XVP7mpDKb4LcEGyg9oJicIx/bj4
43eRF68cD0br9GQ7z4FzXg8V3Ox7Gve9FnwheoCerqKKbhhZGyCznUE5/A+ip6l8fnxTilJfvMvX
PzD/VskJjQQcbv2w1+2+5TN47nYNr2oKX92yF6uiq0q3qYmZzaVYKz0x6QDTpc2YS9J97uZ+JrMC
FKAWY0Or8QKLhFtiDz/84i5gsSAreIxkG2zt/Jeo7Urmv9bJhjBbt0k9qaHO7eTo40cOPp0lUt+V
/jvIkAZrKCKC1sgd9BsAAKFjebVCCuSC9kqob/JNp4qXhSC+67AQVUkJPhwTNdOxZECSzT3nd5MZ
RtRtYNUt5b3wfNlqe4Q6GLwC9eFHDXW9cbI8HYZj6DL9BBMeAsCZuMN1JutP9WqyMytW/BuAg7Xo
4YdrhEJT+zCe/oEXs8ylICFBcYouoYbB0nruTDgos+EjvBTY0Bep62E5SH8TeLqzrPckO+Skx3pa
JFKsLtvARmL9V5s7yfLGGdpN/w6Uwo6EIRRBe1dSqGnYuRMCA5CrHvWxqEDRbuBx/VrAIKhpqDW6
EHciJOC5UwNQW+t10vAkac39o1V1OBmOYqZaKr0s+cIRQIr0cdVMWurNpuhNGoZWxdpgD0rpHt4k
TW9q479qUoVXSu5YaLm1F1wWTgB1JK4NT8dDXcXEaabSkFW+yikS4cxbzRW8riW8zSB8wDHQOIdD
sbUEDww8ueb2k/Cxddbal/yYhCXU+nruBB33/DNCnV3cMQK/nLA4AEJS6ZY6MOW5VQlMhYEXP+Wa
xScouEX13KAtPXWsLv5Dn8NUGTPWf+cAqTRRHR3O6lnuRrOJbTmVjcyBjWWO/jLGf+ZDcZ5HBvYa
3CJmgQ3sRuDO8LLTROPQlOR/7ZbtIUi6s50SxNm7a5vP4+r+jCovpa8rK2kmYjCmFR5JfYbDhuMQ
U30xZIstWtAaZmA6MZMfEvaadUGtVPnKAMYq9TtlIIZZFznZTujHPnoTdhw0gTHBnFIPzsLPje+Q
3TDKMEfMzNVJylROmvFO7E65S9DXSVx5KjsM8S1PfNNu2Apg1eP7UsVXBpMIS8F5llBdJnOIGm8n
7XDH3cosYtPjIo3u6PjVPUYq5vCJakDameAmVUkS2Il9I40NcugC+OAUpxw8m28EkBjmla0BneOx
3HWSOLW3Z60Kr2mQE4KzotRak3C1EFitHtKMAnW8FOzGPWSLg1x5nETUTmD0S16sW913yZV3S8+N
1uj0FRzTlVryyqEWGpNq5V6SQK+OH5h1ubc4cqdZxc/x8wHsoSY3AZ0LqeYm5PVlogt/WAaaxmIQ
VlpplkWWzOx+kNuspPi6bboNFW5LUPEOerpH+x394xmJXRUh/IJH7Ia398zNOMn049gIBU9RsnmN
98jvtvuVeSL8SmUxSixPCK7j0gBys/8LittdU4ka6isVscFU8EO/aTo8H55KSSScMoexpaX5wKgp
5E+qi056mMdUBp/Gy1XcWC6PwTmod4+JPC3cwFuA5TCqunfbCUNSjLbS+Zg5XN4Vlb6sLApXAISP
UPAY/paBtxEJ7OqvaOkVPoOKaYpU9sJfdCjwN5GZZTNY8mfJfmuMux0t9I47jYVObF2RwZqPVXH5
nKIXGehzk9/NdgS1BElLBLRJ70yB3/DZsKAhm99FWfUa9aznJAC9daQ4TPZrI4G70eNgdl5HYpRh
3V872P2CiZLgjQ9L29SfAwtu7Z7d++5H9yqgwOk6xFvwByQ6F/NwTIEzB+j1goPAa03L680Dadmz
l3MUtoOjXEfeSMxhe1EW7E2zGGcVEvEdkRn7yf2HiJe7qdiCN8igUXLY9pEwseH4Exy6PMYq2Slx
6Ya/Sr6O29zptV3GU+aJt7rMd/LgdVhGVBTXV5fuU5oLj5GGs6GzMKrwgv9/tQhR1Cl/ndw492K5
LCvQ/CldDgJjwpXQa9K4aNq5/uFT+mdWooUSxNZZ1bI0NagfdzlfDglrC9kUUO8lvrAnwkcKAkne
IDrvTV39xMD/WK5ivuBpn5vtgiHSqB7ifk5NRbVuLiA/eLOx+k2hXNz8VXsASKr7ip6VlbvVAnDP
f4fCyPakfL0Jbat94od7N2a4ROIjrpCzMv2glGt3cMB3U2VHRHcYlCS7eojXaANz+yhK41uzG14U
X4jJdWytmj5VavzayNB1BvO0jkMxuvEXR3+Ikbhi0taPBVEMru0/LPVddexsJBKWbscpBaSLVgtR
HtWMw8mmPVQ8doMYE6TccyueyAkI6MMKvgmcHs+xVASJxUoUaNEJ6KVPQ43TUbdu8cHE3NlZISUu
i95KY1KyuxdUjmHvNeUbcQHFYprpgFnlCTkAjEs9uWlqZol8Ur9JSlawqGD/FFqsWt1sGyVKWIlq
R0wZAjdaWGvqr2NXz6w08bh3z3qsmbtQ/970+de/ckLYom/AmXJ6qLjBSqFUF1qf8YadkfEKhdmG
7XowYUk/taOrkpI5k/3mUFgriMNHYUduEC8wRtZ9Re79wSD60uw+TpPMFVBsGIP0TTx68XdMTdzk
eYRyTBKspCix1YICD7Pwi3e0Z3u0e73wAMO46bTH545TNDSzCMwUx3jIDtLrV/xb/wdgyp6JLBB+
6KlY8VirOR+hDuWiBsS972Fbs+71JWedBlkKE6AoLStj3ekkv1SdWZ3WY+5oWclmYrqPoOseSdSw
ztHwmYTMF2sIeYYguzyZp8NiUktZukJd07X/BFT7Jb3jhhn+pbZQVchbgDvz6zaL2XhZ45zlHOxl
gJ4LGKFrdqODwYHjylnbuddwhh1Qf10vijO9ZRTEEPzZs7dbB0GMEizkJejmB0l+GS5Nm2TYuwfL
kR7I/S8JDkW6g/ZPGEBXchN7CeGDjEm7U3N9qquaXgQnJA0XMfMae2zPveUoAolVjC2/NBt7VgJg
5O/gP8zwss3rozbeW7osEnJIdtt1gHu1aCCBjiblq+g5b6bKOKW/q5V+FLngGWVvraJMiWteDkru
zx+Bsz3rGV7IvLTw6SYGaAGTHClQC5Bd8v2dfCpwwhUwXiDQ4b55YC3xoSJRYmOEeNdZL/mDHpRE
imnVOJKUUArWqIzB9vwV2BF5fuLhwvIkON91usaCkkpfj+YO87UJGjpsEFfd47d3RRYNX78iSXDu
upIU9y8bVF8DDVPGq1X6WQqKTyFjRUBa09BsSsJ9Bef0V1KL5489CDZ7PfFvfr3/U7Wx4DM3ggZ6
Ctlw548jY1FH7Qe0y7uJlP+mHmqzscL5jeNNnCN4FQHIqMFJ6eUHENn3PnNLSrE4E/1bWPQKMFss
TIgrXFN3Y0lAQ6suVo/CLIiRQ6qtw12RJOcAqvi9EH+XcWbCIqtbtU5/c3KCw5/gGTwHaNa2tuwQ
95aH6L+TEbWxCS8J4ePAx7jkwg/l68ltFj94amkzuNlMl+Ceq2AL1mmcY01qeG/AH18AGi9V1DlS
qIHRZxqeI+2GpcxnKSlELc26LIC3GYw8iZDaU9CMeinc5qwAt3On2ONcJ5QZelJ7nJjG8uCellck
sAblKNAHn7B9dQihL7/y5Y5fC1gEbgEqYc2kA9BCquDK+Nu3JyuQQcxReVL7Ky4QgR1IU1ZkGBkV
6FZ00rhSSZQAYVWUgEbKYG0ZLW0vp/W5K7wUOFat5HfdUxwEf4nnsCfoC5r+pVE/EKamQZmz1X9x
42m0LSzkshfP+2FctzxohLa4iul89R9vgw6iyRij7aNK4ibLVGuaa3Ejhb6Yfs3lPLlnULGqjiqI
es0KmFEeFvro3MV1RWbQlaIpUVogH9kr3D9TeiXHVsPpLtrMCkCMXtvkLKvdQlEYkCNrYUVPY3fJ
1InIWG+8AI9D7/6ynRkyZSDVIv9Nzba7YhJO75mYHFkhjEPCff3IyHfZQLCBmtVHP+6eufGzgl/i
4D3ZnPXcUvjdN72iaxvO8jKVTFeJbc222icU0iqflB/tjSA6Z9abn34UEiAzdwYQU99vlg517RDG
R+PEoXssfjQyS6aH3NFSqOlrlOAFwjwf6hzeoIe0iuUgSzpYEBsFRe0ORjuiP0ImJ+P6hyVAMYwt
52Bg0SQGuRQXi3yqtvgxPFleE+uR/2OdA8OLwyUJiQdooONkFVGMv2FoVIX6f1oYkB+JOnRkO/0u
Sj084tW79rSgFE6weOHMmGZXFmpIGO6M7grWYOPuVbK0h2a5X2U/sKzP7XhhZoniMI6tL9itLvj2
oXnJJqYaTjw6AiMYOP80BiuObo3z77UBi9hdLEGay8Pgp3WM9386bZG62N4Yao7h2XKoZI8a0rR2
ZvBySPn96zcRuCakv56DPvhTOPfn9ARMGgx63lTt14e+bTdACWufvobKNmCRKF2toD5lOQ9qJr1L
Fg23jfMsKJJELYUTmL9DUI/04XIk9w2rZ7v5UcylivGMww8Mfwcq6Zo9mIm+On/c5IU6CmaubevI
mCL1BA6TOPXOiLTqpqbwAj+yaYNKERlOG0XsKWyG3fQRmYg+cMQUFeQ9DepbyP6kjalWGpXYZy3S
qOuJiCdDLKRPWaPvMGCVAvpVFQYSf3MeI8SQcIKgScYSOrZMRZ60a5Pd59Pv3gP9OLcqjr1sBt4+
0yiLe/2BioI+c9AcSpq6daNMTKXIWWpBtZXNpsz0ORNz3G6yDVhiqXKguXaXUcMGZUTuoXJxxGJE
TWPBUVqhNBZwlj2aGym3mF1BMHMV+mC5owT4FwalwwaLmdtqceq8XaT+0dXW59b3RdG8h/NhPA3m
uwbe1CGDT9Lf82nOZXMosTxVKGnq4FGn4hio4NtbCodOb6M3Ce3PYiZWhCD884YBb9WxTNWENS7t
1nuhEfsCPojsCgrSg8tEF8nqWUpHA2OnRP1+7DVS4+h3nRYBIMYsEo5N8aQhWZlHikBQlYmbeUwF
A2bvt29fCCuC0YN9Od3nFKGrhAxGzowEvB2NVGIx+CL0TWOkgTxA3daGZew7Y+h5vJFf/MKcS9/h
PK/v4x1OusSMtLsqa7OzR1WcrlNc8IZyBQbcCer7kKxWFMG+38o4e9x+/E9hWnestDeovYRBIexT
M4jkA2GsRB3DJfq3LVNneIx7bfLl4eFjAKqz8uM3zccOjmm3P33dzLYywoRJULXLs7IHXMCy7ibi
puQojQC0JV5rgauGGBFsqS9fmQeeChsIprSyN9m9MhAbLPQQ47D5AD/dgOb5PArZZC+6OB1y6G49
wi4D6IdZVGGe2YGno+9AzMMFCljPXJSlmQN/nWcsN76TM8yD+2e6QUE5TAYihZNA7af+8jq2LBMo
GJWzzzI6xkKDRI5HKmad8fbdu8F0DIxYaABIGWhS10rd+WxLWe5XglX3s2QuaBJS62OwZ9AvXlQ2
NjdFwEm5BmHrosuoyGBoH+mbj3K5b63G7sH8FYH2CG3e7XW0ta6hyhyVfGz6gnRPZwv0eH7uiQd+
05gnSViayG5w4H2fEBtTlN9mpNpVXrYgB0PnlTtpAm9fldlyx1byG0O48iw6ngkC36NB9BQ8SZ9O
D5ig+FnIBVURIfHuvPaG7wb6Q52SArn2PTo67dXOkLm6e6z8W5/Pd4bnG8d+/19hxELOtgvkiKj1
6QZktJ9P7EsttVMWHnDaA3+77ioDt3v4Psb9n1Hfd/Y66y7AGa651x3ZfOVWX4ca1e6FW6KcGeXb
piuQn8jo1Ny1n6bAMxc3eOwIXKCbAwRnVUtLqsbJeKqcE/MpqcmSS9ml0fq6mxc5TF0ZhE5nV+lj
6ZYPK5L0ZiigY2od1fGIGVnXQg8MfqBFjDZexDTGhzxYMTUvBl4w+xTUEbIDQfN7/dnRP9VmvJ1u
VfHGM4uw/+wxdVelZV2w0kpEb6jZBTsaQopLGCwkGa09fyS7+vKU7Yg9fcUCxKhMw9o5ha5IrKLZ
k0yLa21krJt7JlLQfBWSvTmT5FCxMBR9hYO1CTGxgE2rg7Czc7IpjBd4KbzfA+0JC1RwmSHhtsus
mO6DVqwxW6e33bEmeZJ7FJXOVkoW9RzGC+OK66xtH/NCpooySgdKp5UUDCVBih0AzUgTsUdbTSZT
ljy4DZrKTR2DVQ1nPN1ueIoprbHVHFK/WLWk7cI8QiZblz+5yYkwpRQ1TECnjM4Ztm68gA7mvyUc
HM66dBhNn8wORk29hQu5ga06ldJgzJJ/6B3IZZ0Ol/uEWthlTAlnfBG2vpS1/RQuSBlQTIsuruKM
6CC2yuYZmaqK2zHj2uZQNryOB7JRQLCpKbPUX1VMuaVM47Tj086nWoWPjoZ9PaL6JaYP7TgglBYt
HBmKgmMWfW+whl5eEZ914WhjAt4Kx7eSp5OZDPVIXdVLv6R2wgIOpWtOszvyQwWYuiz+J6GgTzOs
ovgPCUxFwfWC5GvU3rB+AroVrmDpe+yLtNBPXepoFWcmzrQ20tjB28FIita6kkkwFYCeigbIiWyO
i3a6wOvztRGYREbbVl8m2tjMWM78Z6Dg7vvv3IQdriiy0Ch2kBmF+B0uTy3/yO7ryAr+q8QfknqV
r1ZMB7O4K8fxG7VPY9vf7W/H/VYMzimo0ZctdlXuJmvT5dsfBrV4AYLGPYchvAOrrYAebVAwQ1T1
T1+HJdzi0vebgSmzzZN1Zsk4KBy+tfA6nNYnuHSKjirq1BWcJF3Sno+soS2kFtGEWeH0J2jxzp7Y
HQs8fchjnHnshG9Ud50dy/AY6CQFpNSM7liFmcWYWiEWp95FPyUhDeN5QhJJIaWYaw4rg5RH2wJF
q4/2rrIRKqlIetcdj7D9KoV/I9RbsS9BWhHnylBaxZzi61+P8A9vNMgrRk4NInctKD0FCNA5uiBf
MeCtpFM44Mpfd4XrA63qNaS4asa7uba1ucKmDQDHwJwH6v3DOloWaHiEbXbULDOWbPEVQCYH3o5r
vIGGNpMN8AtNUrN/5uXCOFdWUBzaN2H3KM+zeXCYBMqfNjPzDxBhBNRfwIG2qhFqHqVbcQX6+GUq
7qUvARuO7dTGviAxP2fcayHQD0QwN69419MhKSwLD4XOAfS5ZxLejPVfgW54dtFvRGlCEVdS30Q+
sa3BGmFSNfyMh8pQNJCREHEkwDH40YB38EOYXDv+p2oXg5LidePL0gSSMWvlW2ACPP9X9WNm6/VR
jlsYNzQmKijhkbupcRa3qAuCxGmwqxKvBgpwwutdcEhG3k6IwDx7jH5IYyCyWNNFW+031VVsQDz4
FhcAlkViLqucrhLqkIUeXe+JXPLzOd1l8eLztXqdk/OoNdUEab5NIw02imwfvTaehm3Ti1WDrmrH
8EBMt5Xa9eeXPO87BC/EN7V2Rsz8+tBoe55q9i+zKy9aRZRbLR7uYADm4JV6JQjomLfPN+MBh5Kb
wWJ+gA/uF1DmPEH23Jo4qiSCnk7P1Fz7DrEvYNmyf8MD3MK1wvKBF4pKlwgF9eiNYEC8CK+35Xpc
eUvooz6j9fdGhcthvPYohQiJj4GRihDAsKBfBvIw5texOxPdRk1fxW4Ie3Pik4Yd1EdqiiRvviKl
J/HPLJfMF92+iRgsZE/9RF3HKcwtfGKXIhAZn0ZY1zQP37V6PlqoEHdxCnQGPoqNUyEBZYxwqO8c
faMBLGHpgNAs80pvD2yJ0wwXSxj5yR8nditu5xc85TztJ5yzN4JqVAGw9rDyWQ+xKmfh7s9KZAVK
7RqwfN1b36G6oqxeEhD+rSVxgE8/J7vO83VdN/YVDRMM+UYvEPxBJChXAuIP+VcIScMuR5qR5aT6
7E0TyO9B84ckIn2emuIXnAYk/6gJg9TB6UmUjz6lzJh+soTEGZ0Glp/31UGME5un8xd1RHrwj5xH
adWd7hIdI2S70sjyr1wV1DcoRBq9wPP30YsX408RTOB6kvDvhKrreQHBCFmK+u7CoVKrGhBOHG4Y
UqzS9vxuu3RYYoWZGMfpSvEuqC+SjOxEGzYN9CplngJyC8UWlw6kQdwOMtEMJkJG1W6uIQgPxAZF
hCTpP/J6Ae/Q/Icavc/WjCoKdjMBmnobQ/wMGq6SrToTulx0n0Vvm0qC0S2d5xkOavGAG8Ax/okD
nT3j4WQzPx08y+rXQUCtkgzlpbO78WJ77SGafL/3NGnJjnVf0BLzzI/a+S3eVAomh348E6Hp+iPC
W+5c/0zxYrbv9EUM7uuPd0ZilzODCaNv67QBfARu0UPdh/BTPR4gnH7yWScWmL0y5gk7BST78N2x
LxsR2xmyVsiT9zP1P0xV8wdOEbU/f5n9lJqFacf3+PQkgZuvUNou2JMKlcrfXivRi1ZjA0mk9VfN
MVQjkJeqMJLLSzOt6+oA8Ph4YX8j5Oo6TcG61PigIRTFnJYOfYRrL/hGsox6BqUj+hGvFlJlLvC8
eEj1IuyI7/5rer6zHIKO77oKTyHdtv42VKCslkfajNbyV8lqP0jB7Vq7ma6j9mTt+Lf9FeZxWRCV
89ks7CSiVcDelypBBpEY5y3CuKo/gKr/REsIGyrFZvv5D4t73aAUeHwaEt8Uw6cFZ7j2JT7WDoQ0
EQekhwJNJ8LJeO4r3dn3pIhoPKBKsWTvhsM1y+UjsuAlzMJL7nUlW62HHKVi0D8iDFdqG2US6/+y
7FTlFGjdMbSV3OxP62Ma1mF5fyGobH3Zb5eA3kiy3+gOnFJg9wxfMaaStdmrom2MkHViOTLYlgxT
n3PEiUfeKJ+IRQaDCvX51MZnwfSk/6gsM0Djfx6lFgMgDMw+LrHo8SgkHkKpOQ4OnBQy6B7tSouO
eNKDqEU/41bwwZ5GqTzu25psqQHdYoyH5R8tTqOA5nFm3lq3FPFnAKua/HK1gVcRGSmOlaI/gR2A
j5nS/coSJH2R4Dxa27EkCDjh4oWSq8PSegx2IdLxhEYOLvq+ZIUlB4WoQ1M94mI+LkBgAaJe1dKw
o6NSBgzoEI4jsEU4l18qQViGO/MSiVEMUM8bkQodoxE/HR8kjb+sKSw2el7shRd09zE2k+1V/WCm
BpLOUPnKw2oiEOYiOpUfNrM1A4x1r7TlwA0g+J2Q0sw3JkvnzgsViTtnIbyXpzpaRa/rQnWO0CCs
U3zfbyfpKbanuVaOD6powTXy8z+hoKefvx0ObKokeXw9IcspbzWb+8f8uo7eFJsUh3R5kXGozM2O
lO39V8nITJZLyJALnbd1eIEJWuMMZ3vgvgX7QAAgPsJwC3J5uJZ4TqPBApNqt1PTLkngPXqcTyU+
7nB2adXOnd98+hxCE0KGLl0lElRr9CrQsGbiVh3cNYs44uUgnM1sr96mAXAYHi/gTIfvVVyZnHt8
OuI0qzBjjkskJ6YrcEzxcqRsDGHyhX3NRzdF/rNU0htoOokeYzQFsnBzXHvwO0asa8Vk92diUp6p
hxSoFqPHKS0aTKSUwMgH98/XNMVlgTTeFRjW9VEEzfB9z2UvhcVl6UL3uWEC7TA2dD3jswgE40xR
oxoUchV/BTvCBtzyW4bumUBK4GHjCi+AHffmwssNIW8Yy7BDiKLuMVVRftV1UL7GYHEtZT2z+1ms
uah5GztoszLwiWl8EVAw0tn2xGdePxeEUYjwqTSpzyZu4anZzVo+yeSNCrSs+BVXXqi+/icyg9DD
pG0QjJmbe113A1y7HQxOLGHF6YNy2nz0Q6O7t+J8sDJ58vAgeXjR6mFlTplE4O199T2Db6QIAQ+m
I96XFsQ/MvjEc8JUuWxXI7NaEq0mYsAtjxGv7aRSkqc+SyWm+MUpIwmHywRD03h7YsQDzyv1hI6Y
I3As7HpGzJCDXzbF8PpkNPoYJQBNqwqYrG2Hm0MC+3DOBMwmcvuSHTKMTHSMpdFPUmxgZ9sNlGbW
Q4Ob7ahXzRVs0SHyPWdJhO3ghqsB3fhKi4y6SwEjDlycT5qSOFmaT4zPNsbEOV2ryq6rA6rYpiBX
t0zMlyo5why+MzahZL21gxXCMCX4ndiT95+Cm6geyxmisXg3rDOBBy/GisQzjO1PDUaMtiMiGRhu
XHfV471PTAjBok0hgROZCwJpxExG910u0D+jO8+CWYlxsV0C4oB4e74wPhWXLOpbCrXfJJHwSKaL
8FAG8C1IfJ57wS3EFLkvbygEz4CKs55GT1yLROKZEa/lsRtcy4UFwbciy+CV0e5qwR1zKrUdRocA
Lg4fWx8c4gh5FBg3DAiaGLrPUCWZq3Qwwv6l8f223cTNWoQ1C1O9e+KztO+YCCXH8BGhY4DEEdMU
uQGXSZewPceLoOcLLj7ktTI9OZ39NHXZE3UdHLfwMccSh84Sgf8VEPCHK+FzezflDjxie1S1gOSE
MiYLYN4fVVyapLAC1OG3y0WUSQDw6WzN4ET4V9WnhIamu7UlDln9wAuiak1fWpJKNmTDnim3QYlz
oyCqvE9dwEnYkjERL4eEehxy9wuNIBwefaARIWnHP/QApWxhJt0LMfZTCL3nlryvy/hjLsGTSYl0
sOcrercfkafk7hllypSBPAiwnKewoPQ5EQ4HWCjT+rOcR0cromM76ma/NkBsiX2eEyZrnTuFFHnP
tEP/MGjd4H4sVUTtIXIdgg8uSnieY/NUzL3YCGtJGb6NHuzGSXHZMONldx5OxDfIA/ZK0dEWBm2c
/HlqfDJK0DNi/16u2pkbo/WpapzjNbYPhjm3wfmNfGq3mAY3EHaCFwsihUuoKuJi9q8zPJS9ru4I
vbPZXy5ze3F3W5O6SPwE6Bta0zOYn/0v8ZKwcU7siQirhZwS8m3gupiMAWMfb7q4sI5ClynVv4sg
3aqoARfQofoCRWr/9mGumMpKze2ZD9MkhlRl+cX+y3mnUvdAp/7VeEwWZOsNw119b1ofr1Fr4vD8
eAmGvImuLb/54N5CbC/wnYQUBk4mWAjSxLI9jMn0ZOKqgyNiOEfqqKGW2UuO+JuN37amOqt8bDVY
DzchEyxvcStFVrcBvSsaEm3EDjwSK2a0Ig+2uQjL2vS/5YNnPEJ1qrk672wy6rzNGxV1luePAmr6
wL/WLJ4AfarsrtNYbz359K/9YhHO6C5EBAdeTPqFYUYDO1ts8Dlckq6Yu3Ci4FKm/Y9jlTYiCfBG
vmJoQ179/TA2At4FcqCAZ8GzKP327ztOTBe5auFdg7YBNQEsVQVhZGFsHGt/GOa484z4etRNH3Ps
KsWvxXt/RYTg9Wwe2/XbUgRK8J4St3JtanvnLdcnnrRzfC/6M7/qgDA6nrLtWoQcgjV9j46jiMF/
n7m4eYNj8Ym+RbpH7BAKV9mKpB76kiVDcD7K88ow/wfOuh5g9Ft8bRkVoDHsF9bd+eWKXR8/WZ7h
gMMGgKNeQ0dfxEDwUGTWZVBTje2rXU5MM2GhJfFhkPNwaoXshYKOSeQA7PxjkPpAox05K2+46GQD
qGP9ZoAvlsB5MMkfIq2nWozAjTqCzUj8MW5qOIc037ky4uqhdTqqeTKsmS0I8APZbI5vwKKj9bXu
YVNppyv0W+3dCl9bp0/beNtr+JRL2ZCGvnxXjM87bLpRFh2BJWuoB3WXOmuQvsCBZT6sIWRR6Mva
7OAMQuIQVBa3Fa3+2HZZmDqx3Sv8hHntWg/zX81ixT3e4Pfm3tckg1rSAwTMyFsTT1A1qZqpKO4E
oTtAv6LMZGytBuZ/IGxd8FQml34c64qetXrV9qgWfwp5XmXWqh1jUtUXMHTHPiyJ+0bWinqFYJRq
Nizt6GoeFoiJh/auXyqAdrEQCkT6eN+AFrWFBl2z165o3YL7NwnI0LyxedSEe/Coy5MGmY9iksbr
30bAfLc+LBST2XLg3DhbA+6dGa8fNS91zbFtcJyLRey1UvK67CiADdJ30x8dzN6/qLc0BoI9Vl/U
p2dSWGRoW2LUroyCmBUNHdXx1zMzaego5KkAqcbHD5fFTPT4vc51qBAyRiCzYnjUiDiBG0OEOPjv
UT3o1l+2fleSvPUcEvklzWbeDJYYOV0j17+/NTFYc6rhsfQSUqPa0rdWkduVS87d3MErOMzslsDm
LcDrYuxUvaDYr6rdHDXR5fInwX5FeuCCcHdh9hYe2NwH6WLSP+AUuQL1zXD7m7Yrb7OpOuN1GvrX
9zeSBzTXjUjrEFpWgwSMP1LdmWyOrcxfhAd/RTCP0cIr72YbYJcdGDnpX1jhwtR4peW7W9DkmB+z
NQdc1Rp2mj/rS9Xf7RCKnpWMBLDFFeNHaHknEIkUQou5JLMxdCRvQ2p2Y0pc6O9VnGswRru6N+i2
bPC5yJ2S09MDaHZxxYUBHObZ+MI0fmjTjK8ckfEWdI41Zh3SwxOSqDmnFZZIb+aTH3eH6IyOuLlp
mqy3zM5zjUkEbpSfuLoiHn54y963QuoPKuXDo8sKnUYo+kr1EUbCcgNA+FGOSVPiMkNTqnWq469p
xxZECq3608DM1z7+IzwT/0xUHJc0d3y6tHmpeiuHTYjnaLLgrpcI5zXKKoyUNWh0Ayg7au5RLq36
zW+suk7I9FNcC1LNQ360UBhYKkGs7TTFsccVIY9mfZn7oCqGn/YzBZin4yTVdyG6IkDVguv9SCBM
9ykat3PM3Anh3tLstUGJnE6rdhUm6LIPAJlB2v+xm/ZJSn/s3aFG/2gqhPvQ6fm/Ek8g2sK9BGeA
M9HBRvbHdUIw7MkeWh4Rx3grNMqul3sWwVlLB9cmUDPY4cm+zEPKHvEKlFEa/u4uuQD2jR+n/ln3
CcLm/hncDX77LNc6xs/u2pmEvDAEMcs3dEm+GPxU4zwSIcdRX1ruGXKbKoeHrbLhhkIrVMe/at+f
mJIlicrYcMDrAw/0AGY8Oif78vAsDWnwDbKFxnHNBBOwT6l11WOLkQzwN6weMglgoXurx6lRkfl1
jRbzLdOuiOjbgImJTXwG4PwV3evJdQTM8UOX0+4x35XTh9chm+pF/XfzizeMGM5NRo4k3stBJUyi
Sg8l3vj1WxEkq9u1ZW60uv87XodLv/UKfQEjDOuTf+CsPMlFzHR+Q0K3l8NaEKyxzKTFZ6b0toP9
GLpeIncXb7NFKkjpeBSz/lxeTtPV1sSjgJO6g2CVxa/aqYaGb9Fj/yYNZiNUMQN2aOyyuui5rUo9
/YQ5NXenYjynE43W/ljzVj2aBVXTQHZ5ivdaqGEIcWauSZ8cNm7RR4vaDdv0fzwzKv28okfqHImH
QBLGN5b6PaClUIzSMKbs3x2RGF4UFcwvkckPtGv0t3e/ZWvBjpinIxxB/7LvMJqBqXMfem6WBlis
Hmwk1YED6APlNk+UJhtCAbXF/BLz07cdKy9O5bsYhGmgfsa0MoIGucTRT8/zWWFEZ/hCURKe0k2s
6LgR1DqTjeUYb27YTzEYExtMPlKm6AC9suXRoI5H2G0I1VihWUjtnCt+2Z7tvd/27HFoy4VxfYG0
kZw78/qc2NlPd2PsKU8QnXdvmgjVtChxqAt/d7x/pWNZYLbv2a0RMujuMuX3YDNi002gwcFrPdl2
Tubmz/DFV2zxozEG26MalNi7G5UknrWWYe1mpyZbUasUkQP6ETJR/yqlRZh3zDxcjWKuDaeHWSg5
WA1qDuZVMtdcIMXpcfPIOvYEmZnub00lGfH/ZffxiBcKTNS7QHuqLsCll4DcfagAEgy4QCMBh6fe
DVqneYQv3hHdhI1DUedt2vY3Qe48g+2dkjVyXV+DksXOdQJGZeqnrpMsOSOIZrK+84QcSC+cvycs
ZPjkpGuxu+Jg1G147JFQ0QbZjgFw+h6KRt3jErR1fpG9UDgOLDo+GUiLPkyWrkNxNYXWj/awW/27
FD7BLwFkrkHpDaZiuUH5/pvEPH2eXPwP+iiP9xqaqGMbe94jhKT3BX07UD1uj8GY94v9mRzzJO0P
LqPobBN0CXX+1DMJiVLOVAqD9u2gQZyNr+B6L7lJYwPJFVkwOW44jKCU9P6rjpP6pLjPk8L0bbid
ig8nqWIFVmG2jHPJtf2myMQqPL9du3kdE7vwVci1xhQgFyaPiaNw9EA6Xtlf5HcIxVtfrl8pCkho
TZq6fzNmK3HGOd3KRW/hIAhph88JBVuTeyLiR/MjJ6Xb+Rb8fx5RSCYRD1be+dYl06YbFvV5cr77
27QJN+aQO/rEan2cV+MqkKjpZsXhucp4mMgUJhDSViQ5axb1krKNQqzHf/jX3k8KKu/TRXpzJ3ca
JVayDRSHptgcw6kNG1DZJhMwpprJMx52QtGYqA9HadehCBtZT9G56Rbzx9dM5vB5vwmiZeful1fl
jLcaiFNZSQnFBqSXh6YEGJ89FBFMMPRJgtjTmkl3xSghuCSRyhhGYSwh5+He3d1Au4FScTrReEtX
GwQtQZtbUWdZuW7Kk8Bv2P64oIrcWpt27BzP3ImgnU0TNn0+aEEA9sxuicJG+U8UOx1i5mB7s8IU
TWJ520NCmCB7FGhTPAHNUatKXFag0PEgxPiMuGC1UFIi4oeFLHCqj3dvyir+F6JAuSVuqxLUZnhM
MK5LsEtjPBLgnBLtzZSPQkPWI0Z7PIXi4TDd64E0NrH7hVy3O8qAydj53ev8bCf61tYOs3Usawaw
mQukYUxFmNiJgiJhlK+LObFjn4UyxkuZ0yMZctoCevs4N4WL3/4LCPqT2Wch07pIC9rVo5HVXeij
aF3mGMdDFGRHOowJ1mV03nrPP6zv0ExeC04Y3YeSDYXksx91x6u3zZInVftiwwRYitree55+v6sb
PYrqLXdewe2X12jF/X/+K/SgM8FB+mJRap1WUKephq0N/34MMuTmZJOHByeeeSLjLZ0Zb/a7zJrs
5cwTvzcFUsOo6S0DaM+UNfifpCXvbTqGZ7BhJH7MSTc1clQWljM6N1Czf8YcyxC9PgmlWsmuvhw7
crUkLzuqbekdZ1z16D7K6Y7EuE3EDAcM+7l2b5uiJah7Blisail/pq8H63figk1cD5PYy5nU8xhs
eC4r12WbQrbSkg5pceSq81d5czEChPe+Zn3fCrsOaLAbdbycVT04RgO2z5kgo1RC3gTpNKMigpLR
UIKpqG5sp3yz89cf0sOxHSBP1hImoB+qddC2AIghxJsDi++/bHBu9zGoIviBsOJjDFwnaRPLa+t4
wLtVVS10K4PaSu5ZOqRmXEi2Guge7mUXHHsr6iaRI36kmAeOXIhmwNilXm3UvcwYEothvLPrGiQu
+m1lkFOQC/CajJIDuQyLrhb5Wf6WSt9tl4dmxCoXYnZ86W63OL+lSTjlVj+0kJZVMgBkyW6p1T6D
PXYR7fy5gNj+ZWY9IFlgVvxCvSxikAXPOGGchwNuZnMqyknmdblYoOS7kNifvAGz5RksLfm1Zk0u
3cs0q5MIpiF8O2PXp8//uKd7kXAvMuUGu7gEAIPumctYYosl90Qmc5HOp+535XPEBvyfnFufuD+N
YBEG9eCGs03h9X1yRyLjMsHg1jkgSUutvQ06J0FUdsTe1KheKZ4NVQvT3kgyLQUVnWdLRW52Zk8I
W3NjSA1l3Y5S3yXzHVIwuJw1xEVelxfSFpLXeJnze+sX1lWc4FvrUPB1KPc71FCrKmUDO6L4e4V0
1ai790W8J6VgSlIAejvhSmAqkPEDJJH6uW9LO7VXraJwriDDpP/ZHnkRIvCZY7vzCwk2AVFpaCBo
EzZSxfXdl0+Jk6p++ScuXLeejud42OR2WG5tizfjdOoOu0y9GsDlhKX1Udu4xD6vV4JhQ3E4BkTd
Qf/ttzcjPapolAfdNDjw6HK5oWI8sXl/sB7Na4qQSQxSeaZ4n9CW3zk0b8zEwwN7j8y2PjeJWml4
J97tOmWrbNI77LwECtSvVKIrph7PsemT14WW/Bz3hVhLBwNtM9aqd6gRhnVvIeZsvOGtZlANVHuE
fm/HGBCFt6rEdTRw/2SPVYGHKlW0DSKNU425S8u2HcynYFTwTO/qW0vAQQLKZqzJlPFNQqroVesn
+Ve6eavf3bnExmdIqOAeMzNewK035LFfmWl7IrGDMBQzESf2N1xc9i9r8QuQ716V6/tvFReZR+MI
s6ZXh36aHljEo5K9nSi6unerGXGGr9fRCyuIfafDiEDCrgqFN6gSU/0fUlbJpBoqGYY2+z5D183x
4XzWDzoNJ9BWYNGhudlnEkuY6Eeu87WSwzrgjoliNGcnXYFnqAnZj4+ZghwFMJ/h5AobOvP9WMpL
YVIQNgPHEOXvBUtZzEEMSZZrgvdIxODhrhlXW4LUdREW1fFnlQKv660vpXNKUIZRW8b4iI8zuSmz
cuHtOl5ua39Q0fA1sMPZOqUpUPEliHUmvY5sCEvtf+RXH4r1WZjoQf0Yj82D3urtaiO+ibtjJzMy
/B9QS88hOqoLswtoTyDsMZ+CXNqcKPlzBGShZY9vopVrBeYf5M2sDl8SH55Fx6t0GSorfceeQNBI
surzH6MvPzQw40snPiw+h7wHZqU2XCkXOhU3KnSkd8jNetltlmwbgKeD4SLgotZEtCDvI4Gegyxo
vcM5y0a+CIIefXz7xCB/1PXl9Y2kEZ2reuapKd6sUVT9K+SE0KCddJ+Fv9c/jxF0BOGHeJX/fVhY
uTW4cr59nAZaF+2q79T5UveTFLtQcPgrkhGIHVWSZLYDHVSwhrfJGQGY3p0r0NLzaF2rhQApak7W
cHwiRG9UjEyubsinsL6PtfKxv/wwXbtGOiX/NAJgYk0sk4zm+QbDb0EhKVhHG1QsV+htypFj+5FO
GcEJ6mtri3tXy2gqd1C03+Wr61l0j7CotLbqpWt1TCI2N5FsWqZhsQQmhxw/iUZtWr0CLg7Kph04
Ilh4cbPuG57Qj5tjXgndrei/Ksx9fGJLQ0+u2qSqKJ1OVFolteoTHAKdy8HHtsUTN/iXR1tjS0rB
/jLRuyoHaMHNrMItepoxoZ2YBR9Cg+t6slpAtbcka7S5lhOyJk2dfSGPgh9qkRyhrWszfbt4i269
7rLVRHR0uO7JFMvVM+KeiuYBzYQhZUXO1ThAdMUiGmSv5P8OegQ5LK/R+TbNpEA/Qi2LkZC4Zy8b
01ta8VcH8jVloqXPtunrVuK0ZjAHMTH9Vn88/QwpLf49O9ds4LKipL3ezEVirRD/T9RF/i+UTKFZ
jox5exBsbvr5Xu9LbYk0KsUY0DxXZuRGdAKkGQC7rmeC0/kCKtwmwrIxewdsf2Q7mRJm1xY1EEJZ
nxRL8ZWKC0T6SDvcygoFg0t+TabwukScOtZL3AAGTFT941LKzi8gwS1/t/NLzqQBsQQ+Ri7oJBWg
8Y5KJBQFkIXnI+IvZBDiwvoPDZ20n/7NnisJwXwFQ5QXzNhkyoCNKt6VXt1gKs1vuuMjRoBCDoTK
FatUcCcSiPRIQoNxPsf3h51P37iSX17QdoIS61POB4TYILTFQh3qTwDHPngXl+gTCHOghs+Hs8xI
AQTY2PsX06IWupNhnBSKsoLTL7Z/HGTmpJ+XtixQFsKyT7enF/1C6Phhlmxrh5N9sqnXV2FlmMrl
ekFYvg6zXfiD++TxWlb2Mv6VpeXOrqmbxk1f62hiiedQF28n42lkgziyA7VoJR53qt6qisUHoFQg
KMnXo9AQFDQZ0OrXNIR7snlB1TOULZY65kVQu5K7GIZOKiYmjzF8kQBkXWdk+Icb7STOpbpcc/ML
hAwpakrNh/XyFJHtNzrDmexjTqf8cToUrK0FABxP0AcG+JCb4bUo1gyxQ9wElRM1hZ9//CpmPNAn
Gy5Y3Bn7Bo2Ua8y9RUaTzwB8b05YrjNKF1vrARDjKmhX8kDaVZ05MV/1q1PIQe8rw5wB0kgYgtFR
vQGP92r/zX5+jDBLtzq+awdTgHcjd5WfzKDkO7DUu5niRLn4wnC388PHq1r2BGnNTNJmioVYCnca
N/kD7N69k5Sy9zm02e5t3sT1q18um19vdyxHyHmf51exr68X9o37yl74x9fLZvV2PFJDGvUGRTBt
vEdxarnqJaYo2Yic/o0DR6HfMSBQ/aouzsqTyM6KEQKZ8qDPHT76Yj8cxG3fjcOpwQH9G7ZFssff
mM8SIjXfAUsKqVs41RGtSpZEQG1yLnpyxkq2cHbNXuseq3oFuXj21SqmIVHZ3s3drjKb3BAABk9Z
ykx3QD7KNoSJFTWAcUTQhXx4xJw4AwBK12IqHEgAnwqfotiGgcUfnxPARxdtseYLC1jJJdJaAeJD
0v1Oqdzc3vci1EQHoCTLFtHGPoBbaiwaGKx++y/HFhhKPxeNh5Os705sufXzqpa7V9KQ1on2A9PU
t5R8a1U8MhSPptUsMQV5aqkHxjqZNnNPapRPAKeK77mAdS9xTciYer7oqhw712QehK5ts8jbi3m9
r2Rk6hSAOM34jwtycbOQL1bc1YRxlReohARbUmaDtEOrB0mpVHHrox4pDDfd9Rvgk13ZT3O81FWH
DWEY/8dwrefne3mrExx9ldnV8lbST/6XYAENhEpFgpE75nTfr3/sGDgjAMKrTWodngplDnUwGTSK
Xq8c/GmqqmYMzgmLYRf9ZPKtQhekuLj6MSPHPs0zYG1DV5JSJ62inWoRZIftM7aI2jui7J8UgsY+
cK6JwQ+hRa2PIH8aY8u7p0lO8jxW3ghKhwteegioZu7N/w3lST+O3uSdTQHnnkiDWP8v9mEU+eaR
W4sqWSrAtluycF97B/mBkFAGaGd5Ks0Rq84svxeJCZzfUpOOMp1jBioVFudPhZV0J/mclqFGiD1s
tuHFrIGSix8gS8b5AQecxYv6IojH2FyX9q5SkIo7h/xL8txlr1U9rZglPyUP42f+zBxGM5kDyaei
viYig3xyu2WN1Do4sFvS7jEmlmenhp0tFyMELqjwddjoH7nH1W4ZnuS/pK2lBcq3IvQVZPITOtAr
sfvsJHZaS1FaXV7+V+7DDsJ0QhBeUxjq4rSBUm7CwiQ3yC5N9fiy6/cXL00LjUYptfxmQPlceTl2
DpIhcdNxe0OLZ4zMfuSBiQ1lwRYmY2gCt177GwNOTxSp4jk6HkLarx2hN58pjP6rkNzZUJ/wmoCM
GPY2H+tHBgaJBsn3iTKJBPWJEfWN2ELZmhM+52mQXTDw/yYgXjViuVCTrlzleMTxKY4jYQQNEabg
rq2HsWHlXw4NOirnStz1m4GwPKgDa3NPbZ0uxLzcEfDoaRBt4tFODiKb03cYDqb1YECYmNvOdjwN
+geIaz48WdM0TxB/VFgfjry3TmHqRKjAvI2Od5Syo/Tb6yxt2/jm0BZHE+n8MaKGE23dM25Qnyg6
KmrxQl/BuifG7+D7qD9/9ejAg57k9QLWyAWSeuFxLtZcQfRI50hIhvRRiX93UUVIb6wSc74P0Q7n
arZvMlciFlukHK6bgZP6CCPk7E9GIfnD6ItFwcZ2+c8Kp8VLQ742csLUMRZ48bQydW1c2DBI8TBJ
DqNbqwCzdee2r0pjHHcjpZAO5CGKoge0XbzxxrXcvk/79jEGf6YF/gDljxSI21/pD1FRMuYJup5j
/oeEuP6mslRdk+8gKljnJJV/cKgs3a+AkyyBFzEgsgvH7irdVwnrmTnCyIsZjpWQPWL0wtVT/pPG
dOXY8UM5fdbxlqejgtSm+etul1eCCZt33dmMnv5O1wHZ2kmPvzrLBheJ0YHme+l10dSb0o6i4LhG
B+MuTzs0ZVmy06d8dQZFIzmio6h/IqYwgwfvPBHujRmcDdrkdw+C6mnPByi11CrTq740jUPwmCID
H69GlTAgvdkmASfIwNA5evxrwoxYxUIpcdrRdsIlN14zOTghytpaGr85vboxL4RwRTD4wM3fzqUb
8Y7+xmgfCXUxgF/13Zb+SRu16g0PiNg21fTTMYuTaTeP93dIqlmYiCpYMiGKfjjNCFrphqQUik70
EakTocLwRjQzIdwH0Ou2lp8LGED4kB1cF1zbC/Ag4Y4NnrHEN2bwHtXxTIY53lCw3vSI5HQ9j2QB
qLePPZMQkHWYcQQY1YT8d22dZsbH6OuYz6oqiKrYtT2UXI4qNTiE3Zl/YeYNEvNwavvsQkuGnXwZ
w9srtma0d8tQ/g+mHmwpBlhXPdBHFtKOJTSqSOGz3DjxWIAlKvUAFsXwY8P/DRcaJo6Qjq65N1vo
YTalZ7ImJ0M1xuSgp8oW1xaay7IPZtkJQGoxvC7OAfPydINTNiExeZnyaAmNcgA02q/F4i+Xojan
afv8p/slgJWJrY05HEHvkJWzV3OGpDNO8wd+craq155f4Y8uhIJ6/ju2J5okShgb9BzuQ//oCdIv
vTRNN36geKnn7SORA4cK7cDtDgYCNgEDe8g9FKcmx7PAL124O527rT/FouKaCZh9ywChd40fSXyk
UXcet/rxyVpVB39/q14Ma8B2iNtmhAHUgbFFxvnYzq5MkKCBE9vZeDwr3Pr9fs8qVnQNNGnN7eld
IPDrQqqzhbOj+8zEMAvi/ms8CDmoAiEdoZk+qaMLrPwchQqtE/bnB1PjNggeAjOt/oJaMh/iObjd
af0B0IpjD4fmSknHHcZKe99lZfVEniBIO9mq6e9TH6zZ4WOJPbJQYdl6+CyI906WFzvluRJlFS80
z6AEKJtUxMBbToAkMmo+6bLj15zHJZs5EWIEfGQCpeaj5cZcH3VRqa973xbDh9mrOHFDt/VSBVa0
gGzpnUn61lBg5gjCCBBLFlC2f+d8qbVPP8fztCJIit60Y/Oum/3LYOarbe1EqpHUgnt70UgGUFI8
Tx+l2ZXAkRO19k2d+luoKz99MSxNjWl31Lxx+VzjQGLT21logvuf1zLTWYLen6OZ6iBhm1MLWN67
JsPt6wb8vCpkhNC0I8nP6k2QWJ9YwgmoFg2UMLs+DPwmW67Sy9+Wsu1qQ+YMpjjpTtmuGoGYkkTX
Ab7gPJP/Aa6zsbqkwQusIa5qCbUYdZncl+M18HwVQd1IUgL2Zh/nu2biyavk8ZWoh2SEvbgruZQe
Qb8DES0FbPu11c/J6E/01llcI0wiPunOeIjRR7V9NcltlXyM9egaXYiimooqt4XcMip/33lkS5Jf
fI6O5ruIwCGa2yObPAcQHWiMYd8C6nu+7PEdftY5kpdnG46FoIZY+R1RTv9JloBE+7gqGJGSVxv9
kSZM7p+SEDW22NxJP+VABYfZboF6/QhUqYBTpeeS3IQkg1B33+k663AV5xGit9Y+S2Dfi2/gvEuu
2+8yS9plFpmuC9t/dha9pGfew7tnHWbsS2HEK7sjIMdMpBWIn0l6MgPw/fA4jzgdoNEuAQ2wpa/F
8oao8u7VUCbSbYO8McRKOVWN2RTSPwoXjKOgQlCrDmGR9lstk2IW/LJY3cdRzbK+xpE+ac5GaFZa
oKmDtc3Xul7TC7cKpS6RSu4g8ADisdcB9AZIRVJE32DwDLHU00Nvrhx/+KQ2uCtZEnvp82HnCtWc
RLp/VBsVdbkb3taUnNejed/FJBdztFtnQKvCXvDipQMBw9fQM3Pw2ymQZKn1++41wlrAbWBZnCKg
iKxn+1adnMWpTma97Cqht9KIMMmvxsGIyupaAuxSHMz2zBIlaYLy3vtP7MhePVxRH+vmM6DMv6Vd
WLuDaprThzLxvgUuK2RuvfHa1oY917ZOHY/IFdJcJMPBrMJsWyVnXKqfrOGu8ws15Zvjc0/BfY+8
mBQXGFlOFrcwQbrM7SZZi3y9IjqC9rlg6ZmC/4EpIKsaDBdDRDma28FqqRikZrnz3S5sSNJ5e/Rr
Gn3PNQwISTRRio+0yFQtHyNb0h5IQwYspDOxhVUPCjOHowqWlB/12nB2oMyRA+5jv9wbexOxh7AO
Ui/VcSWp48PLhpu35q1KA2k5KABtV9kAxgC1gYs15ybb1MwfuEV5ijyQ1k0Xj0glEcYISODauIDh
WNG6vI0/aLa2qlrHSt7aDG+hRnlBnNdGcGimgz4Ft4pzzK/o4gG1+7AMi5C3CsHeO1WqOGabiPP1
Zq7d7o8YxFf6egTalG9Uegrzd8xgnmOikvViRDJmSQ3e82xS4o9JcYiBr1tcR5b6//8RlM0OFBQe
Dn6VFNABM8+d5/xmC3WEzAgR110A8p80kWE6KGjPwwbwm7WlmnJMowH89PKzBAY5kh041l6tMaX+
T9t2lFxfiigbG/5xvJxgx6Zn+0TNqIsXDWiqdDfOimRWwzWJk5HAwgBdSZo5zm8m0OOZRGx2mkaN
SL/E7JlXC+Ffms8UB7fElxzVbf3N6lNAcFtaqfgo+AFIeaj1+P7OCRAZ+lcoyReHzTE7kfWhad3A
PHI7LzHdTJTuSQhlDLmcBdkW+YU517ymPW7gD6msE/8chgzD4zbNigE1GfgRvKoF1gA/mzwuILon
31nHmvuNN591puzImLkfNC48QoGWcC51hvbV+rPkK4vVF9RyCSaF7aQFUDNYmS0mIRkzcwMmBNhm
sJkoNtjkxMTLJm7+VpOEmOcSAz8kqDRcvSo+iT+7SYFdPkRF8zwMy4dwaWboIf3Sd7oHykfuPghn
uUOiZvERRCIwboZ85TUyHUPQxLdIgxqcz5X9kZhkNZyECfqPhYLYd5G/de/ECT2iruPxD/MjlaUS
egsg/uFwwB1e9JzURNBCPU5lhXooZqx4YlZdSQte6YCj2oTLxq92J3fMn+C0CE6CK7gjtBM2zzTt
rlsnnhYPOG2Zor5AhzW0eInBKXuCPpCxewptyKDulRPytObFhZW02UhDZ2EFgH06P15KSQi0fRLN
Pj1oRu1hqQrutan3C5vvy/yih+edV0fD6mW4rFCtA6z67yEN5B43lEwJkBUzg9LitUuPQduFmjZW
er03YSq5fJD4WIlLlbpC+6zFRxuQYkYboP5JD8kwnL7fxrwFJ4Zj3cVAQ7x6IcfjF2+XAMSL/R0Y
SUrKivpGy6ujLx9Fv9EtlCoUU9G/19+91vFmZFte5bOzqg3HCoOA/dSil2jluG2EBKSGBYCMra4I
u91WBoHh2Zr5nhvbfqVgd1FfDOglOvgKXkn6hJivaIo9ktqCr9260AJLCNRMmnGgS3NMYITeUO3a
csu82Nr95EAMti9LvJXP9v0Il0LYj5+C7fPx8qO/3A2j+tQjl+aIxnGgV1kUC2lKCVPW/ZitKdeF
W1PWKTtJ2jxj1Ppz+gm10HGwRYzFD8wCC0XnNP/IgU6ptCo7bwtIGdU9XBjpKB2WfugDfwg5iSBm
WiWQ0OacraMqMbsjU5GBxZOFWBA+vrJBwUS/ycVvENhCXEytbu+kNkVH0J54p62KCPdTbpRD8rrU
M0hxhlGg1cU+3WQEfQDsxV6/Wk+aJUmTUqxoc3t7YpueWZEc/HVO/ydkewEivhRX5oN9+krhhqnM
xvUgMpF65YFpYaIZNCqfHr2Qmg6iQdR1Bt7Q0GFoa2ErUtGsx8MVOUk3+OZuo3KvcoQj0kQ+oTeP
mynZUkQnUThCUVovyAVCmY7dX5sNeXAyXL1Brge4pAK4M862khiFrgmRmbFYZxn42n1mClr0Mt9a
6/PB1hgz+XoJiVeQPl558V5N7++XnsT3xEBVyuIZdd8SW5n4laL7MXsVsyqojePEmKTrMS95tkKc
iRhr/173hjkbWhz5ux0Psjd9nDSjxxntLwN2QxNQlTIdnqnDxd8FHz52AhbJho4TFvsQ9IUJYohS
yFuBhkMRDq8KE2ylaKmXm+xPvYsl2jkJu8QRr2uSOU+f4t8NW+3wGQZwItw4KMuUKH/1G0jjgIMH
gtSq4dy0ImyvuwiOrr9O0ZABY4C0SlCPaqu8pV6mzcgQP+i7jEuhKVlTXKGHN+wX0dNByOi+yFrc
+s1n+wIa5vqC3zVV0Ox+0o0YtKDUlj/V38IuY72ydqD8iO7Cc19qmt689nSR7pCZz+KcoEycmJss
0PwOaIgyt6K4M2D0ehYNRLrR3/e66DWqxD+5ChB+GJrMKT1jq3Dz63IoqCMoq9owzs390d4CvEUG
mMqkrafAmCWbkRyJOcGFJYX+FJhnored5as66C0ymALB0VRGdlsdFq4rUucdGbEHtfNoq0hLHuE6
3vQOx4l6EI2adReYj/cfLoG1jtaZ3t9WuZDr9zICucWTPfyOAFNjFkOFTK6+gPpbzWoBMCAFgC7F
utkPkkY0HRLevCj/STf9HaMVPtVsrXunfMo4uer0PZQXhhJBYLMqT/oYl6G9zjwXXo7tZuVYE8/p
ZDI46rS300fL0L2BZ7yTwCHrSTidueonj/iryd/D0elfIIyYQO41gpiGjlNNka4XOmDnAS9AJXMW
e8bhh1e8cqyzDHJO9d7APKjsxXE1/sccE03Ntr0RniztQm3N3GplLEgeZvJWzwh/YytdASfInf0y
ndU1W8REwkXO/w7xxbeQHU+9OKVY2tJrDkjYxU0FY3X0rjODBIAEfDqICeas3lEwdl+HClC3HACx
Fzo8cObP3J0bVkbJMkcJ1g5CiD4l56P2vmcy/dv86/g9xqpo7eETHC9xRJ+I74UgSwU5FT82pElU
+STQGDHpapnmY17hBd1tUFE6XgrbjtPNzqEip/Oqz4WLJRwSa3V19Z4eEUvgBwR0P5BAUpQI6+O2
JE5ZePWmNwgooaa8rnBeWfGj27M0ur9AGckBvDyIOwCWnESh5UPaqmHqpMgCOUyq5Z45sLsQY/v5
SUolHRIRYn6Rvkz8wtjK3mdGai7kuZ94X8wIpxh1KSeA3gLcBBkyMXoaL+0RZmL1LTCqnKNN0zFu
OUWlu4sOAd17PnPGZ/bI2zEU0yBeiLHo+59uF8tgB25mp6rCSI+r6TUcIoPbrTBnDktfKK+/jzIg
Lf7QoklQvRZoFBQbcxH4BLkL5HlwAuxx3QCRGi/iwKmCgY0rHt41P+Kzq91eb7a/CQPoGlVZ2C1/
RvNihE8UHhOO38ibIzpQaIjLHmZM8W0k5MC1f32dKyOgg+Diz/Xmr2yQi+2R/kmT9ZWy+kgfqLjN
yWeiEKt0NauoVpV5+xoc6mIAAT4ZqMAiPX+1e/3ude2P0kPfUpNtTPH4XLiBAF28Oo4zPdlwyn5D
NArT4QMssIG95N1O9UB7NyBhwodY8c3PChEbXESdA3CllUemlkSEFeZxijLgekVJW4v3h4xb0a/A
xNL12rPY/cvllA9AzemxHKNoEHTb56tgb3X0WVX49AyFp4VQDYslFyTtoR9IpJ8Bg+om2EF7sMec
YSaafiBvOeZh307lRPz4BJyncFHGprCrfUrm0/oki/67r3akgbMPmSZHKBPDVh0PYPfQpBpWvyr4
lMKopX8ajKmRmwhc3xpSR7j9mKP6khOj2C4M3n4ysLUrGR8FGESUL+mM4S3tyr98vylxmttSCx2I
PU5IVbPRCs0kSlItwcVnUXa7Snx6hvYU/fp9EkLIsKMtYM2o30Eqg+dLm2vnzhKHNDGzokj2Fhui
4nn11HhJJhsEPFwcsMvHdyXRGMG7b6IPnJmv3CZBVtKYi8WK1mUFEaldczkChhpZn4D1s+iuxVf7
oX5crak3CbBuU4Z/gxVPRA0n1ld0QavWAOBG08lhFopxcY2jjJKbLUidT2agDtPoRmWra586xmHw
JN5j8QC4vi4eh8z0RXiRF0eyRIl1T3BrJhhRVpOrmMR/grBZerrUwJaqrpKY8VxmhuXF6Zhf5kJG
/a3sAaHGM0ONHg6tdd7xKZ5xm87P/tggWG0eqXp5V3+ofZ3uVeDTutcXNEM5ECAB2Vj7OrZ1TQSF
SCKswUU6KAxS5CbqjPFOXFjvsA7BNFrzQNu8eki5Px9Z05PLAKp59g1On/T0CKONdasMfSMpcSiE
0Co1lbHvXkqy1pvYU5G1QiP0vZcZlLMFpp+SI04WR+0Pbu482KrdYFqftkH3aNCpEIvTDEkSDOFT
CQP+ICs0dGGOQ5EbRtcht13fyvKMFwCns3aee7uMVgiNp6b/y+YDMlW1urcdbAAaFMcznloScNNv
0ZCy7iCByI7xVHC/GAdYVsJxArdnwVnShPE3VIA06qs6WkeOQH+U2DPUcEU8hZn7xzUbEakNF0lS
/rxk1TZW0cR/nzE6NMoWHYb4NEHwKQWw2lSND9EG9DhZ25zg/8pocQKeOED42L1XxkhJHQj5x07b
S3hKsbj9KvPF+5QtH3FuaItJclVGE7PJHLlq4yqhvH6crgUd4zYQhQNd86mNeOW90oOGj5QmJfhz
TUSAlrBlgNcRwozC7RFXPTOSdi9Po2hBcsWF9fIrQoDas4+y21aUjU8kJynk2jrH2lIzV/1/BuGc
HlmZOTxOvn2udVw0vlE3uljskzlg4wnuCgEFK5YVO3ZihHcDwKxl99aaiF96ksfAHGGpcF34d9jC
vAXi9LhVgf0Y2pgW+qSLu6DnIDgjDad20Ev5+yKyGDXzWUET2MdDMmqYRzAZFTCVYWt5Gsam5bKl
BKNVnkHRHyegOZ5gqgwv2+OGqaoCO87Dq9rWpJA6FqtRKQRgKRWkZ1ytHAY3R5utTHfTjUdogKmO
1KqEuCI9DXAjiPAgvqROPl2dRtUfjkiKEReJpCNmVM8G7jydKCCDkjK9YeTevqFQBvqX0rDc6bvq
jWeYAmz4zRgyBBc9elbZrdfDqe7R3lqJfGLMwuX3PAGEmIxCJbNO3mtZlDUlzUfOsZ4BnWLqj+Lt
F8MtvlMoGXiZKloRqA91V4Mx5MSs+4mJ58W9uikh0AmRdTu7VYYdHWKc4Qlgj7Low4JRGJ5WshVw
W4bNxrxsI3klmZjoJkDoVOwZPBfYXxacqkAwhHBnnHWLYdAWuy8nYDyMwDU/jQ2O7i0FP21YuQbb
qofneMLLB7boNt4Nqv1d3Ujs1ZDhXTFsjBl0LlbRWZaltgiKRwNJWp3JtC6ZzpAPGhOw8OvPeSVs
odEBPUq/loauVWwgRIXu0ZtdVkVg5jDuR0JhkMkdIDTL7MCCx3puc70Nk0HWq3JyiqFpvV2ake0E
O5OC7M2j3J4BjTXdtJsAyXXni4NIngg5exy1e41P/rW4n7Aum0FA+1wkyb15Dx1W4OYGawHZv8hZ
ZMIvUNqiQAaLJyaiN3YvVWEKUJ8pFSJjt/Tf9rU4uhmeRHR27Fk7Dvl0M1/7TZoNo29AJPp17qxA
egQ2dE1dDicW4fEK3YcjLQ8kb0qMX3khV9Q1Segkc5Je1jjcrraOVor7YxtUPfQG7dYnnjJb4d1Q
ci/toV6LKffJQhnjMT7563JTjhNqx6hcS7JGyN1ISBtMJdc5ONy6Mf0C6wwCOUEHCym7+Epwl35X
NgIuo902MP5qztCjxLo6DzLJln96RzJkiTdllK6kcMbPE/sw0QqR+4sPZ5DH4BhuPKB8Fi98Ujp1
J5EDSqpXH80KTCw/pp1zh6nlPtU5Sna6AlRnlUiUOOkUaEl5JMgjRZ0mRajwmV4tAuFepUm3YNmU
5iu+aLjZliE2iqGX+rKtfJlGmv3lBgRcrAwGjHeiZBqua38y1/tpuKe/bLdyK0BSmonOlA5zcdrR
Mzpq/P6fAdFlH8LcvGTqjPFPfWIl4HQDiDPqxv4Cwo7CaODhzKBKsa0ARmC4OOu1jl27tx4jV5jO
stAWkMyyd8ItLxuRsCFrnEsVwE96a7iXICM14/ZodlFvfHc4i1dZbxUcJvFuurqwxpAa0sVZpguT
XzcL6OPq4z/YqjYzW622UPfKiaWsSCE6MIeXul3rEtdnG8Y79aJbWXjsMw0+mh01LizXY458VWkY
F2DGgljNZUlrcK61tUiP+M4oDHkcao/DVa3DoN8EAoIVf81hRil6oChDujNYuevoCvL45luRgzDq
yCJXXHR5nMp+dVKMJgw9P8LwLOYyuqG65MUAVTK/9vosd6FlgQhVxNFO3KRTcZWpGBbr5IYPFRGh
A/JaAhHGhSvfN57b1JPxcNB+0z2gC0LwvEQJh5AuCxqUUiKVyHnmhM9opJR/P+lXXgXmyb191Qav
cCe6oM72zAQnR09UMMhdAwhRMlZd0tCxaSfNb4HcSmrR3cnP+lZ4nm8XaWYEFbo/41+nfyC8Fmrb
YFGLc2W4IoViJaPH0FUe47s6sLNzbLfX3z5X5cmEyLTOoNh5f3B5B91kb15Zlni72ISnrx4Uj+r4
+bVI4tfpUxyQ3z3ozHWl6/OVz0dFgOOAeVJqdrRzsdPiCbSLwKaxxul3otmtbv2Q44vlUbACID7y
5IECrS2uoWanrujjpK1gV06P6biIz0cokKRIIAnaaCDsSN+gdHXdASmDebYhyZwRHtooeicq8H3W
9ZgC7T5zH+A3Amzr09k73UKxPv+wIvRoM0G5R4oM5paRBjOi7dXFX3LpJ9aWH9FNDjy6F0sFYKjR
cLp8ISrszsbad9Xn4N63UXiZmpnC5Xvy/PFOrcS6gndd6vkNoC4wi4y/1mJzahITxxKemaB01Jzz
ReXbait1IyjEfYmNbkIFf9SZ1pBRJd3qFsuTb8VvMrB47Ns3XnoC8Q2IFZI4UNvJngMqR9g/PsCn
cAcYpD9McaFcdPX7/9goaE2AkAlE3V8HI/klB7/CusHCLcZlVBzOJULzJOFakrFfPZ8XjBq6ERqL
rypkZeidoV2ST+obH5vdRt9wWXFkeZhoCvBrpP3x8yXsVNU2XQ5hCp8zHUpCsBt/tXXfXg7Hs5/Z
QFmjYjaP89YqX3VCkpBjeOJADU9BRuuC8j7ZyMkcQ18V2cN7QcGCuG181JzRCM9J3TVKRa9abNU2
ln2oup6VovFrdqxp47hENw8pCnth5+pR6N5hJFELd9G4cCz9lLCDeS4TQAywKwR4YYJokZYckF35
uRLnXQPQS3eCsY9G46Y1/cCnu05g0lbF99i774hOYzNR91ROt50c1J2cToETkooJB3SUdOgPx194
1f3MeVQ710ysdrlGc5vSIgFvV2OpPmUeQ+TIKCZqS4CHd3YEO+OOrLzruBOL7UuXNiVQNXNzdzUP
NQf4Gq/w/FjL7m84vfVdeWLt/Q9OrwreXQCbDUwaid3m1Kinu7eWLtdoNLKuvUBuf+qbB0ZE29Sd
U2coygACCxKA0i4vFsi3F9eq4sCv3Vdv/QxRCwRo0SOhbZlA8TsAY5Yqts1NgJ4KbELhg9Hstx5w
naM7IIdqslL/74ziucBEkPRvyws5KcMAm74hD9gCKV2EUfNrqvd2Ll3sRyo/v2DKfSsalJm1t8yd
SIt2WoaUUfyQ6Q7WSQty8ArrSjwogwuUrGpdldmP2E2dka5EpfybtHy0VMpgsBQQ3u00xu6fVysU
GcxAOsUrB8yqSNAM4hruQqtmTkuR8DYqigkIWRn97HiC9SvAxB+yY3859WEJ9QGGVpHSCybYFUEo
4pKks7ET6XSNPFANRlkw9hMkX9VRPrqzSXAYyeY9SK/mzbbTLn/h1XZkRXFD7Ervl4WBtePRsDai
8AG9sCpIF6cCDaL3i4WdHtqFq0uiXOUnQ9jEpDZNA4SLwO5RC9m9WlQSEVKJxUJXSBfJ9GX0AY63
NOVqQoMC21us2CuoXRVONrvuqyNx9XuU08NBNjFIz/4hzNK8Jr2cpNnTHNyMMa4xrTrPSZqrQvE2
CBG0OLTvpnKf2K6ONQV60fSpZIPF87unGvkuJ/842zF1Iuu6z4Ir0fNQj584cl0Mlgb8gC5l699z
URbpq53E/BNESXw3nQjAVUBU9VU7T12Jji0eBxpi/sj48yT0bOZLNQLJOuf39HIROQB5TKUgHnzU
zKw4ujscFEuCp/pJdbXs/BvT2DAqvlohSMnZ11BGJj4IKXFzz4u7WCIEE1wVhj+aboGzV6HZzScY
+19RR4ffqDH79N3vCFaRIYmrsO4clcK3xGANSP55bhzkOuqbbjh3VC1Y76hjJYnMlNjngAqUkg2c
Unq8eYVMKz+Rj3qiw541YDoFO1xntfDo/CI7PD0FTQCvUBUgxXYyjkndhvyvw7CEMr2XefgjnNMX
aRdfHGuV4/w08sfd5D3Bos1+UXGdnoRfnv7LXLapJyd4ysnDqTslvQR6ZAvF2xrtWlsCvUV2ubtq
0CH53BScbl6VDyX9FSchf4Q6uRojnsjz5HKqOpkjWmsD+M1OVNqJYw0qU/nTz82wdr9O+vAXA0Sf
n7rzA+Lg29gPUl4yiU3UzuzcipIuN6gz08QyZfh7KOcpNsCq9q4FDIC9+FYSiFDoF5OWkRxNiHg1
xdp1SFYlvapgidhKmMKYe9wMFvfANup1jo37A6N4uoFYoheLNWDYiFsAd3+U9hUvNqwgw2reMhGJ
c6CqpgjyEf/wyV92yExzjrg2xaEZFKDxh8MdVseAfJFUq4xsu32Nu8oWhKzeZrj9yJcbGTCreXfR
uDhnnwkqn0K0ibzkRh7rv6O+Kww+6La+xV6NfChyprzO0iTypoJT/IyXm38w6EX/WnZYVum7EcED
ZiDxqPY5ub/xibZLhWCaVckeAzJZI2OIxbhQXhgtC+ZFcrt4wZrVH+XnxMqkidk97HnNKkAEhP5n
MbqJzaBPkOcKfhguISFa1qFAqeStJzy6pXEHd20nL6xkDbRTMs6exnDGW/cnsq/6TlEwn8p2UNfw
G5//N1LlZszF6L+aYvJr0O1XjgPfoBCBnlZkfnMSrsHBbpulkJB0YJrMq5hH1VzgtUDu26NGSA9s
pBORrjxGOeRMicz3VGA4vUSJ7NnwMMJ/2N30kMa0sryyu4YPMQYVjKhvj2X6KoVyBi18wAl0dBeq
jPoljiGUxcxQrhKjTv5tEdMUeEYGG66SXcqzrHAdow/WPhYT5REvLJod9UMQc2YhRxIxOx8VS+j5
tdW6rieQ4VKOwEF4f+BXhmE6nCyKh2fU0ygDUDC2VhvRC3o9jTJ0D6UI1c/kmez94HfHKPv7lLuC
p/tPTNn1cgWSTuxvol2ScNhfMIsdZWSmbnm7mg//mJepvt4cbZM3JRyb5/y4bKxdcOoRPymiwptl
J8TGyIroWi8K2qIAVlG101pwLTsIbdjqrzY6hntLfE94Fga2Y9ozSAxvLZn2rmlkFj313b85Pm+r
4oJjLFLH8WUFGODznDLIMxeV4WXIwmqe9LIar2eSB5TgsnxlBazBnw9WKlFS2lIXOSyC0jC8s0mA
lniNwolE3qslkT69kNor8wN6KSGdeqIZkCTzmyOr9d+ZB9qPa37AAqpt07l3rMEsij00cpbWZqpf
An3be/WtcdIC9xZVrJGEXe1rsZCo1Dn4NfmRM7TX3sW+O2AR4ohznMNwkk12B6rMAHMwuazowhLP
qcLy7Hz9oS3GG79/0hYq7Wfl14t2srPk5/9XCVVzXZ00oJ/OMa+VHPaEtVkS0a7FAJTOu0ly1fGO
0m/E1Wb7JiEY4mSIE1q7DTtWE/e2aLDfM5VBa3CiTtJ0QWaQgxzW4s+/vRpQq2ynFAOcFwGPtHAu
SVn8VuSWo6owLFBK4sf4DVH6GjN+0cO/sIanBH6mCmnwr85WYtwnRvZypNr1v44cWQyvWXD/NmpD
o+JEisoJ++5vJoe5JkyZQeIsqgC13JcftNubJ1QugAJrxjv7BR3H/0P+gw6nlgiYsDoqVMWPVBXh
mbvmntuGma+I1w7fYsHBn+JqKsOhhdNRijmK49S+9Jou2zqfLIsD+W5QEFp0HkkwzQYDWmpAOZiC
N3aahJFM8kICofl5wblPpw/CXR0xBro4PsGhRRZAcEgUjNGCXmvz1ukmgxQUmpoZpaLok2VqS3Hf
SBly0try53rMpZFhWEWjd3BAxOB75Ox0UuA5a3zwpsh8F6MBYZEvFsyop42yzsxvhlP35sTYYnCR
Jn5CEqYKm8BB47DHHWtqxcupLKJ+Z4Bd9XT8UC6dNBi4MUmQrHo8xr7kYTFbNN/1CFlqEQn4SofH
6RYufmBFAxS8o13/3O+D7NFLWEUZh1hrOTS+ozaSvSkSO7nnr1ItAZZwkA5k55LbW8vc5xhOuupQ
+dTY8kYLwOnpC1qbuIbZK8o//LmuDm3ALJG7HM0dF3GgFicVbfKv5OdCMNHJ3eDphNXi8fXopCo6
9lBtFPlRQTadlGft3Ep8Wp01n0Efyy/UBFbJNal4zs6WS9+ALb/xWvs/7Kv/wDgX5Qfy32XFwpJB
dHZSe8+D1uM2nFD2UgoLtlAiwWMVfkFwScqZTerMezBbroc4W5tRfouzYQUKcnnw1EeOS7VzH3ld
owNMW9awtqps13bvTUzq4/UUE+rUN86rNHNeyq05cnzseacs17SCV7IWQwuUFudm6VrJ5iOmuc1H
ojTQ50aq7CyfoCPVAB3V0VoqhUDWQ0WXXHBOwlq4fn9myhFtWx3nV1q0wKS7qFkpzeq7HvFgwYQz
fRYSeGMuUN1qcl374Jys3cCou+2aNCPRuvAUmXRxXCQZJWncNDPDkX1nwQFlMjwBLaleGt+FnK4r
R6252BWt1twyOltESjJWAL/KI9lDO7ZRcwBzlvejMjxxwYC0yc7m2uikXhnhtI9Iwk+egmHzWPVo
xcgta/Ktd3eBvKxxuO+J+BcvOkHPVTMzTpvrTM9Fs5I03F/Es2kik8M3wKhxyD7L5COSXoYGmWe1
wj9Go2ireYs5yea6IsGXDjNvG7TL9wzKjsEZbIP6Z7PJPu3cWrEpLgZ3XD7zSlrnAKA8/UxeRhDQ
7AmMUiY8ZPUDWobP9QK3C6w9bO4ZQESxdXZMdFppvqml4ULCw4/76w2sXy+1Mz17/FDV1WmRF+It
O5DFhFZiV4fpeO5/ozQbqmifRic2GHmUMNLwtY42wPOPl6fuxa6WDTvSNigYYTx7CbSoC0xwDWpd
maQgo3wNnTHgyIFVSAyTy+T/cg4+L6EHppYyWHTYrpNxlaNt46BDzBzjnTYJ1jyH+F+fIHihfy3C
aJ4Eehi6Sl0imjxAoxD32MAabYveguvTOYW8Qeb+g9XIy54C9KBYWiUzDWS7iTw/4WIllyOAmTU7
kBN9xXgaDEB5q2FTTRi1Du0IEYrWAH76j0UvGQmuL6oVBE+8HZV39XWbkE93B+x74Vy5irGhn50D
Rgcq/Wn8JF/EoN20U7uGy13KdPkOTY1IuSEJquCFFp2Njed0KZ2lpVaRdiG2oBoOPm51cHdGOS4F
8hr4t8ggI6qL1MH441rZelG8OxprFZjpJVvr6FIUdXrG7Nn/Ooymeh/OBVl6+dDCLKvqm5ty8YYY
wJh5lUQZEa9FRlcpHxqlrL2tTZel5f/QFxMTjaIexF0C5pBWbXmwX0ALLh+1NiwrNd+hHdw4ZQNg
sxRQg51PJPHFXrwHEOiAQ4OCgPyJXDeYpZU5YHuCENOtP6d0Krin4yI1/6UUPLD1sFBlwfxq4lZw
n6A+vjbM+G58STs6NvOs1O38UKwX+DEGexyt3dqrpED5jqzRX+el8Kx4f3ZIyjcr/3AK8OSrFTGK
p7xB1XQYTWRAwUAz95jUlYZ8G0d7vpGomBmLxIkhDrcAjGhUfBWp4xDC0FccnPyAPICHuVVMGyJs
Jc4wgc7uQCUhF1lzUwUTX2Pd3T+dR2a7nvUG80Uq7Fx4SQkF9FeKwGClTgbIZNRjQb0Hvk9wJEJS
mnGTEDf/twRbboWPpyt2DeHcwXJHWzEnZ3kYbG4/UirWviw7S083dFWL/VjsksXoMLrm/ljycAuU
3WxBNh8F7/vcoOaP/uiGRJW35pIZdw6GqBPv0NHE2KQlvQh3iL+Pc+RQVnWrHNA9RiVuv7MPtub6
ybo7YQ5ohOCqHB3InZPBPKYUKJOYvNpfPTPPLkAyZdzS1vvu2F3wSPmYfUN2Q4EAr5iKY13KkSjp
mGAzSRsWganBniY556s1CUyj+GowxrtEGpNMciptrJ7qmCCgVvTqWYbYyy+4KvSXpqHAgHN0EF+S
m+ClE735l2eS3md/s3kXfDJ/NCBPvVa4l3GcHT+HsnzqBuiikuCZDeeBY56ZJmksGlnXLxsMTopF
oZSwqkzXyIFMRWQTA2LEU5okqQqCxEGgsc2Qjy8/JOaZ7tVqox96nb/tFCX+N3a7SCLODLhS56bg
ed2X4+wj1abGm/HGuXoqaQR3BVIDRdbwbKwPBPTIW+DRm2ZAkwmnoOUu9bzVGGM2TsQsPAXKmWQ4
sbR3suyHkzYq4o7VxNNcpYp4/QlEiCkNUrCc6qZyM/4R5GH2om39oaAjj66yEMv5X2hKkj8Y3U4I
fvjdpf9vXynIr1cFAuUcTeeduR2YjlZiTqWuXsDmTmuHzMiUKTtdCRVCeci7bHVKdt9VWPi7Glim
IWO/5QP74u2E6b5ryk7DvBNeZcIZXZlRem3lUJYCHyOy8N5O8YGK09MHaOqzsPwOA6S6ev0ICV2i
SxpJB7lmsyM0TPrCoNOXZuOlCgrQb+Th9sdwQ90O2KrODm1OTUfoxOnmYf3huphLuUO9ri9gj9K+
STC5Qz4temPUDcD5bYz++MWIrRZTU41lYS2RkmnbnVo7a38mtl3IRjfEsTsM0wBUCsmrKsIZBYqf
wEAToLLjnZKotB+ny5dWF3ioeS0blvXPnTU0ek2o7ifQUC3U982aCmyXbA7JP0lempYX+daRCuFQ
y4E+6abN214o2sEHUDwO3ddKAS1a82hu1mvJpplzjCDJwEN2RjYzYauTIXZ0k9cUij4jPtkL3HHn
n7GMjtJZYZBo7uqsgv+jpuSifLc/xef67/GdhWHCGEsMUQHT5ROvq2zMS/1c/qBKZPpujPindGV8
pYhWK+KuaruzIypi4Ld/mtluMwZg3tFAO8FW3SmA+SXuqscBiBqFX7PLgXAfBFNnhp44HMukQPeI
v5fSLYxIHYlNp+YoCLqjXkFq8Ptzy7FGpCCpGejVinuo+qIbVU4sjjCYRVubzymf8CRyBVwLoXZs
4Co+rWYN/zwsOxHcq2mayLjuzNjQNMxYv+eOWEBKLbnrIRwPAfgNzwkBjCsMfKG6swLMz2gNTo0D
3rHcSjnw3oQzuXa+wn7Zt8OgWLJ65purcjVUoMMEf4HTul+JnXPyAeR88G1JRO45YpAaXywjB5eX
0P5LkeIEGvKfVd+X5swMpVmFxOdijIyMjmNPDJ8tD2DmNwV9xPsJUdQBbG6tGIYGdsQJ55tCrBRS
pBr80KBqawuZrSzZAVChFXPQXSa+fepy4eiTZGVrGpuEeJxHbfRlnPnV6pCiXXbluzscX9KqSosQ
H1taGBI5pXn3qfN0hi2LfnEVOtmCwuCuwind4bDIidcvOc4QVrnsS4mLTbVOgd8csyVWlZHnOFsT
MWXu2QS+ENay8uqgigv7LtWT908mjF/CD51hgAhfXFTvvhPhuw6H2yLm07tqhnJS+G8cgDcG+uZg
k6CChnE2fPmU01rsrTCNxb+XpeRxFExgwZkJ6/nEgZt8WJn3DFUyMg6gSsqARyJ12jBTUoxmgPst
SJ14HOixVD2wARM6JynRKhJJnk35vJhddh36oZgu7veRyNCXvG38c73dN18RqDK+Yfv3moZq+sFc
671q51TQ6N2oZzhwF8HMQM5xvoy1g6yUVcJXmWQ9+BGeOc/USJfWIxpylaO6arPDL9G6iiWiRmMC
pMN0D9orLF6zNEE+iuCw51iUpn2+vqhj8u/x2sqTGCJq6fp+aYRBBUhwQoH0eSVWskoNUDSyo2Bh
boeXElAozr4RsAgpIQu5uDaGmk0LEkd0hnxdfPpuYzsHtR0h5e4OJexWKmJAdBqzuPrOmDfBHpj0
A6CCYUGTZBx5kAt9oBapC6XM58myV9dliUQ5QmGlleslMziwGFKqLKj53Rr2dmG3TVKgRpIfGpk3
SIYeioFUl05jUpFdny8IsESVcG7UslZWeKUvcPGV8idKLUEkfkyLqeJonQpbTgZMlZXfP2vdEJTU
HQl81sm/mAhHCuNZDaiealjHeIfS+CuVsS604j/YhKDIU9ZAwLLtpZzJNGVKj/SdvULgCaKMHdy0
cTdETCxSzsaylZzfjdlxZhaYQO1eDQ2RHNj3kU9/70S0VBnoIclGbSSrLY6SXbjq/fMxMrY3ubw5
B2S91mF5MD4FyAmQ48RVytLnvk53QhLHEFwU6AkHYeAYNMBVauOAp4+X5xvI9kH/pJrOTLvHxOJ9
7pApMsrx+eBairoRI2HeJo+OkmxXgZRxgSKubpqueJu6sr9qw47DoWnkMLEQ6FcyKjoiCBzrdiM6
Jva/vikKf759Y7U9B6FwctQFG2Zwwdeitv7tc8DX1zv89s+910WpND5YAKZOJmPg3dYMUTtaHSg6
0WN+fe04Ce7y4ZJNSuXe+pZE00K2H6+gF3dlgYgnGzHnRroNEJlGa48hsJuO86Ivp73fXEZJ++VE
g290aa/F6pPYcYh4IijW3ORyfnvFjrD6qivqZEt2sotLzNAJP89ikKWuTQEIgVEmzWBZ7Xf1wqFj
9LFMPW7lfxMKwrzN+qfQXDDGsVLn/GuBHM+ag8NQeeH+jcWKjDM8uyiWEqYqXXckhutBl60Trouw
GlNrRka0gJbfCDG5FGwf+vxbY4pvdmZGYEnctzC0eZuedZlXnToH6hWl2A4zZz2G4B8ugEtMJSMO
nWggZ9RgCwO7La7tlUD/iuNxvfCPDR40G89koeGjPGaVPftL4S8mlDqVjF94/q4hMgFI2X5pK+75
2Pf/j4224vFz/zaU5/h7Dhf7oNnOHl0jbAm/nszDGFtNEOWnyG4JPCDCHqt7d5eOyLYQJxPLz/i9
Egh0QW+BqZVbG9cuS5I5lZW3ybdkbxSQe59Bf8k5oWwuQnJbM6kaf2WtnVOXEfjSwdh/4pDZNfnv
FP5C3ATtwomvweMg6+DOtXvh0wvlNVaUg6I/SevqrzHUbdXlZAKbCbUeqv+z3JtyaSO4ihdame5J
/UORmt4Bc73SOkJJA2Bk4/P7WKSdDb2RpwFPEoTzH5d/3TFh8kCXh++5T6GD+/msz7FU7BiuQPo6
YPrdQG3mnqJJPx5vVRmhINHnTeWNqk5OcopdIJvfP3NPuRqf5WXVixH+fby9paznk3/DZ+1IwR1G
og5TGx35q0PpnYmxVZ9D2/HABu01OzCUr3GfujN7szLDs7/G51XHg3lwlfCCp5Ncgx12/AYhMZR0
rR2T7JyGavGMPUlgCEAeUu/CdYYB9ZhM5oO9RqxBxqd6a+9q3DaN9VHhkibw/WFLJwgpm8cC7XyZ
gBmNC8H/RRgbrfpNubUneAL8+aSHLim/A8xi2qS9rGS0n3MYduUvZ4Xt5Np8hsTDiopS9EkuQ74Z
TGJwiRo1I/xY0/w8y+OQEUXIRuQAgCeW/gQmBuCwC+mc/1Jz85IVKMzp5KLz1Srh8Ih8+I+G5n3j
QLd4CitHVBxhjHYQkmiFnBQwF19GoWoO/pOcc4x9dIBcEhidH/OX30tUc81AwzuntCk0IvoA3ofn
NkiYiinf3AwmYVvB6+odDrRCzFQAjegMdtZssJRMJ7Ayoff/MCYEbg7QcuDfrUluyNwzAEJI1zYf
PqFq7ymDwHUxXIBWazqSQw7K967LFrI0iZyoLqkTXHCqK6CRe1ZxQOdxtI18tyB1RyZjq1lB8ra4
MI7cqircdLsxG0aQ1uJOsdKuyNSjtegLZCT0FtExVAVrcBBhHvjydhsC/oeTD48Enn7ku2LFwlYq
+1XBjiTEfonZXYKFCQ0CXsaTR0M0/Yw02lFCUdPnw8FL1KxtyZkwm+ZREOCb1nnIeaKzfCUM3aZZ
UxT5JJgwAaxWAzOT8hsP6L0I6NTgrgopBpE7DMoE0hKTIix+YVrvsbqAI0ODGrfizRbLq7cuw8E/
dEtLOTD8wnOrHHeWAlLBz54tJO9Z4kjy66xhrS1lCU4LCHEgekVwYLga6uGjOfrqYy9dPDglhVtB
0BnIh7t1DK18+UjE44TExqT16oap8js/u3hoqCTlZMOMi5E6zQ7wtpYvRFcd4VEiE1nEupgALbN4
gR9CTbAJRlp/3I0Wsiy1nsbMITmi+lpH32FtE7FhcXLiB1QgakDUan96/kWHVyiJlt5cSI+c7SBo
/QLD31wJCitCh6CjPm/6hZTu9+nExvuAuwq6CrYO8MzDMDKsm9y/jKRRjXbp+8j+dL5Gy3MDL4xO
vbdRRvmVTAeNfUoXtFg6QS/fM67bmykbzaaAQAUTWNWIvaDEywDgFuMRcbY7I/3xKlIcnAiIm4ct
yp2QeT8LoFuQ4CzKBoZe1DiB3speTAFDnooq+kHEbHdIjZ0+dopHnLGGTj5qVP6dS9zMh2f/MrgC
T1KBdK6fUoq1/W6DbSL/phgJcvyiFr7pPo6LKAU2OMw4Ff5epxF3EOFcpPWhO1JK/7FWoyl0lvIu
/MOS8eTOOy+Zp7onuPVR5mMSVz3jtJbWUY0Tfig5C8uycMlV8pbDsp/wev+EPMUguFSGRdIjZd7D
P5vpExeE+c6lXJbM2xlGjwFys7EzJhtKQvwARNTH0/ZrECDSQy4oodca0n8jEcb5ROoK5Jr8SdrL
We3yu0HDEHaJYm/d3U46p7aQ4Q3K76mGYgy5ADi4fwfge8yHNbPrulRNHj2pxcVtUP1EoaTZ5S73
EQRvdg2f9WNl2+MMtv6BkZjp4u0ifIq7QCo4JiJ27xe/0r+Enh5FB47nP3P8s3vC9nqdmQtXHGL7
gC+Vrzt/ZuNuht5UWA/dxwuKOzRLYDrIMfU8L3bP5oQgqSyXpzV0jmnmyVCE1RLOFKNcpKC0OswT
GW0z25+4HraQjxtccQM8ICJLa5tE+RzbLgbEoNF9Dx/RCvihfIq6RSTVbj+UDeD9Jzfs8YrnGFVl
TTPbXJq1ma7HsuzdhYALwuRgAlLlvigfbGmm45y0qFCfqFsmFU63B38xlTWr7NDEUYBJZxd4hqIA
MAmRpk4IXNv/yMgGP74b0V0Vcckls/Zvp/4jjxsadhkwbAftXKtT0C8k8ERjUAuJDQhuHeiZIPOs
dbUDS3TipnUyQzD2Fl5MbCh75D2/SF3iLGKJH41RH2xi0ImN3ZNjPIJMbWRjSwjtAAoR0Dgs5HYi
FC0uK9fkY1JNHZ/kdnhzeFRCwCSeultZJBYzSi8dn6AgFVKMRJpsztr0n9FyLtFD8q+HBFAZTLb1
NE9HdyxewMAJapwY4ylIr0CknX0d0sttvE0NMdUtQg1wdXta5dUImHvWRhofaes43lA6dRG7Py/V
p+uiBqrgZzzc2jb5P7Her22tMBqHjLxuNmFB5zy7NjbXoleNcp7OWrYtKWmhIfGN65+5fWVj55jG
KKv2PBCZbkpNO3K1AVyRF0zr6ngX7g0UuVvTh26d5P3W2v/txj38RqhDm6hAHmXWb12QyEnX6t98
wqVCt4zligb7ZIXF+8soYbBKAaShBGUGOM+sQYuWJJabXQZ1qGsFH3vkm83s06tmbXiZj3vUD3hc
cCBaE7xZ5sqoi/vlIdU0msannp7Z+QQ5ugqvHpASUSyEHyVeEy3+9hQ4kPmU2XwH/Yd6cUNDSA5a
emuS8KxpjtSY1/mM03zSmCpYjh093kqDrvrUlCGpdQ7RQ4BXfhUGsHakXIfbnwEUMwXK7zw7DqW0
3afatPlJXtq+giTJV+X92XE826Fj8yPJJsmoio7eBr96MWO9P0D0TRtdWiQJfw00P640L3nMJIbW
vVt2QKE9if1D3J7GijNhqr8neqfzm0sHSFk6Y9ScO/Nw5YK38WuipaLbMovV+R+Z4c9mqLRiSAxR
imq7lELMGX6lRazuQg2yg054OmA9ITm4DoyAupxTCTe3QOZ15gn63xEoCoaPN0xeTlgQLGI3q1j3
sGgne5TNVyprM2mOXPMV+ZaJkRyYurO4GVOJ/xbUxpVdkphz93plpPggHMaJpWHm7POuC1BdH0Oy
tX4AqGqkLUVSBYKEdrcLdJpsyigtERrcYU87sWEps4/NrCkS0yJlZxXQWohX9t00a1aOBKteXcer
nJ9RNyUYqaoMeUeVCty2hBy5KZEYnyYOaAr4paXo5nPT8zLc67x8AJLdNXoXVJ+NrDQ7glRVl1vB
bhCcWx6HvMS9BL1kj7ZedaNSHOJd+rvz27MXw2LDkZF148Tb8dlALuJ53MQQLrr3COcTRDfBqV5U
ey42tJykXZrUWmvcGx5rt+gTG8sWxPKecgs/j8xcYlwGshQQihCNhKpHrpYSNDlDL0fgdSHzCMyG
S8n6e3vxyb/4nxxfy4oefl1/VvAoD/Jrpjat0vf0E4zfblCeFJaFvdO9PqLMhGP+oVoA8f8883yA
+NEfbd8rFw3I42v2jiSexNbc8xM4c1kYBXpGpB3HAe4QdnJDdF+4AwYjc2s3fWZ2HZeWAXm3xCMs
WCDDkCiDBDtNQ4/OZhotJ1iggjdO34Ib69UG7zjmYcOBH99SHdO9k+VbgemRBZX0Ep5CzaN4usuZ
OfKPJHCcbd03Dl7mE+ZguaAaYcSGL04d6rAwAP4RhE7rDJONlPnDuxD7Yq50ah2MrVQO3Z+lCqxU
wUYyAIcPLY93TPdGqoQoa7sotEzc1H0quhXdcaMx3DynU1P7bIWx+a+CJfMEPkVniCLG9XUWRLKo
J9nJDNm4gAIBVRZj9TJz3W+Y7FWj1F06QHUGkd4xdBKgweAFWjwu21TNq8bvg0ckQhTYW8jLQuTb
1SBoOPmCEU4cYPedivVofd6rX0rYeYXe4kh+QfvGz0zx3U0iwDRcLggmlXhxr2/XtDvaYY/i0/FM
RuivwMvSNAI5qNfGN46+vCQIeY3RXvuN3XdSvGq7hH2YqO18ITL3XYppGV4kmJwz1tUjfGAttUTM
imUmHecRXGsEtkQzDn8h4nUGYKRHqtV/JjA5hVURGFm+hKKIDpwX38OLKENQKNp6WHQ9/3aOQ8mP
+6U/DQRPSnpAv6wQey7RZQXACb9zL0uPN9dFSpbelj60h3hUypzR2K6D+4G+iSOqGwyTCSkFY2UH
Es465iRSRZIGYes1pc370Kzr7q1tq0Q0P23qyw5N0UjyC8/8hrE8xbBGj4qkYPex5gmOIDT9SSKb
AdGZRgVR7Zln84hfaLj4FqdVW+Q+oxlFXw+4ZA4lOeq87ehIAgIXJOZ2OWniEMKoDIoZzFybAILJ
AVWTJUfCTEXoD8VwvK4Sg+GkUlXe6Z5dazbxe8ZOgAfhdvB4X3epJe/fDC2ruTdLIvI3X2h3UXRv
7gTxop45IBbxznBUagbiDFZ8b/lrE6ptNJltxqv2kmhLJOwTm21y0mwU8BJRP6Uk/1HjRpLLCruK
vSEB5Y1Yqjek0uHO/0zZLcsh2vP1b3o1vsjQBVhLmqFb/9HcsEtqjP6LSnwDYvPB9nd2o3WVuqIs
TrLtA2kXObTyQr7va0IuBMku9jjdXSLucXPEs5XGOrJ37JkbHtzui+57AvkmJYQ6H3E0DDkxKx+u
9V54q4Df5e/K6hM1J76VrXLbqBbNSQ1XQsN8YpF+3m0efDhtRGN1W5nomImmVXTAMHp9trQnoz/Y
9OUBbeq2yHx/5oYTAEOLrYPETIPqRUyeRACHC8QiPVTxHxDLdaQthPLlCxb5yOo6znUOxJK9GThx
0wW9Y1ZOrcJZIu7A5Ygco3c8KFcxKYsS1ULd9nDZO2lKkMwBQREcaDKLyOal2wycWhnouEWhJ0Yb
SH8q5nFtCnly3o04uosCRIc9ZXI6+3LwEpHBwxa9UtduE/UsaEiYhoZXhgTtMjMS2IKIot4iru2Y
dq5tLeo5HnIOPSDTbqK4D4UajU526TLgHfQ0dATVldYa/Fn40Bw8ZoaeUcl2e/yBWaATma2CmTkm
vNpMMlNipD70Sad0i5cPa9RsUtPb6WDV/7aRugL4mLd5L/gMAIMb4fMI4zYbBDFd0pqt3u3X1QnN
kNir1ikMEi0/FPjgOoKmHQBaP15/KWolRbTm0PnMlDd2xpyAhB/yZHkmEVFejDdxTdw++aUiPfpT
XvfsjxaI3c8Ow0ih6KXHgzjWM4g6B8z67hqmftQnyHDCzildvpmLSybK4e9GlliBlWwUo28UN4k5
uCGf9eedrhRQoLoQcw8apy/287HmuAfWv3eDXG28fbA4zQRsnHWW3QGQbGVr3G+qPx4DWODFk5YQ
PP6sLejOzYbsKkgkwU9IXRluTj1ZCvk9jvJGP1xJ5DDdaN2wchM9LH5qEeFIvatx5KG5M8ZNxR1/
MXIRuvi5gIWq8Vvvt8W3yhlfuZRxYKQk/DbnetBRdYhpxw37HOHlANVDvtoFCTsZJ6xS3YuMH6Kh
vMxQBNqJ+URg9DzHCkpT+a+w7i8R5kugQMvuSeypzr2g5ZEF/TdV3m7W9HpDdC5AbTeJPZdf7/8u
OogOYg5azisiCqsYnrqU9ZOLK2iaF0UPZ2Z52MUiFKqeOMfXHleRYvSdYbh1U/3ueVADUgqx8HaJ
Gu++rETOq/CSgQtDBnY20b//uioj+wm0Xx4Cyp2KprIHG+gudvUoLHb75PQ19GoxB1qjP8+znEH1
5dGZWyViRni2pbzOBlrFJ6vKITL50aRnh3YOQJhyLRMMOxynl6rqJaFN2daIbx0v1QbnB14njY2W
HFBN5tsPJodYXZoAJ1U6+WhFSB7dhYhuoVjxiagBsGlGQFBbQEFpHJi4PDm5RxzYhOUszkmPVniT
BnSQE/GjUop24ujLNm02bQgC5mKihAJN73v/6v/tKV9FoxVlG+q6JJimQ24Min9vRjISMXcOF51W
B8joYRAuOZTKwrG05SfTTrPjQi9xWPB5KqcADN9kxXFXj7Z6o/zMpGKgisY5aGvzKOq5MapsyvIh
dOVPf6ltdb5y7+Dlsn8XBKFi1o3zFlrFsxIIPjZCPdTQ8kWZFLjfC0MJLlClWxwTLT0jOMHJ3TCv
9/wHm1dkOTQohB+4FYMb9nKqIweXCdToSISEnjYmt67OvnpWup6vFr+0SYkZ7uFi/ygXyHFkKVVC
nmNl0IEcH3mSzWtYQFGecWAQYB8KC2GqYcbP4N/6PVdR++VWFrFxUIQYOUJrefKGLJ7VzJ859bK7
dNieeDNFNGv8jAk6q4uk04CpM7A4SqBswZuyk6QQi0Rr+cB4DkBKjicwWOnf7HfOT34jDzRR1mAP
zRrbbzvWtYJE2wkD5EN7+rbsznm1FkFhmBkYwHN8H+6ZgWYjZAu+X4H2ARDXOgBxD1n8dQLr5n5Q
s9xcoI7WHjW5EaypASJDeyj6l3X1a+9uu2/JRwqLxJIDLgHEbl26O1e24t2Mo5wC6/cvHELT2bqC
Jq2cXKXdBChkn3NUOjoHGaKe2hCm/s70+TsKFzWu5IG8vP03+4Y8qadQUR44mf5gq2QM95f51UPP
KplNU7kP3PywcuktoVROPxZ9/F6GFghvb5UZ/nEFly0RrdQX7pMmoCmSrPP7UNy1bjUAiUqvX7Xq
ZhjzL8SYTf7vUm0yj5MWr+/YDw/p9JCbDuoaU3pKxxf8PEwNeBonsh0DdF+ccvIZ+BiaMR3Uf9vF
P76xYMzgKWa9OpQHZfw/AhihICwLmNVbbusHms5lbQC3aWNytBlic5CKQb5jvcrW6+1W2pci6BQX
a6Bo3iga1bnKVYhu/gz178KKX5BekU+8h7g7qzYQqdtphWaKRae1f2KaSiJvUC+475Dux531PuYU
55rqCYtCPdJC8Cj2Ajz1Dp/PyWQhV+9qdYqxt6f9pHPsb8SCgan3aNGk6tTciGdFhxQhwmU6lo3h
FmzoxDHwKi4Nq58jLZhKuL4/Aqn6McvbwZ+Ul8oEgnbO/siGHmcaRhXvt/H5I7BR0el9t9KRRFhT
xtu3aJViYGiPp9qemEu40xDnuTissRzOxxYzq39VXf4sj/hsxsfN7ln6b9g4KhXEa2PIXdrbyI4b
1HVXWfH6NaS0fikzJiIESXvAcK8k9WKSVslnp2ZMUaLSCJm12OIZGtXORRUT0tsYb5dbVT4IRPyP
OZDhjxinnyvev/HU+q7ZgOqKvVii7rL6CID5cemYB+5cz8k0GASj6SkCxCUyA6URhNEm+JhavXk2
Pho+S3Mro8xZ7Dr9QumRzjwZIByMSgVzFmImZqG6v8M0vKr+mf5GWpYu+FJx8pP9hg2kBq6/S8o4
wNLLGOWe4poDt4n8OU1Chx21L3Iv+XMriGN8qAZucApmHM5BqwCLEtXkM+pt7ljgAfkGZbkCD+Mw
dl6fMZuGcZSYkLDybe53BpqR4bUD0sTWaG6icwbNZbUwwC32sGgku2omDdBG9ogBXhT5NgagNzUS
KA5IyYKEBSajYQwL7PjWslvDwzEarQEACpQ56mi9tql82U4bUI2T7mNpHyDpkDAr86k5LE/FhTh+
o4MZAwLpR03YcnXWOZHX9cyu35RBt4ciHdsZOpobH8GsesFZbXJ6YOqQm21rV8bP0aIEJX2D6Z7S
xNXb7/wkZqwObpSsxw0STV+Fbdm9LpHz7jIWz7tvLHI4n0FUU7eP9WaUAi7FNTOFDWa0eClIGgJ7
4AzWMotWdMkg0cvhJski4jxy2qHYeUvoXD9CkP0CdgGTrUJwDrW7l6tmv+PLL7c2IvSDVnJ1U00z
c/cdpuK/tISMXcjwRtfQoG1YG/3Ru39Mv0vy5nItgMB/hn0mnWSSngUgkzitxbwduHi1B0gWu+sq
V4qULhFdfRW5uqMbOw28/ySJBXFHx68CCEHJhT/x25idEMXc8iCW/j8B8oPG5p8SlZeN3uhCJXyg
3KroTfxXgOyH//3zH7alwcNyqHa4IyHm+lW8SoqVeED1Ttm+JOsZIEQig2IaemENRCXP+PKptCtg
jUb2v3AetbO5FNoRXpZIopNMwMaLpj4FisHhXWjErKRG16O4XwJXkllIthXDxWiBTexnc2jm1Ap0
m9iV0bOlaCZBxw28RSZWrtkZcXDcETbXCc6fKjuBHaveQVT1g5qmTK1SXxiyhVgzqY3CcQWFy7iV
mJQSuAvguHOgPDa72VdYWfpMwe/i5jvqpGNsBalJ0WpUnbsd7XzzCHaRNA26wGaF/5J3Niuv4XGh
SBCnFoUOpk7W/T1lU1DkmSM8/aYHJleeZizbx4TtIoFv0ywe1PNyBt0Yxas0DetmYaiNp3hff5FG
9U0XSaMM9A6gnYtLp5G9qQILudbJhWH1KOUtux3dS86NwRAqSQvKJTwXZJljhxn5RHWuiG4MpOSJ
n5VRkuNzC36DkFXPEMYyp3jnYsucTIP8sgqlVqjV3UEsKHPg68fGkEZiv76turA7F+RP9JTBdo/e
8hKt5hLEdDgA21ijEa3oeR7TOHRptSyvJVY/ILNeK/Y7D5Np4MWTUXkmJRuwgf9quK/Hr8Bd43Ac
PC45vGCZLd+AUGIHlq2AUJ1z7xhOaYjt5BKeMgX8vvdgcIa+hGCrI9Ck3RwVYh7RuVqcjw7+S/Q4
HbepF23fNOj0WyL/BDWumqH+NudAEgZxKhTNB/dpIr8u/F8NxWYznx/tP9wo9yaj9FzpZz+oEN9U
WB88SyAE2cr5AQW0xSrUxUq13Mgg/JHKVL5JpQy6KOv84nIGPMT3UBTLFCQ8cE1PEbp592zqeADP
NpkVC1biNW3hpVz5NMutyUX96zWONRZQK368zSKNNkzU2jB6zk0vgp6YrfpT9OhNASCSl6OrANrn
+zWkEUAA9oYJ3Me0+0DGnAijrbtrDYD8/FkhkxP8LtFoiudN0OMXMr31Ax6nnHMV4U8o9aR5F0aU
cXew9z42xzubfIcmrGwOvjSOxrNd2EqVFi9MQ+vQ4Mx0wo+kCLtBwg7NKdQ5u79UsiTWS+mIe76W
DdvBC21EkOL1AJ8rzfEkWHE/zlATNBl/FDtmjM1qp+S4At/XL/yy6vRic1tS998yOkP0Wb3YLx59
Vole2k4/n10DxZxvCZZskrsWpJGWgV9TxkSgMIaTahu96z5jURzqDkk4f1yriYMr2OC5+5hTioq0
Gkjxmx4EierDY0JKTXf7rbriRR8bC2lkgj7VQmSNY3NR/WvE+VppN3NS5VPM7exjgP7ZLRfVnVDT
VumXqpp08gDn2aTY2rEiKAD3z/ctUZH1KFb3o2hc9NjDRyFkbAabMZy8SOKp4+/n4TNtZzLKpLN3
BvXg1sfQ3DgGx5waDb9k4zO4gmWnfCsM1hLN3/AIL8diNOF/YZbmH2XJDzNQ2ADwMpJScEXBRRU6
HmuDSGYxcD+LxmywE/1Jpt7q61XZyGT/MdalH4ynwMkpog/abJSOZh1AfCCe4KQfUURJbpuolA4z
v5SJlLK2MHoeju0UpjLd8oeCqnO/LFAVPulmTcc+/6MdObmoy7uIQfnqxtsaZGzlx5priit++1l/
j2CzbZcYX8nPihbGrI1aoqasp1zNqpiOmX83ZD9/wXigaNr7p5VZBSylgMv4YylUs1kbQZr5Xj81
9QXrtU35+obk10kbuuIn2xZBg4a97KVafH8WUuNobqa7Z/d8Tj67tisD6X7OTCxFC/zEkH22TTYw
NfUZt6egQ+e6ccvMrsiE+RR9AbC3zRPFs8vx3SYszZJ7sQpBXlm3VUrAHlMYE0BOB5i+Th8ub4I5
nSxRp7gNDPpVocj7zA+cbVo/iPb4Ia0EnEYNqfU8RfgbB0vutz5Yt36HDVlfFdVVulsoRUqSqUuO
JAfNeKz0olaBA4oCGFUHzMCYOE4H2wHg2oj/9OzXt5XxCR9gDzwWaxPSMRRyVkBAMdiC6PEueXq7
tPlCjqk1BSGQu+LauHHv5Zfoe/CRAdnWkJG30mcSGXm/7c819eTePfK+L7QIp17oA4q0l4ryxJ3A
oDtJiqrN1tVPrO+xpeUZbBhiml/guiwCm1IZTzCNnLPsa5rPEWrrKwAnQbpmtEVwNw6QbMt/7TMy
9WjKOOXQkFrEtKP+KFRVusQLw0QLCjnqlD5iee4MZwDrIvTcMwMucwgIYa4++qssyvCX3URT/GoY
2adC89rqXyxaQUW2WffBf307p6+DoYBgXNYul1ImgNHcCI8Ezg7Z8VFYXK3AP70p5fwEfpj+/s0Y
4PNAnENp7SxPob/EUeX1XS7oSiIwNadOFdCDxGtjtsxajpunUSiCPTHRbz37jsBq8bMFZbEqiijw
dfJ966qhMYjhJjKX/DyWAJv55mMdJ5On1xiKffCxXSe/klexCxzxHREVa2EQgeUse7G/8/XECoM8
dGOAV85mSA1Lr+YjJM0SFt7yg9XOoZT1eQ3SaXt5aoMxE/2F/CZ9qwYDK0Lckf20SiklEkl+XHL7
FE5Ncl5WTEoOZmULV8DgDswgJFIfOfvcJjn3UV7Gdy+e5F0RiinmNv8BIM6GuCe+Y4GcqJxzMmEF
Q1f4iuizExzqrrbWsJAm9l16xecJ3EJMakEDK/kOucAtLjF3O2WMeKmguD+aULXJw1srAhjLD9gH
mytNOQz/zrAq+KdnyugDYLOsxMwPaaY4emr/Mab3RrxV5oN4vg4KfDvPu7aUdUD0b0dbu34NbmkF
YwlBY2Olz3yEu5rJCq6MD0AzwCjZ5emb7gmeK2L85MEKhD5aMYPaq9oeDIKQoVPmbJm9EAO8mRjb
R/4/PP5bgWS2aHHUdbCKwnhTCQZeq71fViJR9JWS5Q3JID74bmKCIVRuYyMmahSkmucgInEQoHUT
laoFYaozCrCTLX+VRMRVuFLLBZIBO+0S++UNCM7R9AapXTmLYloKvCyFovLTjFz6MKnFcbp9FcUO
+jYf+4qhwPRGHred/Q0wBYBh8CHwQvqu3pAz5zbZKntm5ar3yifjoPJnjj0c7PG+e3BHsBVeqmqk
yolh70Lb7wRSmuphNsVXhZpS3K4l17BlDOqdMIt/xYTD06hsvkm833VrC1mnAhYnNVQU26lIx9vW
KQix1N3OG7OJ25dKQwrtmuGrnDG/PH2G6ngROxbWhL8B7UV7i/Uz6q+1mfp+qG7rVTXwbnAJh3/6
47cxfpRhsMkn9XaweEAMe2P3BPk9UZH0bjLaPnf+u9GSRAdDgwKDxD3p9q2AIEqibb/XMfiBb0M4
vrZgMwNUPHFz2GjuHsoX3Xagg1DIfeADQz1z87xjPQb4fnwfBCsaaLuBywyfOZRg+fPVb8Z9BSRE
w34C3vJ4R2j5OVe8nFsyOeTlYEOE0lUJWBx3ofDWxY0cjJX/wz8tj8rcnvBbmaKwMlsOwyebB6Jd
16zbQmVrKYEhtcZhNLJSLUD2k0Vt78BsRnWMMbhUZSRidVaJXuv1EiqacViqCAvnsBZ2cV6ejeCW
/mLGYb2l2jC9SIeCLieagyJeKUaS0nxlYXoKcWghnhAsJdnWJh1Q4wuW2v1Tl3Djz+Zf96Y6rT4y
Rf0RcqpKcAJ3VfL1xiwaRi+WI5vF9wgCfAWMKbWGLoQYxihv4XL9/MikeCk0NHiIK9HI74s3ReTX
uUQdnamt/u5J1E09m7BKEgl/8rrTiaQ82NQdbT6iG/o7+oD4p+Xfet5iRqYsyCfA8J3zYERGd8UD
YTmuyDwHyeIXLiOmkcHntZGzPXMvj2Leq3vnmGp6xUmut82ukdYEUUqMQAKESXP2aELzEY33P9RC
Ig4SREMHD55NsyEU3xIN9zaVkZk9jijRczmNCQLYuAOYkxVbpFLe3wFRPVVimdGVgEOF+zlwwnJk
OEqPrEIM4Yu+rZpUV6tCfSXHTu0XETJeGHjz+lR9FtndR/bi+GRwfA22rxsCQoQyOzSnSAyiFlgf
Bp6tv57UWCnIY4CH7/+Iu5h6a4KQCbczyQ69EBQFnb3Nrs1OfuuuKYb1QnaDawjwvtIERdz3RzL1
fzxmsBYCWqwHBhTjvP3vBIsBBYPux5ikAzrhYFe8F06qLeD9k9mgRzvBAOuEpEZZOXOPKRG4fryq
tG3L/i9/3jDn2IGyiAYCS0iuyiUXFsOQs+xNYkJSjDy5QnJ3Xcp/l0Q67VntcLPVy1vIjpCtJ7Tm
In9w443dmRpCgYT+zUFv5lZJJErQAs7HagCnB4gC+mIuqo1MzznfLpxJhrKNSou6GK2e5F8wGvt7
pUKcqoNxeztI95ex2U8QggvtOeNDaWSixxANqUu5me/S3l01vnJQKhjptOgmBvgScHFi4tsxErrW
kr60so5pugmu5oUTdFGQd6OaYMH6kVOha1gQPfqACEakc8dWWQrE6IRANds2bDMfN3yAzQuN5TcK
Lo6OOREDdJuTBO6EPXVZCrZh5G3NJqSOeYx0vqeS8i/MLVVDMOQSld1vT6NAFiIPXGkB7RIi8dbX
C2u2LetgHeZEFOrrIbMOjUGtAbnTDTLpNi9yHWviIKbfgBGYYa7r+N/S8vd1l0LeqPZCrgLgS1RC
u8JT9YSl8dP101o7kT5w3+O6vkRg9EYXM/NEzoRY0HuB7oB6I6H9TcLAcaqxCB40N1ODTswO2l+R
6bLY5SUzvFOZIj82ogqXyd/GEasUOs+tSDCMetg5jrBNUOZAfWTQBTQon7xOZt+E3kF8YqA/YSSX
UPziRutpTNx0OVBWev7ZZSwjELpA5unX3qU79dwtklUJxO7XxxPoSPgDF5NL9PnQlHknb8JH3/XW
V9O/iCha/kjKzTRmYZN2CHKC0H0c4RnxpR8GsC3tD7er8muONxI9SLK7xoNNoahDXAIAQ6BRoCSK
jEyBC2bVq8Do8dphDhWSub8Sekk1n+aIlPye/TO2Tqbh6H9POKhkkb6i7lVoyVWXhov0PXvTJYdN
WxYq3NuretX+Qw+bLsgayEgZae8fTHcbxXRm+7afmLUEHOkaBdhYgex1R+IIWZHZTag8a5mwKNFz
v4I2UiMoritpk4KRP4aDNpsHAx2iWPKsUkmFHz+7TKaxUUzu2scDflcN0vNzJi4Kz11EsYmUBmL8
rjpfFCXevFxkbx6phF3bzaJvM4R921zcK/iZXZPPd7fdnLJ39TJeV3LpnnXgtr7WqWVS1/x01/0j
FFbKqvqBvpUrBFX2e1OEp90ZFJqv8HyPmgQx30InQoilQXXNCyScgNuP98O79FsjXuYIp3a1CGty
lscjssv51cz8pNKPXQRnI9bZ35rkj58cXwyc/zxkogwk5Z+lvZYAzgdkT/pKBzC8SNn/Y1EOsMj4
oRNJOfbqLr5RctoG5PD7EsshnKfr1kpd00zmK5XI1HzTgNk/dm4IEO4OXTpb/X/kEHHHPpzZg5X/
aCIWQVL6ZBLGScwEaGI73hJolLDzKkA4tjcTMyS/dtnGNIREkmS8v5+/gvOwDSsEP3MRBhgbik8n
f1OT1ObTaSnw2Olls0K0jJKm3g1agpXxDCJ/ulHoQwpedCzFf5K7mTMAx8oB/xRL/wQYfT8Cg2k7
44lTt6IRBAGZmCyIy6yTL0YF8DHiMmQwtBv1Z0qWYojBTnBBvC2RRqKOcDPqxZyn4+tHjcojoOy+
wQeXNJaCo5R+rMMj4/Pk4Tyrkp1S0LTCeN2Y1FjA0NtADX5nMEMjokEqxTk/yi4O3O0/Ce/nBvbt
DFHpmAfEsAIHWXY5NaGrGAyJlTG+GnZHMQ55kEqQLQHrOYeMIwJoF8jpEUZYYmiNAz8aIuPpe51E
XmxJPMioQaaJ0e0nfT8sAZD1D+NEuluKPuYKg1yP6r6RrkvGkd/JNCNE0mjl99ShkwFbwPJex/sT
dZtBvji3rUC4mKJdbK+BhmMN34LR0NdabZYWT9rkt7QwF1P3z1J7NTdiYeD464lcovWnqqxQ8JPm
bgNlZz+U80ixBMT5hRwWL4o0iBGcLzAzZsMYYdNzXJLo+r3sP1pzozsytnQIQbZvDfxlQv4t/qPF
JCLSfqi6OPQMESOaRAe5+cPAk+5K15pUEbeqG8cKzzET3POnqVRHkMlH7XEUiLTl6MuKBnB9bTRk
x4DgeeUGX29n6d8AREmfqtqK9Uo3b37JIG+3Wm1xv7ynfggsjxPDKCqaecbiohWeMuBJ4eDQ92/y
rv1SucGwpfN+d3bq9MFHLLCHmD87vXDpppbE5rXCL9mZAmYOp5IIPJziMhpL6T40gAUFFXWXlSnv
DykOiN/k5FIXXYjw3q0yi+OiAw0yOhOJG1fM/Bl/wXwvfwMzvuMNIRU/JrIryH7xg82Mrylxav42
BIUmomTYSKBDnXMohuUebuHsu2qSq2rXkXj4lM8T5lx3S+10m4e+74oQ2AIz1OZLCFzu49u4yYgM
Ft48CByudJfUWR3qvVBh1ixcnCILzSwr73+9/B0RjPlTpF1HR4bNedH/B4MA/56Su5V+j4AhCx9X
bzsFU0PtqCA8egj+j/hwDT4aW8ZUgmWhr+0rtz4t/H/mX/eQ510+QW4PJYkDMj4+o1sgAhRLsN15
UB7puQW5jne3VyJln10539TSUtXigdPmGWZkC2teVMwB2kEWThzYy2b3cBUbZ+RpXjaAs6c6Fkch
xYZXscrlttJYVFMbK52Nl2jcCDJ5c2gq6+mPyBMhkfwSpvXZqamDmwtWzXK8qRUE6RfQwIhtzMBF
zZyvx2RJrgiJFPptsSMkUuAk4xcwEDWaCDu5UCz1esD1pn8KHgRHQwxoxLc/zPZCgbCAqAdTUDP1
6Y1p6uESA/2OcdA6ShN20xQISytWbAb5uURV+8qL9J0nmgS0HNPDmgtkeRM7ZlFvFsU41fBOa6x8
p3JHxa2LIbRU7Lm6SRZGr2fW+MPfv0jvatpAQVOvJqBa0N3AZFfrDKnXTb535aWfTDo8jOKBai+b
Nm5NaU4BTF94d4oL1e90OG25X4GXYvMFSyC6ADXNGOi313EuuuCrK/RXy6NT0ZbiZzkDfT1cb8hg
X8E5rSXW4nStgFrs10iKoo7kKUxsr//ttL+qJslnzNEd6GLPW7CqlXL+7elUPG9sS7RqEcBRc4dV
aOfQvJ2wuxvN2nVllAoM/1eSc/8hSVg/d4zypB1g84bEX5L0+iu6cZ+slkgQVboZRYOXGg/rgvxY
E9vjCzoVeaR0mxubeaxBFjDJpYCy3weW00pGXihZ77KxHqwpPzyM4dTHAhurmGgHyH9SrE5Kl9rZ
yEgUEDhn6tbq7/GFJ0Tlqg6/jDuvy8tHxAMBHVuVrnTINuR2O4zDc9YMGf910iOuBx9twYkGMTD+
sMndqO7kstjxXVO6bEaG+eeLY+DZk9At4VtKVd0IXZWiY3IZK6/05asPvVwW4XQRcLAnlsEZppjA
YBcM51DOBLGoqHjrbsNVA5a3Li0fHBAicPzhFGcbWvfzZ5qQxo42q+rvH8fiQ/tLo62WxYKrR4hc
h1FFEwoJ7/4GE7Of4W6Xz+0MyyEx99dLnDia0KZdOOI4zvbKZ05SZ2uUOPEDHTrKSHf3jEV2zAzk
zFA55NVGxJ96iL42T5WbI3k7g09ZS2jjpwqEQ/il2orhy1vVY32D11HFUrEcEDPP23cy6DwYVxnI
SvVYtvUri/mfQ5VMb2PBsfOQIe+C4Gcgx9LE1YZbxMhM0F1M+FM8NO5uKDHAeT5YiDi2UpUx7Arf
C1GQWgE+NHp+h1SZvNy8hpIKfKH8GLVKskV5BUdBXGDZJLcoH17BYfOkGsCUOGUBzmVxGVuJaJ1Z
/0GURHai/aMJOMJdEh2TVhAInyNydXYNRlJtrpnEz0D2qpFxG3c72jMH0ad9+v/SarM/GeG7d9Mc
XjqJAJNfGUqYwLv7gErl7tgRf2KmyR0zXmYViFGGpk5gu05Qn2Is79WEJ0uxgrjuCVubzUVMqTEj
0WkSfpEvRVP7hvrp/PvQ73pGlvPrSeqTkFevj5GXgPksRV4+FIQg0faf0rB+n38+SGsKwIXEqelK
s4Dmh/bJQSr/74rPOuNUc1FDETJL5DOTJVh8ctyjMc3BCGjxK8p+UeKATdXcsl77/S2grRG5JLpZ
lbJYfW8BfSwiPHE/bvn5pO+11Gi6dZd2tlYSmVmjQK8JJrR/wLsPYfJUUfTTyx8CAShkZKgJIbMk
hNrnWNX6+eDdqxyppB0Yp7XKhk0qcQzJbnb2pTRoVrAvGw3WregrhZQdkLyvFkvjbMW+BspRAhiL
/Jd3taL/dQ0VdVNdRdsg9hVl3eIxS9mMLgx13jjprBE2VlL02FA0K//rDz3SyweNRjNcKD0owngm
UyEZNDYIkRFAhIV/EFUpukz3VujHoOznZ5eHKTJeeo09lyV0rn3+hP21Xm9q6C2hcvTWD0V6euuB
2zkB1vn/l/osCg6nw5WD2AHombAdMvDMXr/ietmn6A8P4Xh2On1nRSo1pTSjaRTbvI28BR8/+P99
5OmP0UWaLA/5qZ/EtLzHTiqKr0raubQCAIxi+/eq0NVmUXoT3HKy9i4nw/WKX91UkqZeb00RR8Iv
sf5823NGNLfrKTNhY2YtvnmSM0KFnT5tmHqKfcNUJ1TP/iJ19b8VI69qgz3PduvcPvFKji+0Ytns
mOZDFuluFb2dCiAV3kw9KBB/CfFjy3MHeScG1SXYkGwL3hAvAEODUqx0rkRUnxtNx05l4L5MgTCm
5mC4m8eO64ZjIIZf49jghG1kruIKEVjx4SoWy2xy2/nXcrqjJhuqyIrTTL37S4MBPDGY3LztRRno
3TnlA1uUURmwTc0y3foVTXT0wW9RZjK3Ehx/Q0BbZjZwU/Z61LVMh3ZI/UQbno2TczsnRRVeWpM9
qYY/bX0vMCBHXD0hGwXpecBFjYWR24R73+k31YzIP3bepVT97PmATV+0PHUqSAkxhx31ovEjmrSG
8qGPsRh7RRXimsnZE/+WiExGWkcHijnyIvJe7FmLoO/R3YXOms5x4sgcFXfPv5DR5ja+GnADBOWG
tHUGsiPjNCdPfK+RRHTZ7Y/ws7A9uyXj0GrCZB1sjthA0pFyQ6cLbEgU1FpOXeOqmFjjgHIY9PIW
P3BCzLU7DEkrjPwNDNEmFbheWb9YKoV5wTF5HVOgXe82wukWZAgX1DDFaGEVT4UZEvCoR0P5HqaG
J7qdkbqYACC4FWO/IAS8uHG7s3PsDSi4lAoZ3XniuXMlw+UDhif/h9MnjcHsZcjewx5cY8s6/YVI
y9zjbhapmCLsaEAGfqW+tK1Ha3x87mZ5rdJwaSJFypRhHGwnpj8qZMd7EFXuZ7jhgGPanr7zo4No
EvuGrMjfySoANq5ndiUz35DPPnGRRAu5kg0t1mPtzsC906lGZhdv4G1Uo0DyrqySqCuemexpcO5/
My28RdSnV0B31XjIJUFisJugglNj9/EezMblytEdvyB9crVJnD3JdqmH+3zk+LFDy1ndsphXGZOw
xIDfWG9bCbbEmpbF6IRK7XKoJM1lYkVqNVzLDfn1eGwG8FnJhNynvkmFFu679f33w5/rMXkAGYIU
F5NTOfiWNdSyGj1KQAD3pDElk0vPUSpZseWefNAikelS5MrC1g+lYAW5J+VCt0O4/Tlc65ED/d93
ea4Sl8M8uqGkmYR48FE7hW0JjIq/DXlVPAqU2KDeWqJBqsHhOuZaK/snhOLqsMXJMGRexbAqKE5x
dMXK2x/BcrufGf5lJNUbNLTfKYjZ3NXt5E+ou254OGrg1l/DaUd1ojuYyCD+Bp5p38ZPvCX5wTaf
BBlxwpS1fmgNfW0XzPSSKft2sQ0Idfea8wwJ4T0Bk9M/OerxFj2uh0qJdIPc4f6XJvMr/SJjicii
2P0aC7g/PfV9BsqbDFvJVFYpR9HkSve7KIrMwKPO/AvK68XetJ1e7389twNuusZ4NL8d+bp6mAJX
GhE+4BFE1G6AApqSS4vsqYrIHIM3wzmV6l0E8zPcRxpUGD3gW3hZafKnSGxl8yQ+0pQ0XyTFJjjQ
doB9cVrL0fck3+WyP3D/bjNS/EQ/JYr6mCt65Vbw2ie8HIl5iKQ+Y67RwdY4ih1NZOLAWtlik3uQ
HHv6N7Jox/hD2FCWEr9QHn9DEdPKsMfwADdi4rh0vAHdniRPu1gqmG+NvOS2odnO9Q8+4K9Mo63H
jy+Bcqxjxv80qS6Y6xDi/604HLbZoGAXQvZVD8f7gv2Ps2iPw10XnUwGyi8SxjkSHiNQ4Rqypf+S
4wQ42x+3b+F/6vuZHDO9VsprAd7eHZMDLteiyWR5SzO6qIDs1dIsVrf9kucqaOXjfmk6lWB6+WUe
Y0zl11dc49RlluxXcWPm249Pfl6WDrwOo8YlQd+CS+sA0SVb/UUFwGftNqDnLt0RiyEtIpM5iy4u
iz3KoB7iWgoHzW2ZQ5EN8Ld7oqq+KC2KFwVbgK3p4bIym0PBKqbOsL2rOhvf/xPDN5FqYDEt30WI
VSXdlMH77JrWJOTbn67D60aSTLliRPMI3SMWMXgzRGWGFabvldYjpXWjbyrAUpOxusUu2ok453Qa
vygl0amhhLKAcGoSY5LgP1ox6B8kJsx6aplsGsSCmZYsk3TtOLAhUe+jsCo5wFXehu58Jr7Sp7Tu
WLuclXOt3eVNEzO38HnJiZtL/2mi1v7Bgbpn9HkfsTq3i+eJLotaGAvIg7DeZYP/OyNoJbHeatid
Ra9RZ86T+mxoSzWWebEjqQJ7xCMh4CWp5GlTe42aDB1jvLOtTeIS3llyU1qNd7tHr54u7WCCsTPt
BywBfeb5VA0tymQSHmO9sIYDMm7yZv4UNxz/Xy9dEPv/69sh7jbiSaYWv5RX13tUZ+E7DdDz918M
NYXRGfVYr/wY8T0NS7kcxqEApJQ4mhzyiiYyPGSmjFGqjRcqpS1iCNe+NTdOKJlaPfertjmXR2cr
i9c/dKELTS8AVoJxnUS8B8JfbG0zryTbODuczBpyBqgMacT1xSvPC5qII7R0gFnc6/tQxl/xkTq1
XQ5nbGqswk1VQGSButSA83+l+PXv0qEoJhZCHVMrwOlrpsCRIvw9gf3ErAw6+dBaLrLXPvFCCNEu
JFrQWnk/rAc6WfoHgn1UX5D0CxVeuMST7QIPcWgFwHRjJmbtR11SfAGX9cFZr5KneuWsYeC+DPRy
QBEOc54THwneJ39kn8p7qg6vfgMeZrLrs5ojQLRlrYM0uRO+9yDNxM9g7+GLDubNmCefIMHWf800
WuQj+d6KEdaeGrjy3Jvu+ho9OIopaV38nGJe9tzuM5TbCRT3Oac9mW476jS00E7g++n1uRmzH3oS
a4ib1ATT8VIc1+90D9G7l7ymeX51iJ7AEHV7DhXRdDOPZb5L9CKdGsgefqZ3ORcY2tPOWtXoiuKB
dzT3OxsjyBHwf94NZLcK/XicEBUrZQVy+8wuuui1QFs3YHDhEtdRAb7mcMq/j3l3hwvj2VrsNnsI
DYMT/0ywtlLn0xc7iLf41unhQ/OxYDj5DUleSZ0Vq3U7XE9GkYV3I0SzGKjQIUsgfqN6cSMda/HN
bcYq7+zq3jCWjHly9tl7ZpAgH/ZqBwTfB0dWkhVgm4WYmEaAx5xUnOhsqn2BA0mEY5+ztc+G0CMX
cAHtk7w284/NtbtVQvPcw9gu3AK0tjTJi/aMPuIiyfzZNpss2tPbJSJQhXblpqUWMTmNMJ5Vhvep
3IBl5V/WIb2DcGVJuKXl9nQfjFy/1JekCOcq3kwmhT8Xa+VNQIFJff/DcpVmJcjLIndaTfTaBhl1
MbDCkFFt+b7u52AAVLxGd2aKact/+NV+MmlBEGCuJzURAbFowKAnLalWzgXIWNZtm5uH5jqWPV9Q
t9C/syqZPveRigKG/Cfz1o18CwCqu1I7VTg68IU8s2KUSZMCAKxcjBxeXXjhsA5q+bb2p96ZohGn
jj0uNI2YXWqTgmmkExiCK6UnzDBUVJ9J2K0OIpFMg19Th/D1l3j13c18hWJ1vCp9YwOAFtMI7mYg
gahPRAKdm9MAHimuo90B3ilLg1ORfHLYEuSmAI3VuU31IQW7+ZTPXgSDKN7LzQBEEKJAWvIqP/h6
47TeOsphjJAM9iHOgMry7TakfUhMOhfcwYxq7d6jqzvYjXcrZb1xsAsq0nwuSToBvbeqTs01U27j
+Bh58NjO1GUkJ/8h0lDAv6fHAhv6Gb8Za0ah2hq1NjXF7emNCN5VgPQV+W0UXSLePkvXwR6nm/lh
lCHE4eJTDH7fo8gPJCMxPqHdtHRJw0NwFGUJaIM3D6MbjxOkQfSc9AeM9qWYFruQvqBmBxmMrcza
0sTHjERlCV2bb9Ev8oDl9QvC5GOATM6gPG02hmjBKv2zfedW3xqVroNUzcAOgtXLDaxNvw76QGmJ
UCmqEAIlDrbriKRTuzw9ugVOU567eIuVZq200kVsttuR9krrND6YfyJc5n778SkhKl9pC8SEq9Go
V4cKm/EhgQeZGmGxAuKcqwSYkk6YYDzIC1vo2em8AIwgu7VNSDhIcij45Ukzo8OiFVaLpOsHyKsi
uMGWvZF8dhb6f0Eox7CtCn+14Lc5fbzZ5ap0aJvID2DhqJpeCkY5VBnQk2lr7nHGwX3wpER1kkHL
HSWZKdS8dXa+mp3OCxiji1DE+b4IjZRBKplyH04ku8rWitHf/ReKlIrQxXzGOtp5JbjGqsnp14jS
3fsNcZ8tXHicBcqUClYiiuXmmuQSOEYK6dvlTXAZ8OjAHKj47+4XNOtVSi0HxpMGjC5E1WvmG9lE
1srkPrc/fpuZIJ0itcmDGGrx0hEySNPdPKWocUeKkyO0truxwhg390w0T+S2pMfDC5nrxTyS+ZKQ
rG+bu9gBXYu6PJEszNlP623g7AmTvVKQpZr9iv/6mEeLnNumXO7UWDT6BCtzyrIun44L4NTEfL18
kJcNereENzz7B2eO/Qrrc0CHAOMlC3GiR5s11nfDoL6FuiM63XxmqKdm4CIGDiWpnU9wQz/8/xwU
OsEddgOdeHqMadU7l8M+/isukX7DqE69UQzhZmLxMNLEAppOfBsChrAudBaSoHHssg4RHG2Xq1Er
WvEoXUUUQhp980OXxxEqtNbmuI4uCj1r0chHltnBislD3wpBiRvNFurju4+EeBIibjbBiq6P631M
kDZ7jQvO/F3US2DbpNvgpG0IQm+hL8sXNZhOJhzHRJ0JPIju2XP8XM15hCKA9ZWywSta0Fa8JKUl
eF1NxBob07pd6xE2PHKJaztRf8TV0UGZft78emAU31N2QqizSTU0ADx7LPVZMJs4Xsmc5gsDRn1M
K2TqCVl4Yhpuk3F6DZfnJQHvpHYaZdQACM12ahoZ+P+3r8gvn5MnY0ZK+RgprCQ8knw7rtu6vFh+
PMfWnjHj1vLTFNnIkdlqizTWXedkNwrkVkNvkShrhGed9YvqDbEH0+2DlLBfwA76QRPbpBk7BoVB
OpQbXaT3qv2KQE20jaME8nuMQXawn4PxaSCI+aHh3yJNxcHY+s4zoFyvE1ugo8ty8nQGOkXi2MZq
Ad7bwXqlBguq10dA9Ixkxgb/OYBc3WqsXBNDGpY9Nnzlti9wb+sC/IFV5gU5Z2H7DzQl61/4JPIA
1uPkgk7oL4EORtQQFRkUOKkHwyL3lzltNVqHTBYwRIiBI8xQcg4ID7mYEoTvDyeMcRDzdLWIaHev
45QuO7w5hSWYu2ZN1VDOGU5v7/8G2QO6NIOCx20Oi84AeiSfT+W/GftDphOdTML+BbBp22lWc6W5
o8RET14RLUKBCFnE5wGHlGYGIFep8reMNZR7hfTfUKENKKKMfSQYBl6GhxEwoEr3v193hS3JJrvx
mIdJ/PiTfDoeN+BCpmZTZWdFhlS9p4Mi3ViwnCXByh6RINqDCzxgB7YZycR6MMP++rtoz6yYB1AV
taLspTFHAHLHdV8zUxIVhgY7ImHEPa18uBxEs5fLBeEY5Laznq9aAFVSfYIhVOvHZ5GKG+fDJsfF
WoxzAV23D4fdP9/ggNVL8MBGYH4jRTxy/OmwfuYawjNyWse5eeinodlfvl4cpQKkOm9Adt8GMSeV
kpbx7AmEwbWpS5TUzI8W0bine7T0ty3h1Qjk6ZjdIBxXv+Y4hN2RwUgbsHO3zTISbXX0Qy6F2AW9
Pzfi4Arn41BdfSTGXbcq3ZZcK9z05Po9aaXeogC41KraPbuIF7R31ITYFu5ZALDFrL+hLQ05/M5w
jXCbVLGYOYdbolT8P7/bcug4/tBf2gdW2oktcmCcoVkGrTCp/5Ph4QyWGqhQruTEl7krJ09BM9qH
RZCGOPZjP4k0ypVCTS0b5sCN9SsWfbEylQO1rpXVJWGKheIqPjwnwJ9gEDEeroTgwHsMLmNHrUYt
aU8S0D+QL7+tkJhwchYcJS6KXcZPsbZfcsQnVyz1wWpYA3f342WdgL9dT2ELfZ17GEnD7cfcCNOi
/Ee1yLtulcJy6+TZKRupzKzRzB941f9Vqk+txGSeMDi+twXMqajVhyb7AF5HNLNTm5tqkwnyxIVC
+0nSSZyk12ULl+9Syulg3RpgkXkT8KbKbpUvGttNBNonewjmfOjswF9ef6hgwlKhPuslrL1pwZPS
WlEmdJzg8w4FxUkwbcwZRhLtfuBIk617lX6bTr8F0IptnBmCY/LfnoD49CVrWz+hTNV6tiStOb03
uKdYBe4Uzi0ija3xlZqWA6EZfa74/KHk13hqg4L29Rwk0QsipB6q6YhPXkKw2C+Zwkkhyps8x2q5
SjRafTUQVt93VgNsHTYuVsmqsj39/QSRFUNTg7XsMPnJrrrGIiDmH0O2UHnbARTt/ODvWCSRzoDu
8okZk0dRUBJC8JCSBVkvf9udX8ocNpv/Jw6fS4aW7XVQl4deUr/AKmL2brCqPpTC5kD2GlOpu8Q+
fNuidcMlFu9MVsW3YvMbu0hcsR9yqGLAb9OEMdP3nmb+vD7KRydAJLO1DJQhxKJEC2wDCWnmQFLd
ljUBVJOeb5bOaCAXZsVINi+qvyuUQay/tHK44OIaF5wQ7nkLjgg+WhhS6B3w68yZnCfzSwAWaamk
LLVw0PIfZHSCIz4zZf+T77QCf13WXPKldNrH5P7xGKjH9JXGzBPiJZlLRWixJanWn3U/TwCytAeR
QqHFQ/2keyjQp2jpUU6AU94/K23+r441WV9f9J/FCaZpawGBuxldU2g1ZHg3jV4mGNV4z4PEo1rI
RWGp1Y0O4/haSFTzymnID0Pg9omjh/ixWZfVfe09fHDPxkAcYv80pvYidVZ1u8waU8+QHVV2i7ia
0xiQuAptkL3nhQ/ReVU4RrolMEVKbgLKa4EplZjAXZsMK5Vts2lL1DKZMu2Efzqn2d40OjqR6hg6
nQ2AXiBGk/QFhs+0Uo1qsvanVVzVIaQvK5c/EtmSxCY2YfUTzACUtC30ZDiiRn8HZjFv5E7lj2vh
m/c4EF1E5nQCltbb9ynHrVBBlFfFbfXxkHYWZ2hgiuYzvhzvMMf5Acym50GK2MVf1p63VjOMcuq6
IoFwpZk43uY6m3DazQ9yYjM/A6RGmez9oN8AAD1hoBekhradGs/TAhXUUmuogrwYRmYOmQ+zgzFE
o9SIF5Tu1J1sIGH+GrCB/6WoMRCvZObmqTz9DjSJqaofg9/Wrik2OVN4Yt0wCepyKOEYzMC/MWuF
B1l6mMXU6Jl6iUxRRapEn571+m0LbzYeTM4qLy30llwcAwjc7ooQgcqs/11FHgBYOQjTXK/dDBAR
e36LiIjNHCmf9bx9ZbquhKQnc67EmyAnjA391SZIfinp3AMlxetjQ4ia1L0kWFDEFNuNhYhvl3Jg
jGNGs56qeULwXw55UXrfMUx4u/OPMgQda3mcACaFQfQYgHYifUXGYq3OmZ52KCsEw8aP5HihPCjq
pIxxNnUNWXPfH0YtmHkqPAQuNzENsjINRqtrOVPa9yy/WknlpY4Upqes+776xUecerAGLVgF3/sF
gF309aiV02k8jvLVdFL5nvDD6meSpNwaJabqzVzUoHwKfkdVa2y1eqrwo+Pt+UomKK4qUEX9/feL
500Bg2lJMRNs3CiWxQHKg3jl7AonBCavrOWrYz06yL8v2EzstlvnOF1VLQDWG2Iwxh4VKnoAh/2A
8cYRuxtvz+m+3NvEhTBNWn4hnfZ4KEnD8a1mTNAuHJ25OfyoRUsC6wiL2FuJ5u2/wUF/CVZktjIj
hcqprzTSLxG0BMpveXKQJnYESi0Tu/YocqoxUYTf74PLBxT5+mF+C1rSgMSuFWYaPk8wmcylfuAc
jE8HS8BkowrLhKyAobengMwYQx70OkjApPijNT4lYFtKb3Vs0gU1sY4jqaH69LzZFq+3XCbSJRqW
3Al2Nv3Aa+DEIdlGi0oGg8vbRX/Fnou7m3kLhAKNzg8bLjUhE6lvG4PGdLaL/I8/LKL3SpGM7v+8
qLI8aM5FaVTlvov2Yzjkv8VMQrLhCGxb8ZwcMhyoCfUtD1j5MQTXdzitsKRRoLclA7BlmZd7MaZ9
KZqbuaS8zIrv441ROetBGnP8aUXyRw/DpAjK93rKMFfbMi0cU2HgNIpdNRruYZxvgCAN5tfnYA7X
QsWcZH1rT2LsDCOi8h+BGyyK/ClW/iuFvlpcsNaO+4Jhq3ku+sjnePwjqdQfnuBaXbG6tO56LQiH
n4cIlLqbmI2RbEE8DeC8lgu7brcMSlLxcy8dcgH/pTl2HxhCnBJumuInoHzFT9UOBG5bOGovwwVP
OLlOtV7V91jzJRcTTlhA2zgIRap4SAUt0pzZh8V+7xAFrfgRu/uXekFto2eMhPySfSTZhUgtqpVj
VXpFSWoOF3nBqc7MTA7OQT0N1BIaiTtE0or5i/coOxZha/bvhrWWpJfnlC7Lmq7imPZUIkF6ozsb
+EAN0ZwrK9iqhXnIlzWpFtU6+N3uIFYOqzELTW3zCOF6g0vxSTAVzPHUihiC+NGA3dg+6M7cPmt5
luzLteYPvgzgHyvrOocyNwsgNZ5phRdeOZjXhXSNwWCFFZOGZcHD2D7mKlHISjsKTLu/ww6sVIpa
l6RLoMCpMq657yOeRF4cjt4ks2iWH1DIIK6IFd5K5PB6oZi58kAZzaFah6FFyuzAFVpgnLTajhZs
66F8F4J6yWnVF/JSoFENPA1Fz/oLs295gCSSvilLIyCeUexEIwSpWMNbCg7ig3tm4Lh0qSWYeyrb
yjDtd7Y/SI1gWvQMorcrx2RxXeTDnJfwQDQgohXMua3N0LDcoQRwRG77eBQ7sDcAraUilL6D4u61
XDfO8O0tpajY5PHdoRKZ8vZeG9dsSH+P7LuZn7BIsIhWQcy5lH6QsGeOyOFBkw7Vw58f34OobbWZ
xYaICc0nXvIdtH353YVStc4JeGGYyumOXinK36lVdzYr/Yq4jxvf4LVwOTX4iQmh2+e+vNfmPxV0
FoSlcxQp2r5YHCrbq/CjIyuoNF2Qr52NGdVCLuQ61+6CYAjiaMfukd2WAehaPIjtaAaD22v8tjEx
wcuhw3kpYg20lNE7Qk2qYLxvEBfU+mX4+Ua51R5mvjBP4fWGg6wLyoEu+KnEYwaK/lgiZI6L5gHl
MhpBZeeF7g59hDsmuQcAEcYn8pfz1UuPTWwkFe+vpNLw+ZP0/zDVa0Eq2ZPxBYN15CBI66nTaWic
iNigkuhJlPgWy4gdThsHY3siJwvdcpipgsx/3Pd9Oxxkqg72g+BOKLP8BjRE91UXFCFRyoLVUjSf
25ujvFSKbYgNymgMf1OWMlicNMGGrVTKvtmWNVDdNVPVZOQeOkkc4h0YcRWDWHefkyiIF08ATQ/N
2Temth7N1QtQG+m5Rrn6wXmJGR3YoJwhMVhU+ZmJvd0jVRnjpW1Rwhfrp4V0+zwBbNPBbXwIn3uP
CIzPex6wwsjbiJXRnuOTkuO/2iOfgR76qHPPLrHv0vKAh+gICRH3hO0s2UWmDQwBfpPCpNtKOWIF
lbcJPANGD5OLpLpK+DRREzhHgzSLa/c6tfd1YaaDxFCft/BZW1qZkLKUy6ZvNWQHlOPHFB/veIIF
XuBzjFRrNYuhxsNVYjqELNRTD1lBJfE0sTiHYGjwphr1aTJIjZir56S2OSFBQSj2Cm0LutQLxSW9
jYaoF759aEHNKS+E9YSRjbVO/Q3Ph55+lmC7a6zRvwawNSmalN/7nXZ3N3c7VVOaEgVMHC7kbJyE
aTbgTNl5g1GWTMwI5yUAuFitOoOxWZg47mgkIxFavkKHO97qCKfTzwwB4SjdIbYEwPS8nN056B6K
7xDBOl2omTX+cCIDmlcGuQ8QQTPjTH2JOm4Yg0Lldq+hc7JxSAqOeLopL+MRbldpQJQ8WGfc2sVu
eqrgIVIVp/OrJtIjMug0kY2ieN9nfGZKc2QC4RL0ovYMCTT7TRlm4EvKu61A99/OF73sC8KogfF0
qREMeVGeBHLgV+J5Hl17vDrtBpHm54KPf6gwLZZCdnqIBZyj3u62YyCfl+22i5fKtCB+K7RkSEzs
tlw1Xk6hKisHTmIdNwSKmh0eSn5mxDeN1fs10Kk+yohaJamSCwEG4BR+EEFLZ3DxNEp2eg6CQagN
8rJqVPQonH7zK6PaaUydmyPUH8DG2yyXi1PafljUUCYUJLfnAzOSWVEh2RtsAIQuqMDaAxMEbIwd
zkip8k8FtjM2ETfXCsLb4YQ8LkVfEQ876EzBuLgAuNBmEcfcA+cXJhXL7Xx6xs1lnb4xoF0hEzeA
Fqat381wuacHSOw5iGPv/VTD29hgX24MQeSxnqxRT7WPO6yezG6s65lCHXQ02qEKHXI/XrkuxXvg
4y8EmjmUypuksEcBhDUtSsY4Da094Go2I7VAiCTTDVmw6rkYiFpT+tYMExzY3pLOAd5aCLax82s8
cV9Fbei/+b5BtxOKUsblEepwPkTcjiJHAHiHSVLqJNz/LVzfzBZ0QM4mxjef+M6HXajz+D75s401
psZ2mH+JXualFz4VWTgAU2yMXDb7ezTQtsIHRAWWy81lI5EX0GF7CTHeXT8FIg9tTFvb+k1hHx/+
9lUUU3ZI83+5nj2vhX209/Q1UQMyaD14IxvozPFTm7AqUk67Pq0eDJme3Symxu430T3V/7HBTIYN
5bXGq3nHZS/Ofk0t4sV4Fi15nm8s/5iHRAZcE7b/6wZWp38SL9AMKmK392zF7txgvZ2AvA8Qm8Of
T+zSDcLwVVQplOCa/9+p3VUEcoEimAdOfoW/bEuRZC8ob0k0Oz2ay4wzTQm5WHwCmr1TAldfGk/b
xHyU7P8ksOk3DJhu666NGAQAOwlWW51xJVcOAq9C290VfrLxU9Xk2JpDkCDFRFHqDIDToXS1dXbf
C5BMaA1pIRt73xNOH/07u3c6oxhjkypM0CT9i6QQQkfxUBg5z8ljTEitSN+nGt2mwrX1BHcL58xH
eNqNEJU6TrElQujYIBvUZSN7Xj1GAPMPl8GY63teCjVASRdCGc2S2Nq70uDirL4AKw5JiGc3rq+O
oM1y9yOl8bP2KTsNs8Sj9CB4f9p2+q3UadLa4RkNLd9DmhNWu/E2DsK29bCk/xhwzMvUPuV4qozc
ahWQvQPt2uThxywVdjo6hG4HEVu+oJ6QcRE29yejCVIfvvSDi9AsRPW84cIVm0PAYJbF1dt7L4Ed
ZKkUdEZ2M0eHw8uD2vSsPWiT8QXqMi3QOkUOR03vYvFVbmIpcCKO/LSAIIQCIOqormgesVMaL8Le
jlqB5TS1EwYqda66/IKVwMHKz4lhYhhAoabbM5Vp4zckN93voL2CNaiWRczJiuCvPcbW8XYhHSKB
c8FvKnLneuxUTr68slkYQ6EIK5p4UQzgIongNxv5BA2DTXSg/UJm4mKcGABnJfUvx6mkF8Rv2LYr
4YJhbXqW+QkNDmeW3ziYqzMNmUDmZXZlvFJzOOpaqxDwZT3/MnD9QTG7CHWm09X9z8SbgFlL25u8
8/z8sAB3o2EShRlWk8DYGODz6osYtoLXwKG7lBdGTb7KCl6Z0b66a10gdm3xjse43U3McGOoGAb6
NAdwKYOpTAltqQcUBa9C+SupTO0Zk1iewU8jAX+Ru48VxZuZLEnwqnPUjHQUkiKKZ+xJo2eExKls
nC+KlaC8URvoekKPTNmafkvvPJLpKw4uXd6gPtyUp4MqjyScXJXJFUo3ec72ZGAWyHgSgJ1rZmnM
D0Xilu5JY5cLIk0nSGhOmc0x6NUUaSu9luB/CycURXl1wDACoXDvgffE7jr04nZSCDQXhNmkyirS
loOx4s1p+O1LSKlu1/lcAaMoWGlR7vNSx3xkmwX3M390zRVdttIxFS9nM6z9s1E0wYUpiVuASNc5
RLc/bG4ne3xa4FJcv4/K8WzsFZmctmfFpYpz1FX2hYki/ERQa781HSOkFqWBdIDpQYhT4OiRVeCv
VRM0DgGHJc3lCFvP++ACNSvH9LaA2A6UIphJZ+eVBSybQycVFlHZfH517KArjc6ZaCNIaMPCNSSc
s4ulwDfqetVbOU6NnRmRsq/fx/mhs758WXMQHQ6/cP1L/mgjhg4i6So8m6OMt4YPyE8Zkv34m+lL
/KGP0frPVwayY/wB183eDPml3eRw++Z39cfFXnfRdMl+56zg6sYdzW5MiK3bQelnNGyrudeS9R7B
fZ9P5rfoe0KxjBNka5ft2tzfdkUYDUF3l1JZafPel8V1Q71vj/2bOesLJtMEKxl2nOEUGeqWIN8l
z/yAQGLgfExFKel9vWzFE5PWU+Q8bJk0tbcKV1VQMm0xXQ+kEIuCjR0O9qpa31/Oc9KAQzZ2DgeV
7IGSfcF3sTwL5tPErgqtXxsfc5YDyoanffHC/Q4Hpj1I2QSVGRKxkc0VofcT22fJSsNuPoYEMbif
7GaDAiPokfNy7CcIb+agNfYHeDxlxmaqz3dMCa1eO/8pwJhoi3HUhtPi1PQVXke+m6DuBtJtu5Mb
zJ2q8JCGPoqtjblWQd2QrG3KobnZvI3DQS0vvl1cmH/6D/k55h/E01iD7qkUQQESHcnfnQs1S0EQ
93tgKMTbGzH+ORsjcWE4xiwxFclwaHlii7cscTBsbU+3OQWngZjh3y67y6M8p9nxKSbiRlS3WC0R
shENxY1K77XqcQxqNSF1iHQ0qQdYY2npmMuDMGfbqgwOOBJioznp4td12ZUhTAMwsGSoWM5D1oai
XYXlDmMv5Qf7h7VJm46ggb2z19MWL9mCn83bxhRfL7X6Kk/T7aKcrH4tuUlf4sDfEos/euAibX2T
e8CQz8iVQQgtrEEZ+uXAfNzHzzjyiNcY98mjwRoM6eAfffqnKg6of1H9cAKzb850cPSwzdZOV/HS
OISsuj74iCyIA37K2+WXsAMKCIEXZbg6CFJ2c9mdF+sM2NEj+aDVG2of99ymFSNPe+cVLiS89qsN
5QwZEnh97i+nr/gPGSqx8igcVsqLufE6eKYUAFM9cQCJBD3yXWwCAL1N0MxFffI1r5POebfj+vSH
amhFxVQC1xtVCalXXtHgRhlSESf/XjHUQ3QErlAAaM4qCT6TlHLJXnNyzREEOwTZ5HlcagUnQFCH
qj9vuzXeKMzjNqaE7maJRfV5fp2o0EiEY5NOOIKk6/vW7uotpsre3VUAYUlfBhsvx43/cpLPa570
8rcP75HIlDKVBVLCmNOk2mKppqNs80VzqGbPwAr+jR21loTeWRlXVEK88a/nI50qIiSPpbiJC3Qm
4IA0GR5nD+IBV25NqQR7XRnr854eQWYHpSzGn6wa582tB35TvbkSgqKPcLdMyOg7L83fmIS2rqB7
8hOWfRVk1GdOGTPloNfMB0MamHtSyXqgbrcVOuERS+I8g75TuHgYKL5VfwUgIUwci66MnTtMIOAZ
1NRVn3GR8I9c8teVrEI1huNzD4o3UKh7UpJQx409vfN33JKbYaWzG43LkPWvCF9cG/0H5IExugf8
eE+1IVbZkLXfaIFW/wAalNQStJzrb0aXKE77xSkbhJT8DTqHPufMPu8F23NGw9skj0raH5hswDBL
XP7YyCr2gH64QJmnot/r4GrBFp4hl4ZWQoWherheJY8wPSYYtXl/iuYN11ggBSHb0o9HgZpFX8/l
/XTX2ex2X2uEGkr2Sjn5PpcVisUSLdBp1sdWUg/d0Q85xdmO5Mx4gi6J5vKBvqNtUy+MKuv01AUv
+HQENDCy8TZ/oshCbqJfa2TyBbTcL0/PepquAqx1hNAE2vsaPU2zgQA2MGq548+FzTouUu34keJU
96tLFUtWbDN7jMKiJUeGfIKNpJsVuc+c9R95l78teY76W7U4CnezVywtulyOe4FuM3lNlQe6qRTe
WP7+jE+gbF/kdMTjKWroFZ3BV3E2R/9OR5aBIyqwRnIkB/ojKOZuSN/HIXvlZroFek2QinZDQfmY
8ttLntVEdaZHWprbDKcpckUfYgGLUgMgW5k9Y3tIeMGuIMWbB5/+OYnbK+T/qvgRXYpp7jshA6dH
LCr8+Yv8kahgYUiOmY1SEl7GC58JCH0V+z2eLb4vo+EtLynnd/75mDeTfhSRmPFi1zN6Yb08VGuJ
29k/Lue0S/iSfMyKkhxayjW/N5UX48NdFhJNRg2R/CoaLpIlR4HvUjwlB4Z+EMjVhwnWJiXR/17O
2VHHlk/TaBcDSjjKRl7TJf78CXLtnWmK5RJC3VKqFPWf8pUfLRK84TkkkaK79o0F0UuT/JT/xqSi
9FsVe29NTM9t7KhzWfZOjTB3+++PDvI/61zYuRz1RgeXDSepA3qLIcBfNycb3rIW+XBtzvqiEjc8
YXG7n3ZrF0EGB/s0aCZPFgMJl/L2c41ZMrP1e24UarL1XuQjQROnyYNEAocl1DLjzRDQYUgPUyI7
F016x2jddALuz9ST5PlgdcSLO/Nl03k3G3kzZHRTNhdF1UznuFxNuwYjeKeCcUfRwx2TcYfsXdwH
mhDAbsS8Qoxfwu2ap9dHAY+VxulmTKVtoBI8yJDsMn7xwSaxiJNuiEN7Gs3WFm2YpnFzSGH22KQ/
8QrxPCtYREmXW7ui0TwOrrXbuf3eJlWFsWRPILgxqaKeuZTX03DwdYnWlCIXyhXFY01DXY/VMQz5
L3ERJbyjcioQLB5FHRmhXI/CAdtZsuRmKOtbhcxqzxowY2Z/Q0OSpFS/y8VJCLY3LJAWUnbsgbXC
EcIh/fXVgA5Xemh4uTCg2MmH94TEfDjcoTmyJWalAWkwhMowPYmmudccmEHMUQT9eO22nrtqa06y
prImo2Sg4I/wKfWwNWvHfd95Ej1MSt4NaWosopOscbHEGpIsizLzqnfyfHp4rbwUL2Dh1Hg9XCUI
WeZ3tS/aNsowgT+PX1nlGD9fJI/j/0y1njZZs3dNFCtPKBvIlOmeZ8Y/rI9I1Eht8FDveglo09jT
4n7fTrob2OHIZspEK1ApQPPby/3KjPuLAu7eBSWT8ustgZg8g5zFaYwowU5eYw5LTtOLouW+xWg2
53vexolZ+NdTT9KBV7pAggLunH2pvB6F4/FliM3BXoTQ9QjTiQMwrnQHA0TAOzWxHLsNBhayuKCH
6Y+bbFHFmk7mqqwuVcMZdPqBc9k9tl3yWMqWVDtViu7w0YgnweTRZlTg1cXjaB6Y+EwkTs9RBmWU
mcBESIagKfOriSIMBG++fgxFDmw0Da3IQT8AsdFi3xIeg6VH05KV/L115MPx+Pg5eNdPXd9ifMMf
2MwMhLE4B0BLDBnn/bjNalmHVpMjY1RFaB5pVFX2oeUA4hWPD3vOtqdwrdXHw4eymJh7l8xkUBNA
HkmjkmKXbyIcANG1XWdeIHbhH+xv51/Ppaat3D8Da6yRvYQo+WyDrThnwQUO3QhRZdyL8SeWEpid
pFpQx1YO+ano7Yr6vfzcq5GlKEKj5yJKWvA2pnU3i1N9cFiVn8efkFo/sBDzRUSh9e0XvPsGaQ1T
Ckh1FkTkDL9OG8xyLSuYc6u/HslKxjA+jcUX06RB3a8GgQ6SP36PH2GIQBnUnUg50oosF9x4C25J
Udnjga9/Gjee2le22Nn4+zGPMbuHUQmgI2Xpg2q1yvD000/kqPL4V/eKSzo20BzgOamA68vCi2H9
TPH6S0uDzYTfiplgF2xVYdoeI2nmwhFKYcyAi/BDYD5FB4Zx8Hjl8Yus3cSVDeit0LfygzVlOMmF
GXbaA49VHecaiuXypxRIaONWjaL25UXkHJMCdWExn/7UHMoMp2E1GPMkLPPAI08pXsAF+jJvPVUG
4+kHxVjrHtTKpZPCOzaYD+F5t1zztN5WMJlmSajWN6bBXYmydFtS9ytQ/0IXTfansPVK1c5/bCLd
gru6f5zNMnyoo0v2Zs69Q88nU2fveLtAAEGJxIk1VaoPAYYTrn0QUzIwrMh5dHe++euxtrufzSPF
4wqU6FGFjaBlMlZwpqXEjKMwvnlMa4cPOJkg7BxN71BzSRbVph1IuYPo57qWHrrPQUVleuBHmjyX
ODPZhIhFXvtl4XfVNn8YkkfcIMvABcKwP28cMQsbINYLE7mzQdwVgZT0mzHDvSiyNA92zoWH66CA
ZaF/FPYKsqTJ3HaQCWh0Y9YYB6KGslwcgtllcvG6NMSsWBDP5DRrVJSeKmpCnf/m9NV3e08gk5s5
c0dx5i93FqmsPAd5dRcWx+J9YwidDmDfaqydSBW71Ab7lsiTZgmQ3a3ZPzrlstWr5tOu+HCSd22p
Fx86PJpdpluiWZ8TMLgM82K3TLxPGWmB2sNnt+V6Z5CBGIZdTSOxELsShoPS0SsCDJQ9mfjdESus
0t4CXxKNcXuqQXpJR7Giv16DemsWbZqAYhh13jbOi/nGqNcAqCY+DUl5QlOMdVUa4E4zIGkmPntB
5+dhxoP/tbfzNPq8vCeWxTrGfK+w6TinIL2C3Cpwc1rWC93LQdgj5zSJF/A5/dwPShiOV5JvrtNF
gHoA1j7eVvm/yT5Gwk8tFJn+eO89++P0amcd3HmvxUHgcDIMfY3yTjHqHa4Udd+bxOXvEt5dngaA
nV/4Gsrtl+M15yS1sz7dnIcrAtdBJRW8EzN9NT04eNncy6P1i0+WS7BhbHDY4INqfnbdnzI8Nq0D
hPhbAZ3/FvnnEHKpucy19Pbt3BuGZvf0a8BLd+ZKZLN9RsWz4IfN/a9qecL8MVdqi1/INThXiw7K
T/Ixg2limZ8jl8y66zrJXFz0SE1kHiOO9l6gAmQM5aO4ifu2EfP9Nv6r0hJKPK8UPAIO/t2T83B1
pZQTOUxzBjgwQC9a/ZQtxvL3VsN6WtVJVf3fYxX6NmViUNv+a5E01Cl/WJYuKVIwgzfxlNc7lT3t
/A9QUBu1SHynPVgkq6eNEt0ub+BubqD7wvwG1YKRK3m+0VIgVJCvZiEUpQa/y/vh0ZXd8C2nO9vp
g+5G7K4fUgWM3ohRQSSGvqUeHTV6TC3rDxbYLLfEzWgdmubNlY76ssXmMUWvKXtHwgfqpw6qZ1Dg
sjJgm/+FWPk0qJbfkm/SScQsnIT8Uwe+fMwn43HO6AKxOjQY+pPvdt75pLThIHYR+kVe0Fz9LL+J
EPVyBMFGWhjANZncHk5oHfh0qg7b9ea2VhyUrDy3sE7QBIhKIWU6of7bMOxuzQpBj49nd3wfqvTc
6wY89OYDrb17/tKvdEuD29sLhWIzNWy0OjsfpWKuBtKpVbMPff19XazC2uUrGP31C/5jh2HlgWmy
8mWRLD2IARc3r+f8l3TzsD21YxJeMrauCrB3VAP0nduLp18fRFYvPNB/5ypvkXuc+WSxIGd6F/HX
O9hUvRUAD/QaMfx+Bkn567j8NiN3aaSxB8h/76uI3vzWrP/UP+vHvH65Vm8hK23sE0cEC7OZbQe2
cMbLr0K+3RMNuWEzizx3pKIeci8qk4L6/kDaH23hf/9TA1KxsRPw5cqvjIu+ZXfkcEuTxk3tctA3
ZxDbP+K+90klb5Yo8ZZ73Vi2JqchbcsJ0uu/vfbz2Qd3izmYpUWfZah8Djk3+fHodDTDgedCMs66
K9YYoBpGC1v+HuWS3KVgZXjcnihpCWpNC/yhxVKBx7yVUnaaMBXjM3j9t2HAn4iBH4Tzv1tVHNkL
Px2mQ7Fk526+C3uSzLxC2yh8MUZ9HhdrQt3tV3BpPOs1rg+6LjLJIy0hob0WRngS6AAlDMKjRyXQ
2Uwy4SYYpuLdukiVtv8JcMVn2M1iOKLEr0cc+nUpjONlI+xL8nD23mC3Uo3s9yNxIOwiVxepM3y4
8au8hk8l7yKni5YH10RBTpb7zaRMzfIEMyD4mBv78qhuPFSw5l8Vkgq7rDTgn+3IGypQPaJ3O1kZ
BrwOjTsjV3hkEXSbUUEcNrRKJwA293jG+ijmRJTkSTXJ7Y5Go4y0Lp+WvpYETflmiEj1hJLGKD28
G437qa1OvkBo2tMiGZl3P6LfD7OSIWOm8R8ZMRx5zSXoKy7Y4aqnDLvq2gGu+P4UMx/XDSkqX4zi
p+ETDd7eyP4j+yge1nANGaCyUW9SxXtmfdU1zaqKMwKdaHA8UHFev2cd8gpc8DU/Vy5avLLk3oCK
NGPdM7QZOfUVQXrVA2R4zWGCJymZGo4KbDAuTigj6hKDRtYhjNgOsD18Iv214byXzXXYHfBpe1CY
/BX//I7slpQXlMz6GB6pRuLMQ//DZDcDtsSwUmpvxuVAWhbciudTNyW0tB6QfrlQd2DOkBpOzgYu
RNRMRCO1uf6f0oOqDSLLUXneJiqp5E5928SlK3brYDWdYNGPQnOl6Wx8i72PMQLwPZodkalIlMH9
if5odbjLi1WZqe0CjrhKLj1oBUyn5ua9ozq5B3KfWd1OS4gD9/llorL60g64QzW51Y1ElWkt4qnj
HG/bUITzrX9AuH8ERkGXB7i2C4ugCPLa5g9OyjsLxSr3Th7drOmYxqUpFt3IEQ7mOB+vMaM6g7Z2
PYQ5RAxQTN6Z6NUVZBuaYQsmWjb1GrGMv3zXN/sOdnyJOeLaaJXQpt/91kU3WSUfqfL8puaw2J2u
pUA5Y+Zk1paLLOsBDbK4rL9sMwa6HfMXrNE3w59H1GEsAOqz28GdnT2rQOY/r2n5D46wPNgWuQcK
1IjX2OuLqN9Ar2ww6kTzg0EWQ+TimGXSj1Uk8aUviyn5+evHmp6wFhgf4gY+WGsdZmrzIQSxwr0G
9GkEI6Rh9z3ANoJc29Q3ykhv6tgbUxPlk7MWLW/a2h8utcLTXBccGmrAAkbSKFAwHAHpRo/zj+gE
ECFlbbBQk7s9XOXEfaPYDTj70mUxB47ZvvhUZ+X6qRIjGXVd71FFWjwTb2n/x8r9LWUl2uhNWcHW
9t5Wjhq+qbGIBXm0roNi3MPYzS9KagdQ+f8Sg7F7xyEfnTm8UF5FVhueltI+fmgyD5NrbWWUI039
mXa8fLQPajI1hjq3mbDIa83XmYjzvjD2j/0ZOyrJxGD+kevvSreOUzayf20yreuqYYubx7mGMWqI
OCiL9JYh5jFk/PVbwiGPCPeX4Ucen0MtMxWRYELXk84YxwGC/O9Sei7voZsWD06VePJmWZFTMcpL
JuR6CXMosjooRleOuQZ7uOe6eFNuMH54Kd9SWV8kat50B2HLZ2NHVrCvg1K5yqI2rsAV8/xBDVe0
zrdzXuFqWa1O7ur0G5XbVH0980rljJlR4w4FriFOkNWbMUXJxInnhQMHRoWfHKt1CDUnrN6T4r3O
NJzxo/FOHvmjQpl1rBzguB1y8fQA9lRa4j8Wd0TGCGWnsskgcglcAZmFX5ovaGwr+EuTbmBZ+/Ru
4MbCZ1gDktCJXlZ+LUd2d6cFtmKUFri9jN2I6gWcPwUQErQbCDm9Mv1hGPu8MTx2eyd9JUc9SH9/
/1qUYrl53rD/mPNVCtgGxLHbjibF8Qp8xHzJpBDQW2+MHrdq0csMlDhapZLavE2Vfx2j5raDzCiK
0DV6l+c6deByHrVZglkbzZTDaxbLonQQbuZ/znjHNC8wD1PAiH+nWaS4tOi9HHva10SJ5DOGsexo
YaZ9WTv1JSMFEPbc2oQQu4FRVbQy+RwswYStoBW+eilao2vJtppYzpYtE2QPD6OhjXPBZwuLWzSz
XvWdfCvYWdzUOGyqL0xp480+HHeGYrjI/3A47P6Ec2L3totavKXVhXfCbFL4FBiwjbFg6LfW6O92
nLcXg3gubv3esuMGWaQNVjD+VDOcRKuVUlRd0jMtybRlSNkrGgblORKBBev00axnwHz8WTIBL0sD
osK3unedOdUtiev3xqYkXlp397zRx1/8Mz11FmujrobQciHTSHpRJsfY+ROTaVMmVxwA+QGhRMDR
OuZG/K8jT26r12sSxUwEIH99PdC+34/iskBRxZBkDWx4o+GSzLoZDIjtbfR61i871PL+mWekyEp2
ySXaE1tmYk8duJAelYRPvpRLpURm0bt3VXc+UvaLYfgCEZx+Q5Pt+0tkMA2uouXb9EW78n2VxEuK
4+qvpR/6cDeuRER+w8vAqdIb1VN87ixUr4wjtRb10tBNI3cmZqjW2YtKz0EcKRhdWOnfuHFrBe6N
7JZYAu5fk6GqyXGcbXmsyBs1VMucGWcK/ZrRoJ0mTocmKgDJeFKp90CoVYMbXCrUG6PguEhVm0WY
/x2W/YfHC8JAUePz0202JKEtsLFWSSjk1eri8dYtSUTqxIhHhlbBd02L60vaQvl43W3JfYH8NgE9
9pG7u69Wtckh5arLFSTfqar3DWBap1FmVnlLi9mhkfnZOI870dE/Zqu3EgxPZmS+TBOVzjACiEHz
jjpstxZvkQ9KVX8+YuLcouk96X+qK5c9ewjCEUzWELEWz/YdsVFMHvntcbX1VYooVsVeBSTZSgVq
mSnACol9DH49unpYAsfqQRrYFQHdK+3VpWw1VdMlFoPP4yJGlhv4yi90Y/UwF/rhQQbg48GWnlDz
0bpJVVR20OGRMJK+/kMIE27Q0kOF/bDXpkfHCGczs3ZxSv72WxB9b4MtAUrZguNzNUtXssEdGU2r
ycaQrniCJeHFXBwOHb6lHZf5SviCeXuA+a7IZ5mWfWpm4ymO7P4N0C/j4Exl/rxXxLwh6Eo4RM+O
hFZwZ9FLn7BxNtxSnjGoqPubzIjNENYPlQ/aNswOgeS/93lwY+9PvPevL+jnEN8UQcFGYjHKFvjY
lBvWOsaQ0z33eWVyfJK97v/aIXD7MymtELiIwX8w+tnhEd3dKvqU/Tx9AEquiIThJZ0mEFbHl8W/
xnoQNoXxtjgsi7cR/qAHPLudE2v1c3UoTVO00/iQ/SCxKbFQCay3Ook97ZblbXII8ksY60fNnZai
ox8jt+NX4BR9FGprxLaactcZYNq98uHdocbi0fAPJS0UoJ33rQQfXxl/ekIKmi0OWIvhwhcEv2qY
qzijE2QTnbS+cOxfcFnMWD3B9pSNcpxuriUAHdlc8v6CwMVgL3PXe4/AkhLcQspBpsxqqDzPUVKg
DCxI/LTWs/BvK23n297K+9prEhtmsLQpYM2DKRFYiTFNk3y0TtffYhJ+lzXex7tt8ytY19HqwA11
SuzFioKdqYJpqKTOdCplnchY7daCoZhYbRNd7muQjzNlIh2EaoZjP9X/lCnUL/Ma1ghSGjaTDqA8
bRNFS5AGVhqC82zsfE4o/cssaarnCqwJCCpWZCODncOG+GMyFlUtptHjrhX4XagTMSJo+GDtxfe5
TF5ff8bWghVbD6YRWI5obRsrAoHPvxQq7Aqh3omt/v2EwdiErAuMYYsUj3WbLWEQKcW7MRSLpoIf
ZcUcd4xkbEV/eju1nzoqcuuWF6fOuS5uF5gJpBSTYT7rxu+D5nW7FM583uC0V3UcElPIe39GiJxP
UYwxUbzS9+z+IaHE1n7D2e4V01Va55hJMbf97R6nD96nGTtuqdjc1gXAN6m6lANjPOAHSD3mYHh7
Xl2Ln6ibUwOgogsaBXE+wLcN7WtFmjzLEzI6ppH0z+uI4RzghQwSRzJIB7bwuOE6LBaherqASStL
oMTmJGqIfzmg+PoW5+IMGQrW3JieYb5+cDt1TjptXIKu9vmENgHttYF+WXj5eHzq1oNMqzw0pJWh
w0zLMA5ef7Ztep3wVgRs9RwSWaRh5sB/LXnNocTTJPUF7Djh+i2/2cTs6hnS1K0GCIvJ3YTtNOcU
w3HOeBzRn2nQJpQKzEOZHTEroFRgbF1+3xMdWIfaoN3foiJzAsYa4Hk+f94TX04Uo6iSUD96tU61
0KCPdQ9JI/uvCmQ+WLV6T6icNf8V4mnftwQ+GA/akFh1DtutwIXd58go76K5Kl/H+gI+T8MxvE5k
kUl0t0oxajYSuE+XfPq8mQUG5Raau9PVUIGzAIHvUrchGKd/2a6tEaLtLm5aRyg+lloFbsbmLSsr
WijQdPjY7DxtHXLC2ottBvipYk7rlyss3zo8LawHEFLM3/okva4PCg5UVUnzXbJnlYjoHV/zIEpr
Z+cVGT7xbrR3Dk6ldNo1zByUobDeaBUaH/zD/G8FGZTeEbAMIfs73kOI9NLRFuN3798KVEEzvHi/
Xu238a10YWAd4dfM7xIW/OUHHKy508ZGWXq0+c0UdaqSsq89bBaL+g+x6jiJM1WJ26tNTf3G7y8F
5CmHC7fGLpOsCrWNu/2fqammWmQGMenUIeH6n2gKhpyiVjJ79xciHeS32lT48Nd9lcRDTdOGO62+
9557++jZRmhd/vqv3ZPrgwH2vwk07cwd3xoPbt3vCmX5yECllUUKLQrR7OUZx/fUO7D89RBYyT4/
nazizdd+6xOaon7BFFABBZhlC/X0gNQMbibIeJE8PP4YZX1qtVrTmKTVU7kWddAASzVvb3NTqR4/
wWMtUcvsSz25YyTtE+EhNzngWdWVPzkDf8cB5E1JW/rgzTxu/T+dG1L6Y46Czafk0O2kjj8GYSbn
7WixBxsRwG/0MiElEYvDzuAEj+pAIkiTvBtKKjE4X6h5eV/FKS1fz9G4J/Y2Spw8GsSCk0nErHBn
54Kdt8ripVqVjBS4CFLyVWoXJyKdR1VS7Fj2OiVAG06B0s8fbbAOFyL3X7KmNf+sp0dKmlcq/gwP
XXiM5PKHvjdVESUGAv5NN2BxVQYVosKAyDCzpBHR5911ohVIYXj68FVFcSE1flBF1fS5z/tiekUT
mkO1eB1fqU722QrJaBlGtEpKZpmgbSA/i8dQVmovV0YKO/3wHODIi9BttcNmndxXGeokxIB9MS6v
daFwB/56Qp26BY1kDddDzpy0TIK7dql0ueO8u8uKDjgH36yVOYvqqZ/jSCw1sl1cfLSZOp64qyLe
AS0HYhEMckjzZNMVlL5F7RkvyJiWhdJPzrpKkmwSKDXCPvjqeqiZp9eWFKIKAbHZWImpTOggPzi9
llJbOgooBLGvjYhMhp8j5uaK87kDSj1B9wPyFdr0QiQChn5FKpYWIindqCcajbxErywZiQvKY1hn
FCfFlc7Ta+8kNlTBPp68gWrYZYoe1HNOoGzOzYfywWA89ImgXCANU/3lkOaTuOQxJn2+wVVzfMd4
RR0U2lXgbuE9FEJmEZwcLGaaAx8/AhZcSSla7Q8LmF9MQlGV5k4/ubqR8Q/bYrYXYCVfKycCzrl+
q+H58F7ByyrqpqvFrvn8/5CQfZZtqzdI8mzjO9PinRnE9gcq32TDTkG5wMFGaiw6H5mhlcs+bo+e
yo4mKuNh8iLlI77e04fdu/QV9hHZHbsbtkEjCn8itCeoopHOGTWkRBeITZypMx85W5u8uXPVNFRP
ecwMHWc78tNaBnFw2GSL7mG/pQ1KTgs+Epsono+3M63iA5zFTG9CQT+MZbNkHRZbAvufMeAwu5/O
9hx/bdWBeH5sjENivEPxyjx1KPDxhEyu+zLnxZ+5pzUoJPTj0iYoh2GAJfIgkeiOT99Tlv1EdqWD
pWZgOkh5OCJh2ZUJWEwHJhTn1Jtoa8swe+wREaYDW0BNvaWbbJzdIlZN5FU+K7U/xbmqel4cGGJq
+JwPCtVhCeqpcdq7c8F0evfeyioPgdJdDiVqtKpk/7aze5lGSJhytUvABBCNdTL4vMCaySTqvayd
oJCSV+aItum0oo9HMQOZrmE6oFArC2TJhoeM2YpYQiMtGNDgmSkuoNbhUxu7K8TlSEYIwdBs5mSa
3g1vIUs1rRvNTP0tL52SrqO3iT6d1inPTZi3UoIjQuzkzfb5U+hChIbfvWTVgu571IoZGHf07Y60
mr9hTMatiVOu85wM5Pe/LLHzzuFmKXSvskK7wHefQ5MaJHWgoyGIJaI+mokdLiPdLOXlamCI7ilf
EzF4hT9Ah3Wjw3L6YdbeeeNuQAdZOr26Rt0TWLSpwEm/2CCAuIhwwAgB+RHxRNPYPTOQbOmZjL8k
0Mgmi3q2vksosXcfGhnsk+qW7lO1cDRllt+Kjh5CJ2uHg0eAT0DiapNcc1TZXaJIw7V10WJjrVu1
rAyB2ExjjauoL9wBsinKxnlBXGHIl0WwSv+RkcrFPQeLLFL70r4mBP9kn/9HG8UUetGL5Ey87AAT
R4zy2ve6yCjQZOwspyJtmwEtjjkzU7l1KEfVB1EynUYVENZWywfj2KsWSPQZNOhrsHTH1cqonp3L
8f6m+aQ8cJab2GuvEPa94JpK2Rmz6Ze8xhp/MPGNOcHouuEKEcQ4tI76n+7juGv4iNF2v4ZYHefC
ihFIPYwQlyrZBCVMYZJItAyXNpoWOzerTRn6LQ8AYjaswl5YZ2/xUSZrFwhmim/VenTMVD31woAP
SjGCVqusxDjUvGUxckg9xrapf9d/428vdANSwx9pR9nR2pP0JFoidegSnPUYLYVgqWDTqwuxjgF6
AmazgOtFaSUohweQbPMP4P2gjIbUNInI4VLc6KF0fnNJP8VFoxEi0YwOfb+WgSBoGB3L/wXhoKVE
ePCmrKq7spVOszdMuCrtcUWZsNf+32Ae5jaU57UK1vwJS7v/nAV/OyUE+OmcPCYCsbS8RTBp6bEm
oEW6lEBWdo30xCuLfZ5HnrKhJUCg9nOSXS+v1l901bRUAOmjdK76qemXjgglns4HhjIGn43XiEbk
i+ibFgJZVvk0eq++nk+aRxAmmxRKkTkmgYwYCAsl85XpwoC6w1Z2rSu7gSebbakWPJJ2Y5jth9HV
22NTvbhlPiDMImHlfMy1w0Q0IQWMGJmndPkjkDRQuK5EX+n8XI+DX8x0JvEwSrl5l//W8DCk9h3p
O2fJJDoOMlZUu6gWhJ+8isChBor/3UNhPc37jZUgKP3PPHIka8w05fHGfg3sLV+Bt0bVYst+z98K
11tO0JIgXma/FaNDxfO0gxNmtMGTN8CvtxZ57X7bjqzrTOdzz4BDH6Q+uXbZSfvQ083ngTSfX3Um
LwdJcXu9LnLO5igbRwnbEp7nb5TUEilEjNwkPJNlEWQYNiLCqDHB20I5tAXbKuJbPbOrugz4KtZS
K7Fj6R0+wmmDqdX+mmcDHejsiIvrOir+Td3l3aUOb+zgxtKxPVlmwHkyuFKh1yA0d6c/gK4vC1Bd
QEhE9+ye4KgxtExLgw6Q9BVb+8J+T8SesHj9/aWdIkopN01w8dyTvQKzwnyfotJBntcRBYzcRZlM
uaPgMz8X8TC3ggeW1MtcFW+RB+LWesH4vCs361iIiesmmy9VoJvhXvywZR/HUE1eoEj5Ga0hzKM3
Zjgio/NWhkD17kymY3KTZO+WUSow25n9gc0Z2b6OzmgbNrU6rj8LKV270dWYtOaAH90CZwAvPqtD
lXeMSO6UjXo2CjKo7mM+/o7SLr04hq7a0Y3kFmoVl3f78kmJyJu3jFdfpWG996Uk6uMUh5bcLmTi
rbdvLm2sxqn+v1zLx+IfGAr/dLT0Smn/+G58deeMGt5lbGJes2QpUUo+okG1NvO1GawnCEtUVWqI
ufc1rxfW+M3CVvSao+sxJR7TlaGKBrm9+8VxVM9jBeJjZCIZkXYQoqlsc0ZeaNL8tJCqtA2yDrln
HZ6GK7Cb9BBZrO0j3NHlSe9D1HLeOHp23RQNFqMcXkr14c87l1xup8SvAT5CdWZn8Xd93HfBvALM
NAaG6J7ELMMB2C6qQK0yfM2okyCK+of0n9FoC26zoqVMU8Ct3uILMIH4JVa8pxlegnvJONE9inK2
EIMlyVXMDL08A6vQpr3zEtmIILj+M+o1y4IowDnooE5WivXgHjJ3OYfZWMF3KmD+0Xkzl5AqubS/
c+w8XmY6+FoWdU8RqRS8SnFbYPdMJRE3p610DcykevA/hJQhxb0cRRsdzcpw0YMar8Xt8+f+l8Hf
RZ3GKnoYrMuWNSP2RfFBJyFxfKlGng4pnZRigwv7zZ79PBrZEubXsK7eeVEk/jSBdk+P7F2P2EWa
X4wKo7Hvm9vi3bwPVz7eQhvXBlO/bKRTy0b0cjuJiq43hBqNxbmalx+XBkh7yBI3ITvoSL38hEnV
NK3suL9I62bqi07ncFfh7EX96wkPJH4CuU5VAxb6Tp37OXCjHiZx+ZwWC4rkecGW4HnIEHo3Q39Z
hxe7F8xYjovHHHNCe6br1K/f8sBIA8l2KNhELT6DO9JKMKbKmiZRY9MHxQSsnazajJ+TrgJxzULI
QfUKHr27Q0iFYs+Dd7yIG79kggtdAdYdzYdE/zx4o+LKNYACD6fd4nZJJpNKNY6ExLer7YVzXeS8
f06/dB/qF/UNMyGdW3e/ndetsmTq7hnaKuCjgDBoV9yPVINoXC6ZgfEilkc9ke0qey0b9xmAdk/t
eSk/HkSBcmWM1ahvZX9dh4pbRAvYzKc1/7bwdYhJlXr2pK36s3D31xsHeJszdezlwkjeewBDSRgV
ZWoV/SLGdhnQRKboyv5QpW6lv/wukQxfEZH/LwwwkD9jAub0JRgdhtCWlQxe/RANrib0nVsG63Ws
RqQZYf5+BchaBXAaO7rwTKYJB9iRbWwMy1ly/36ihlHEG0LX+zWL5DqO30MFY+4yvCgVWJ8p4av7
+5TBVqiCbq7yiRCUlCWprFBFp9AOT50DdaybyrKXMV4vvHVU+zr6Y1m1E/fTCGv/EsIf3SCump1/
LiQaS8oztgYSz8xlOP70RYuXm3RmbeRpXhBngDa+O0fcYp+OvXn1PkSaKeIjJFUWGCZnqDFIJJWF
699Wcdk3y2jiWdpPq+BTmVWoXVJ0qFNL0KPyAt5V/fdmk52ujvSQWODtafULZg5FV0iJhfTODHQG
iQ/j0GFjQ5FMMf9h/EdephguVtF1hbXh9hdc3+C27AQGGa7/BRPpvDijIjdlnT56jGW8Pb9fZCBW
qAeYlU1sDve3kWJPf7PfeqhqB2sd4E+eWutKqZYv3X/EQEmEsoob2ZYE8TjejZiFKhmftlTA2XG4
ynwvKncmhdbRA6ob1GAU1GXwbmR5ebTVSdBtVok5wZO+kR2xJAQ96otuk10w7pEODmCfQlfptVDO
3dObRD2TeehzgSeQ94WDHCINPsLH3qKKaCqz34O/d8m5zwvdWiMQEx1xeJv3dso1OfE/uy+IO2a0
/m4/ohBTKZyszOeyEqyNsfd9b3AMhDYYg3bCCBWOret55GAYsLQ+wgJOmtcsC4gYyiItWNW1jln3
Ft+zkxxP5kvzzhJXoLKcqrar7vWmPWbUUcX57r+222NX/Z6qS9/btHmHrlS7Dxaa+2zap5B7RiO4
EPdwySANehoLugFIQSzRyUPNCV6nazqIYQigUwyWEN3jvf+TLVXFQ2BLbej0TWlmVe5S647wmsgA
2voo9xhDFfAeHlIX+h3Jiu+KyZq6SNuKG6UmnVoPtD0Hu8tvbF8k8ajwixfjelOmBZ+eETtoaAwA
agMBBnl0Xv37f/K7xuNOqxKYThlj+N5BMmvGZFPzGVSDwKOaycDqZJLp4mIpZ+/gNrKi+7jgMdNI
tfh/nT1khb64mG/4YCfnWAZWJqWbKVbdII9mE0w19zfH5ZVkasNQLqyWyDLbyR6ClQWS0qqT7PP3
0KTo3Cjq4zzU2VaVtqo99N/n3it614sKl8YJM3cblGIMoaNiSbhBuRd0YbH89Yxroeif/9n06Cse
rMWOabuhFy2wz+JltLHbPGg/JAcK36QnY84jkRgeCP6JDKKP5MIIC03QTKIxUlvr8KBZ/YAkhujX
lJIOKIqApJoIzTEGrxsU6CPFzppdzyKZhuZ4zW2pDLmBsIbDoUNaM2xexuEJ0fPXD/l5OGJLvf3O
1IBZwYonVlkBcolB3VM3cyzgnr4kvZbs89UdFwnhuMlP3B5QdNZ8zA2xw77cOxvRxMYJLxH2kcNi
uN4h8eLyiVG7qUf3S0zAf7QQi3gRPvjwZ5bhARpkEOchLGFSt8Bo53d84RtABbS/sY6RHkyMcMAw
E7iufuFXyG4x0fi0beDeVAKhh+XXU9LzyE/v2R76bbvdzZtCNm3lSVc5b1MOi1v32NPaevx5rOKE
DJpasr7Q5rNN7o0AF5wYH1ROemZHY2frbEHaZSQkrKGzWB3zdiJyTqoCx+44apWuvQq4Qbv+3SDM
GpS2too5MGvUiEv9BYS93VJA3ekhbF0w2yhaTj5fw9+vtxMu/tdHxhriLE35AxQIIzO7Hah4oLVB
oLwlfO0sTrWPX1OAOcq9UsC7Gvvny9rAcDkzZ6k2c4JLGJQTcz7yq7+h38ZlILzL+Yts/QAgMvrn
npYflMSKGz/bnudXOyWr/cIBRYMFMZnCYCiooa81MtCVGefFRnVcP24CWVaVrW237EwSM/AMA5Gy
qV683LtEIx4HM6Bmww3McmUfpSIBfiEslmptKxmj+/Dvm3506599YfSRI3Hk71JDDHTCPsr8YwxX
Kve70rWqf5BYJH8d5+fSZ6n6IHm6Ycam+xFvHXGsShO6ZuhRaXV1LUnij9oKDxI7380VmWCzmZMq
KrzIj4JRqJ+kvoZQi9igkYd3b08m0wy8VKLm+pqc6YifAxbZR+GlZUOvG7aZrFrI+GO/sti5qRR/
c3bcq49mE5lDflMLmH2ZsWzYaspdrC6KiXWv8DazthYsVttnx5zfRIcJdzOMi9TDkf8HWFOheqfS
eRmMdjpqSoHCgGsqrCs7T03vSiMioJiecOfxQxmN80w1z7nMhhyMlnNjRxWffjT0fX2GNZo+6KiA
Vpb6UUqdhoYUfkBbAx7gw507rKrd0AONFxzvmGcxzZYwElrJNNSeRAhNTqgVq9wEHB47Jb/OqAyG
4kciKbvVSGTlwOoZcSeUV2HqCtA3phYjCiguQH70+s4ZoPEy4X3/9zOxtfGMv2lDGOz0dDYGJ7BQ
l9Kn69LVKU5RR/8WWZogWwcK+ooVDBfKneiLF4WUGu7Iw8TPryt4Vmqh6y3JLDMyNN6V+sGolGcg
1M+aoCRNBHaLtJqKXkCsMFPUA6tKQqoAlnhGyw4o2/jqlh/TpuQYyY9ULIcnrMdCi1QVITGPwd23
Ho6Fa+I31p0HyDoKPdFGkvgqPNLE3Wqw4fNJbX2vIeIHZnKn1oRN92G6iJdNCBDta1U9+O2UqqKa
hyAIvoQkShPBemSHS55x4UwP1i2QYVl8sSj073aq3LnluaxYrSfwcRN6m9rf0HTy3sZvfbWLnak1
v9qPrh6a0FGjj3K2LPezU4PKKMdhizJNpXPxvi0IFrQGcv0Q+9Qcl0OBtaIFkH/ar7698ueqCeLd
rtriA7hX9h5ycVcW/yqwiuXPcQrViXLZbQhh9edMR3v+LHegnmc2RoVzpoMcnbPVLnlneg9YK8xt
uHLJQQXdLuo+CNLVoDdvltIag0ODCYtXxPjvmp646Vxy3PfArsWuhEHYN5fF/h81ZvDtC2Zl2sbj
NC47VoS8NdF2DNZ3SGYWZDc2ndp1dsHTFRxcuJ+lbQ4RLwMJZiE9j6tuBAXZwoqMGQycl6dTJm2u
mUI9UJXiMIIjjMSjaoFlKKNw+Az8V2NeJarl+V6P2fGMcWJXWZZCOk4njbRDIc/s+vIrchVImlE7
kAj85sD4i1TvEeaJHCHp6qrg7jhGWKfR87UqutsiiOFvMPlyIa3psV8dMtkHJhXYVSQV4Lqzarzv
0DMT4nS7WRbNGkiaw8+j8myXl5yhpCqRUs3duH0nJROmlWCAIQT85EYV2v+HuL65R4AohD0l8DSc
g7KuyTBa6YzWsF3T/9jYHk7uupkP70CAojAL6zUwGAF8vLivVLprZeoDeyUvtddpvMSrJhECmNM0
HafTebw+xhwtWk6NttWWmdgdiSbvtbIbK3ef3XPaSBToRuUe+774hqEA85Ibf/cFahvft/OP31H4
0q0LiS3slwBmiNblC8Lq97gn1SM+SsyYo/CjfDFFydENKnBPtGldgkSvA7RUNGDfMGwItBqbfMk6
CwCkKAa/gXFPFhXditXaJqN8mtJVHeKySC/hEdubD3ydFueqkPuiKVgtj6uHxhR/Hie2JnS3XmmM
+pscjhzUuRV7RzZpuH2iAFeq6DjtoU3o81WFrB1MuVd40QitzxL7FgeBTbMCTA9PZ1JoPSfcoxTw
1gLWgx+BtPsPSjm8cicR1Q6AjNL/1D/6gHlSuXWveajEqv6/V6Zo2xADQmKo5+IqCSVP2pAfuEVW
pt0imDKySfHw6zGUXRq03Jj8FoVAtYHaa9BO8bqoEhcJusFdrL4zkmu+miVvJGdbipbi1liYF2Oq
VQeg0xAvYoNijS8ttX0IaoWyHfh1WSWjbeUUwrMlmDxNe2dTzSBXqCsgzYNTaCD5Xu+YWAQSZ5id
npBoL4Z3BmGkQjuKkBo76oaRoSsQ3ocgYLyeNI3/D31csoiewiRKiqGPNNbcbErsDW9MKZisTreV
Hr59s20mTjYSj63TwfPkbaAarCPt4I7P4y63zj1dj6v7HNWrVwazm6JSQy1aAPUwt2FREn0kR9Ub
oaI2cFRwxalWhGLUvwqSYiOENayF0VeIV6cHnaUnJYz5NmBxtR00VVKnekZmPChhqwgXvZhlVTia
qhE7cF/tAhc6Qpff7wZo18dKeJF/CFinBLTQ1PZMZnRTE2NeEJW8E3kIDc8FTbRYJTu0quEuVgBn
mE6XXpuUxYPxugCw4bZ8/JozpTWXGeQgqwpACJShr188PkirG1KDnYHiONIth+CpsTrpIrP7zyQ1
cC1yN7gFczRGcVpHpcmdAsjN0a/0vO9aiy5Px6ocf4SCL8e1Dj8IK2oWrSG1BK1PtbCyntAPjb5T
cd3HCRut1LLYpv4ObztcJG9bF89KKoJyUcTt7bzhlpr+3ttxreXGYfdz7IeGLNueIn+WOh9QDEJl
hZU44xGnZNM/+3hMGXbbr/Jj8rc5pP4txKrMoXbB8qCOvpMhxTR6HgKWW/SZQsz2Qer+j4uv/WwE
GmqbSiFS94VMo5+zFbdhYrTB4MrEPpLimJ//XRuojCjNRaBz01ayVG8EbzHLMkLdYJQR8h2qWUS9
gpe13rXIwBGGv5Afu3HWn33sREBIw+inGZQMV8L11ugsBEBNpDpv+kbZmv8cGrDYsC2/5Hs8DdBT
zXLFX/6LUp7CIzFGwZdXMAYuVErtbpr3fKIcdyyphF6p5FDhnJYg8Njv6rXzgxzSwazpG5T11U3e
sS33x4c7cJszKeDLpYjt5ezbUJ3GwKucSmpx0IR3Pfia7ggiCOHE2dvNEjU02SOOgStw50sp8QkV
Ikhzxn9m3QT+HHbZdkBMb692DlaghxG6xKJujy/72IVd4gM/9FA+oFIoBadNWUrSKYGthCyy5oer
ZOtkmnKFvKJ8nBSNpZ4cwicEy2+rkgxfXJR2yi5MJOLyE5milOsRL/US9ayQjZNsCDyJKtGRlWf+
a3KlEg6bfTeGAjkpTiP46p9UEPhQaN/azaG+ZTs1dNHMFAWGVzSW8rmcyMlU/KUhNxxhL5BSXHyo
YIyKJDG9WjzEHu0QIYu+Yl41yfc+lmu4mM9claA9pSMw6xZCYZpEwWdmhQIs2cNpmy0cFhgdERRt
iPaSrCbJo9IP+7DpnquB5rkWcSmEypUc4BUhS1cfxVi/d/RUajoCF4IOG3pNTfpRZLWWEVHH6vAN
Kb0vhiHkWdtueKyGhPthBAEgIZZlys8Ipy3Y7JhbFEI2aov/LIW3/VB3g7YC7n2ePWS6AxJYvxjC
HrdLTG5RcVmolWIto8IFFhmd8DUOMOoKxXbWSrvNq1ypEQ0icv9TxaMtoMOcl1xslMfdSvROmxhv
b8qPa4ce4gIil26fM2cKMa/Em9Rm2XjzZDLpTIRKSk8wBajWD+cD/jxJRs69Y0rTUqc8icnZAoZo
sFwzSuMqtPLXTaabG+fQA7EOANpFagKQcCRo7sWpKX5A4rs6EqBUIzXyRMLBDLIqemSr0ie0tFm7
qQVlXBR9kF6J7q2RS7DC+Ps9TvvtRqoIg/zl7B9mIol6eAzU+28JuYYBpjHSS2uG2aKXPGZflCSK
5bQJo9PpciUyBF11Fyw5TaixuaHkW19+fy6hS7gFFmb29sDZ+aD3nsbxfzOHoQbU98XY+Dc8miTf
VuXRBkmTHMjZFBnCku+tGJY4KHhXIcfq4hwWYKVM1dDIpyyX8gecQittVRJ/4CN1JUOKiKZkfnlA
XGOWPYqsD4G3VOtdqjgprOo4HxLXAxnQxexKnpAMOnFLEM19BFCT921odp4F5iklAZ3pEGv8CLIk
tVfQ1Az18gXwCBjTT02oKU7JUSh/Q2As5ZcatMrTcqsVdi3e+Y2m3c2Zsj5EvhXSnuksZvDWdOUb
96kcdmoNLEtmPgQ1Ub2vXTJPOF7kyfP5epo20LbQlFKwHqftHFdo6GnelHM9+X19LRXgzQbuxKEy
qFa2lglxgCPY+DM7Zl+AAr39Z6tnLO0y0P8IJiv/7Ly6N2M496m1J2u3LW3JU/eUzRO7nnmaLh40
gVtbgpzA4T4LzwMoyzyK6+h6owtbvMblx4JQt+sdetFiUPA9l6+gUnL+a7GIS7/pwT8h6WSe1uHJ
FHH3Tu1HjSa2wpqIl22GhIEOHoVo8aBI25j7VqqzakJ3aWTx74mHVWTsA8eU9TU8F27P4qDXR8O0
T7qv80JbRGUp2xVuO86cGSg7o7KcMa7DAEzw5v6I8vnt6VHiQKxAz27DOV9trXhRcuS7tY2cVcsx
CEX/SIIZQDz6YNZMzZrPAXhhWXlzDaBZdXDXTEkyhhagJcPNnXlBC2QJQIXPqJZD6Dmp36N4z2Pb
B4lvF7r15F9arTYTlZcQ4oTMFIwbo5JuIozfoto1Ez5qRPijzewrfiKWV+UIzuvTcGGQJa5y4qws
ls/oQb0eSpoYeaKWw0T+3ZsT1HocqEq6hZJu5WEFsCLymiK8TIgKJYc2Zle8ziGU/PQ+599hOfkO
11O2L+TjMG9CZBI287IRXjGVA1jhVUwJ2Lak6dnXhqRAXKCnxJbyUGa08meSFiECUcoMhhqNGYxz
GqHe/yk5Edku6m92Rx04xNuWXtUxiARhCgYTJVEryjPNIU0vHoLO2goS0M3Du41RftCxnFNljwTV
IoVP1iUPiBGy0t1dGZ9lYA952GDcGhCXHjPS/U8x0Lb7xxKIxj6u3hddI8WX0/YvcEiYaLWTxY5T
cbtNlClkdZ72cwLnALShj6s/mcfBNcCZgTIIZhV/32elCaR16EwBYNPMzvMaL4KywGzKmZJm6kMG
bcEGZYi/O/GhZb+3DhvOfagOi2tt3xj28lrInXzCKCoORwOjdK+k00DEsa5Tf1S7roRwKmDYaKNO
AP40fCvcaCHYgj3EPlhp23yJzuwIJajQgUx/nO3pv7XEQ1aAKTY6YPG9Z94FvcKhmqrzNPPJRYC7
V+9f+Xmppv3THfTnwsgmDBQRG7Oc9StUfdBdzk4CSLzQAA042xjwRK2BJp+EbDWdSDAbuoQ4LKRm
ZEmKOW+lT4KexH3R11lmvb4E7TyIq6FP5bcz0ib71DraHAoF0DHVifHhPViJrlQzV9Epr+nY2XjM
ucBIKW+EdDbAV3oSRCtiELS7e9c5yQ7ssu6EoJ/J34uPQwdiRPYVgJl8SP91G2jGOQ2aUP8tLMtc
mLeRlEWuIhQXX/f/RL1rYyyID/fnBs2sNYkPvFrQuKkEltZcZXCotnxQKPfIcOyiOYgXf9/10qGH
u5v2p/y8H6bbL3O9lZ1kV0ybtFhO55n/SfVjStse98erR/HiWS0vUvQGPN5GTQwdLPPYoUExVY3R
ZPm6TPEW35LbZAhd3i68oslvR4G8c4i9vFCd8CafmPDMCKqxOsE+5gqW2b+9dUOnmN/m3hfqKOvB
AULZ+rnK3gx3pr1YLRPS4M1zYZhdmzj3VekniH+9Su+9l+FStkR93DmGrIg72pam2+8mogVCcKg7
SmmgPeA6PXXJWtSlyQbq3wc6amU0mOU4PzjHEwZAhDTYhHWytk5ObAhFqjTR9AMvZghp2mF4gW86
R+5jXLHXPc1RqUH9Mklwf9PUT1v6h/aU6uUUIX6vavFVewf6AKEX/X454QgtLkqPDKCRTfJ9M7YR
O4qjwswyvmxvE1dkZTRFqo4FS3XZvP9ZhjXywmIfLN2PvcxMaXgK5gwv0IOiDmmGqIQEiO6wNpfJ
jUtUcPn5s74c8rNQTr1+X9fiBzUnEBwOyBkbwkk8dW3tKJIPwR7G2HYZz9YdWqCHxeM4k975mWN6
VFev3qefg27W9gU06BsAS7UuaPVl7/qi5+CYB1ewtEJrcHrI8nlv0Bh4EcQd5PrKH43XHF0Umfxw
SaajNR7IaMv2wfZwIPDJQ9SCJQGBZDYppvLIFJHywxunrT2dCHKU1SgZBaB03s+d77In+yZxe5le
ta211sbmNc76kfSOHsFsDUOdVjiliJb9DXLDuWoGzQeoLfiEjpU0sqdkrPzt9ly9vhf4zOV7VEfZ
6EsHPuJGf6caLtmVTnXwgO2u2mCRSj4pERuGZSfWjRF370YYbzn0xUpXnvrD6hAoxmxFU/hvnoiD
k52ySI/1WTNqunZUUjyz7PYBuquHHPf8FWYYiXVaRAyRyKSpFLURbJQpbBOLfDUfqpEf6TM/KNI3
cPL2rMOVbzPOL39GdjUTKGW+KyFwFef39GLfr7KQl3D68ilvfRmh3UQR6HCZTXiUSUbNs7haqwS9
54VCckWGpZ3H1W+XklUAeBfbt1wHl2Sb1EA4hw7nKkxUuOXmCOFajHCm7Ya0jjmT6uEL/GhnKPIj
a9KHzRFvhL/ELmhjlkeQehxPZMIUNDZzx5d99SvWz2+GGqFeZzsd8+/jXzGMk1RkFGf9Gq8AHPM5
gjmT2+frV1TnIXnMiqhgPDFM3H0SveLuPu3deGz7ERE/xb1vg3DwuH3el93qie1VckMW3H44QKME
rM6AKbNz2x3RdYChKNsPjIgMj0JP7TEDYJodnacB7IaGKqtIrzg/AdbkwvnmT9dC8iV72yj2w81T
CbZ1DnrcHoU2/Kc4SkGSyv8XLlvQRxGmv7NBbDWEnTUJ+aJLc7AMKxc2df7e7aJzxTRGcR8H0SWi
qaDQFN4vtMPQQAE9OtkrlYoBW2WF2dfSpD8GmM6+7cgnwUNwwt+BKtDoXd0XJG7nTPOE8lzSYTU3
rBcEJG0oQZ7mSO6u5uDARc/eXL6q4mtoXadMEli/kzoqniQAH/f4OgZ9WhxX1Q8iGr1Nyf92F8Vk
ePz0ikInwiOsbyMrp3iXvKbcWMMnl3MQ56FaU70JYysKo8WDc9mFEhVUaxI/3daayoSTiW+tIWyG
EYPCU7wrvqKcTWRlJFwR5aL4Y8E50yTmOljP0bPmfZDAypVnXCr9NWatK6rzBvIdBhk4cJp1jjab
nkeIj5joGSiochHax7iIc+7qFoOUoUoVeD44dZDDAoDAsrcgQEv/XURdiue0XIs2MdK16rQC/gGK
+K2DqYUfChAdl2ZLH1JGZgjbjUHYYMh8dKNithUQCIOop79+6CVld9XXQEFWHPnUCwMK/l7Xfox9
js66ukszt2ApGJwwCfbkz1yc5qqT980uIznS9kIXzOleMgak8xRmQwwl1LXohvk2Kmza1Mjxq2ij
z8Ng5PZrneQDGyMwaqQOjFzTXeUUH+EjFKWU/3peZE7LQ/lSnK3Z2mpLXYP04De0bazmTlPPpHX8
Z0b3xh2whD3tgX8c0ZwDdgUmqMmnnoLPJDzM/p8Rn210Zwq9rnQHRZX7P88jdkfcT4gDgdejHIUs
lg1Cn5VlhHvhIBUH6Vtdk+6z1yq+PvdjM0u6Qe4NAb0nlMWJYoKjhyeqneZTTE79LnZ5Pd902MaU
8R94cUEKRzGWlDKK2gsy6TgwcUOL6DR0ufk6z6zWqZjsNm1CFC2nbL/6vm79KxenYdImIrDCJJiI
KGYIrXaakujQ0d6xIDr4S/B5jbejEAf6Lk76t0l9k5oPwCbNDdORO5Zo2lkS+uJETo78Q2TCwCfv
YFfwl/Z1uwx4/ZAQe5vzYBG8bW28RSGQP+X6khZrXL8EzoeKPFMeOCPpZUQRoOY36MGAuNGdaFp2
YP01VEAGvM6yqVTdiucSZUtHjJEXM3xIoxnjQIjIIW5LSH/X54gjaHzWMkRh7fyPSoJL+JeiwDva
YQ8SVB/dwbH/OTYszjoQsRFvuKCEKkHKroHVIABNWtTEEVHBe+kWvl6FE0PSBYJVgtGz2NsAosNW
dd6HXyk8aGa4BxY17zPEjpFHraXqthz/o3Mytd33p3s3FarMTIPgincuKcPg38OK0HE2T3J0T9f6
sPmBgsWCVlyaMybz0XJ2l6iXoF7uNCrPcq3qb/gE5U1DdeqQgVvIyhpL31smnGIgENLKXkrXLFEH
07oJCkl2sPNMyWJElNANVS468mzINCMEG2OYefp9z1W3M3iBGCSnpL74NWR5wdbvl7HowdOznRka
IpoOVy8ESqeuSOqe9nUjAY+Ce5NHZAXcQi4aYccHpUrj54Kqxi+FpBKsRqxPS/L+5SBJ2W+X6I6+
+sQ//wJi+lkOr+Qvf2FcPABbmXBtUVageo0h0+ggrCxEjJbc+8cdm+HoKI4mQFquOgVFqGuAn8Ck
Op1FHGPVgHdbpluEshES4ZfdOjbOMrI/GBdrA/30BXHY4wGj3JgUTQLpY8QgO+VZUbYWDYFaAc6E
LvhDFgQgzVrN06cgCHsesnZiQsPBcvxLWaSIMxTw0Vo3OvRGuiilnep1kbSlxTxKBx9bSItcxxEd
2BNvhUe5nd3jhTRxIPfTSBEOz4cEB784C0FpArlPWIJvORq4DoXvV4rdyANUaeTM2d8WWocpX6Io
sMXHgke4rOxYxjpGRnzHuKIUUjwnKrF7GqNHXDTM9vAcR/IbF3SH6EGYvahmIsLKTwkrSspyzDxo
mwV/RKjx8jALbX+/U8e9bZb3Yvctur3RL7XHj2HyVeMw1MFgi43Kauq3jF3ZWRutz8qSZzT3u/FX
pDbeqHDwFqYBbtNgc4eGXpLY7Dzdd0XdPAXRTVCzKOlKzviP599sfTqKChOo79oLGTdV+yoSHlPO
UZ3ccLbNllNXJxsnHFyv7abz4p0k9tIDqb0IdcoknoxJL2bnR1JsTHcHBO8dROGje9Yf5IYGxWAJ
GvU1TfThqIpPne/c/bUa9rXsMQq5YvJPGm8qWZ7dSBOXOwxPf9U9acX73Rfo+P9czTpOCjNCZ7CY
dD6WP2xAnCBHjdAU/86WlolhcikcYWBPtNV5MpwkzqF0LKtZuP64h95AxbdhMsNcGTYhFcoaWL3U
E63EruO1MD8S21C3liwxjCdQ3+9gL+4Ny4zOQ3kT6vQGosAo4ddYzq0tWAtOg646zFBqAKWDpB32
XRGMClc+ZWL96avPyhI4LZ6A/3KYIaCn0R1+E/Lk1gQ78OLroaezprLbFziP5RiIydw158R94Nsz
SuN3aV0IZl1P48Vb8rw92nrt9mBkXch9Fvh4Ypwqi0dzt7Bl5GNgAi5TENk5nvXU651atzVoySut
Yp8D6HUivwK+WldkJzOxh0JbDW0xsrgSL1YOs1zQu5Z2LN1kZ6KyuDgN5Kn1YZR+zvRFdQ7p2pGe
7WwH9p8o9wJbXr3ZW0SnYXe5ZB18ygY6WF//GFAvKEGY26yF9cC5E8XT7De5Jp1Rh/zcYMvmj5TU
bTlJpKENbxmjfHDDXEZ9zp5Pd275zEQodlrw5u7Qj1fRHAuOGoOUNsS7qmestiJoPuNET3Xwd043
EhrxMe9UAAwx0rJZIvOVYK94g/+txPgdl2C898AemK1rViHJ/9CCeIZDbM2zgrVHOOXcKhCRAZGe
ytb41NSToKg1axQL8FPp3pngcSnbte+FliEQG3o5lXjRPX477ZXZqj6Q45IRhD31OqnuEnlAsrA+
Uf8FLzbkZrZIwAn9nwO1rrLLGG7VeykbneWFerv7nWuqHnhta192GMfv8x752gv8CvxMOXfRzuyD
QareOUZr2RhlF623/m4rTibntmdzLeptP68HW/i6w11Xl+84yQ2dCe34xY+9MYWKdb+FAqH2qMMJ
dCGKPCgxSbIvc4B+asgCc32C/6UbQDLq+bkbThJYe4yBtl4VROw7dlV+qA4pkgqa9SeWTo370Pmf
goq/rmkPdthH5NMjuQJ+i6+zKsAXaIQ0Dma1iYReAu3USSwaCogWeyAtPx8tQgEB7+iLd1RfOZxT
OZg7aZHUMQBKsw3q+YGN8+SmC6urRHRm+0jqxQedFVXi3i34lEuHTdTGtZAsy9wHUIxsM8Zh3Gq5
ZRt+f51tDDb48Zfu2E2ipDo7FfBh+WAvhQL9ytFhLgQ7Re1a7fGnyXAZ8cmJyTEwKVJ30OcpPA9W
kZ8L7mThi6SyAXXC9WGcZeOMol/4wQ3mJehfxzfoKsdu9vmJ34eDFjx6L7kHQ3OP2ibIOI3XTlF3
zeaIhTkT5wVKEknrErgKYol1wZCvTsTSnYCWHrBkMExqYgXXrvG5BuKWnr2HjFN1X0Pwzxuc/UPK
/CnbjWCD0vj3mV511x0YwpIzt9X5nCGtutskYCXTwwJmiaqN/DpPKvlCwU6MasSbDRPqRETZXR0q
QNk/6pYcGcTGlQO5mrzl5cm4CZ7zypjQLUnSrK1AmKW+Y2/2QerePjxVvxelUS5z3AXaOA7Nymlg
of+t/OI3TbuETaX/gus+lVe/T24iMs9Zxx1sjfjwFD8VW2j/VevIOiqDZEh3rLOE60wxsCEoWVzq
o2d6rh7//Gx36QA5T93Np/03IBFppdQRk3jklQwnQfhasW8I4cmefynSgFdT3GFaNJzMWCDy5rRV
xvIjG/nMSq1fnXZh2nVTJjHZENqVSHSHh9oiCu5av3tp/lrkKNTQy4hr203yeYB8r504fmuwtxfK
7oKbzymsmiuMasAwIeuR8GVIdAOXjlv6sHA3nT2+xqXcO54VMDoYFC8DFPNMfNy4PtngoXF56P5q
Hryi8u0D4vKJZb7tgateBAFg0LfJp+TPx0R56AEsotlQAlPTvSuCJ3/wbjUX55kG9rlCfumXpLty
SQo0UDiTciqi03y4UCvMf1i77NoGIGlBvQClphHrgLDsvoM0p88ebcSzwTrR1BY/LivGlkzw/fpg
fnyBxiAWrAJfIYhLcSwua1bNtlQz05G0VnmOMB/wQchD1uE1LKdVgksyWxPINBlNP2Pdfni1P1QM
Qb/qVHNDHFZWNHlaRUREm/HAcudXpPEu5C3pkki7yBnHGAlYZdwquoIYXRcqtqXx9C3l1ySKQIgG
kuszEBY5lWB/VKHZsc1wlQY+sJ+ifCaEWvt9PRhjLZOlHDGyG5JBYOlbBVnGcO6OAhssLdbc0yDi
D31hmrLoqbkn9Tfg7/IMAx4e0fqutyq26XMt75M2iycp7yIjKgtuyKAKwr7AdZolFN0rfJQICRyD
oaQKseRzAv36ZmtMJlcz9573tmCCQbnwEcXjen/Ak3jLryXzOLnGd1N+rMIZa+DRYxRQOgl9b/MA
cz1xRM7z26IvADpV4z/kWxqg/DFV/cAclcIJvQHj//yzUPxwGWhiFAIioi9NtNHq0HR0eFyMdszM
Mefi2zPSlWohF5r0J5GYZyVVaJ0IlNt3MQCOep0b59lBnXl5qDxMJ2ExR4yiqBqJEfJskiYqIA7F
LUqy+Uv4qZPe3QHH5tudDsPGLcixAOSIcst43soMCud/XuFRdx3h0iemGY1x8d5JT/GtNB38ZhMJ
67Omfrs40Agz3E5u62FwG/GImhX5MeAjVrpMakss1Xs3sYnQeeAtl+KCKoKkq9RV7krNEBc98HLj
mLoH5odTGgMWQc6oXaPqj+aZV0GFCeSLJ2ulyMPzeJorYeQVBYZApcDjVDK5UkR6qM9fh4Qy+tgq
+h6PadMiBUBn51FNUuo2hdwo6tG0gRcio438DX2r8yVPSIVFCPF788E8hDWebMYocZ4a6Qs9D3p6
60fP1WmaJmI2mQ2p6CzcSoPNEsdS+njB6+ust/nFKey/nwN7zgoL7cUTeDhs4jwQqe1C83TwLU0A
KEje6F+vP5aW44ioT3JTqJMtGEouv9G8c1RixtkcsOsPmjw8rzNZF6QTH+H9aR6k/ih6ImPAvusu
P6HPLv8lavAJDBGw5+mP53aNY+wBMfoW9nAxcw5YlSCG+6n9v74Jl/vi69ZluoYA7Whhy4xmV5TG
6qR9kKK6sFnwfWcLV1wlmB80VpJxEuD3cTjxlB2ECF8kVVLix4b6UAT1CjbD6+YJFTRYYfFWMU4y
/FqG3iZigbccMeGZa0p8xCN/UqeKl1LaIM7Y8HLDhVNqGxUT78u/rlXy7TLBT59r2SKHrHQYndvu
Q4EqBDkxlCVO/BJW1yQyAzgtNlGN96kzGplRi6uP1HWZkln5mo0QV7DygJU7nnyhWrAmweXllvFI
wHN9TmtATCQiEYjmv3KWpdHWQFDOgJy9XbyrR4YKiPpj0Mp4jkJGmOtgyDFCccKRVYMp4ohwOAGx
ck/Lxhmkg0AA/jnY4gb2dkoYvFfnwM783Xh0E4xv5siWpze2vA3VkiVQ98aUJcPcqd//d1pydm/F
Td5wDGWp2vG5ml+AgJ3Eew3dqv6EYuMrhEmPs1ycJkZTxDescyoXDVlnj3iAHvNwHfrboYdfKZ5i
X9iJwO652Ph/VNKFiFqGNAgJLww98GW++yqptVHNr2tGggC0FD3CJSWgN5IBHP6sOjR6Lu2NaN88
IwttOdZ1/ODyCAKhgWJbqZ5IHQwgY0LDdYxX4QdQRs8ws0nvwyU3l+LRQPGEVpioPLEIHjSp9iu6
8EBriIJxGNgZmwL4kN6+X+C3hzXxqf8NFyIBGW8vdIAJBp7aNxuxjW86sDfnVUCcZ6XdSGdumhfB
RihNSMB3neuZqjiMLqu4mMi60qkHCVmre2HwLzgxh5dvfVwLbxmy12eFcfgjrZQmZgkv+7t2YqnU
c/A5g16DwFmRe6jPjAMbdQHd/25tputoT6OQGzH21eGxbDBFLIZIW+rTGj9umzBpi8MTGnNcQJXF
Em2kf7pk1d3pIOghaxT9WmwcM6YBnIQuXtTOnAe7VHKn+VMbdkzM6ML8PPBmBl9REy/OXnKEycfq
J8q0Cgu7DFXIsCIQNUWw9nV0yi+bsHSZ7ggVFZeFD0VzVg4miIr7pGJybdQSxm/TwZz8N956/gLO
Dkn7ZhbfrdxY6FlMhSypco9dlKoRLPSyNtdMQm4AnT6iEVDAdIOkEO0Th3beHhgNNJ3m6BmLvMnj
2IXMlDYq5ntZP4XqmleycHhnwAc3CL/AYh/sqRi/5O2kCW1aerXDSCnJ0dD8sXTulGf/jrxuyI4U
M4JYMgu7NSoBPuX85HgtxgF5q93kzZz/qF4MOIDGLsjufY83Cla8gs7xDsuxCUkEAXV5lMcbDxy5
TpcUMQdwjryWZBl6KcTl/q9MEPhWzm/VVQfnrO0PvPoO9dA96LfQBr6xIYaPafG+bQXc6gUT6tN8
iUt6ZT86dY6EKvdkLuguKzZGNTmsEqOFoBCYjayBB/cnyVkdvoPPUJUjONtYTx8OwgrYug6w/8Ue
yn9iwdWSHBtgam/+iR5LZ1+LZeCz0+jIYjXpmjKK5nTorv2QIteFmIZiB+MjPygtOw0yiXmyZ0P9
6iOF6zf5WsGaM16e6SYuH35cuBkVdO3EnYnbRKpnxBWnHkgpc01aWqu3h7gdPlFyfoPgobW/X4DL
36wvxmFbWjBb+SeftF+Q+7vxp9vZCojoL0wvgNwf7sUp0AaLCFOQwjRknFAnYX2eBYVQhYUx1Lmq
hKIOZGdt/AFoGIVarQB5iQJKBawZsytxzsXqWDetsVvsTNSWsrfR3I3EwoFnMPyOD42gl8H3SZI0
a7/7cl/BZCl2+s+hH74UbMg/qdXRXWhTF2YEMM2BiabVidebAzO7IQfl0tuzCYAmEv/mrBvW56xd
bmY5fZJx1aye3wd8WP+wH+3Bp9Wo66XuzJvVvA/gYgjSPokKpEfyqrT8rZpFkcnqzwzm5eKHPLGh
87j1tio1a2GkgkJr0/qk9DK/n5BwzKWPBBlUV4Vpehdt0gXjnPe7WmaPzVCf+cdqDnGpbdVF8T8l
ST+QiEI3O0OU5V6e3lYUEhfvpT4Fb51G7583rgrQq2OUM13xZiwg31sO6SC1L6gdfSCy+dow5VPw
0G81zonv5m3V6FlU9xXnwb9OEcInUL5EN+IDLeK1/FV+UiEUEN0abh7vA5A9d/z3d73DvvjFxXiJ
3eZb5YvxMENDGW5yzLsaXoZjF2XtgeWqTZEmdG0HwE9u/M8/fB3L7G5YYlfmP08noyi7sO4B9K+2
li7LwrJsf+10FPa/ZFTvSxAbX3zHzzJ8nSPgRF5hBOUUy9GJuPbEzTv46TLY7aL9CRqFMvEUBEZW
10FfaIf01CZt7RIUr4v5LWzX5NU/nbCeTN1fppRi7caZuXo+v/OB5ValYkLkbxQJEwsqjbcDPTwk
6LEv9nfWIRubRP8t9xtxWTbsANXXFVDjG8BnXElOVp1uThWtOf+3djneYK6S4skkO4WTTvPNusBe
vNjAFQIgLoJt3bc/99ao3p6xgUSbLSYV+Vdk/T+4/5eU1C+UajTMu7bOdIMfIICV07Lv/6sDnOlg
Dkq/X8rpwxvVB9sp7kv/YDizjE8AeoHoSSguOXyRf6lFUZn7MApssBk8wpFlpPcIe++39CpP/inc
qDAqjFYs0b86K0RZyOs8ordfRaHdbquda8AkzLaC5LztxD1YKu0LGqtHBEbcSRA3oFPfwtEfLBEr
ZCZBwUsIwVzZ+0B8lN8vbfK7dMdCZ/7byCSex/V2jZOMSwnB+D8IkE+X/Ii5fp6pzaHyhURj1Tul
SkuyGJWVJhVLmaPGqgzcP29Ea0rqJzf1qP7Ye+yiVrZE2J9sE7R1xfZ6B/es2mK+jlS9z/8WK1EL
4AMSVs545PRIjIOK1apv/Ligo8oWnkipGi+85KyQqh2W/Yt7z07i5aWQ4GCrcubY29FvGirutC4d
yT5eEGOMTurgzz9uMmRtoMIVAEBca6nY3ONx2Pro2zsLC0Hgx8bigUYhGDmAeFQJ0TBaoAJh+P0C
eo8aSSaFE33CnwwFolR86j3w6ibq2zdb+C3JSbOF64ZTYYogGbxzNadxRussjo+htxqtsjdSxkbg
9JSE9HWquKf+bkXctP2YzTu3G8YBsFGT/BdknAXa/QyBb0kuJ4GMg00nqVuxL9/h0wBVeB9n9Bgs
dhs1qWz/WXYrKEJHocZBsxqSFqsh2dbENUeCVmAskjKZdO5mBwC20A/RNzBtmOVKLnMS4UEddeVG
cjHUbx00qd7iqQ0j1YKbO2EfM0Cm+oJJsXn2MwLoauMzPSuKq9KxZ0UiawgItV7unr9yva/HZr5j
vNOYqU8Ns56DjDg0uCRncZ9Lps8oezGMuYS84nezT11IXNAdIm/s1iI5/t6V53c4894XvZNL1occ
6UBjJTMfy3/S1ClkR8ZJH1rcLjzShQyibeWO3cdX62wAwwc6nDp5OtwgvmZQtpEjmkOYATXJRnnZ
3j0CcBqGCicYuYKfsOADN2W+5gYIEzq3VpFTURz68h+zfUTeV2zx3mWX6BeFWIPdI5/crbzUALca
/dI4yN06B++vyDrp1/mx/6evIvyITBIjsTVPPcnrvwrbbRgkDjb73ZnzE+8BLryENwq9bz5xfJql
fdJgzRKE5dTUvFvn1CeNDSZpbCSMJFF+E8t32bCzBV6VblfeDlX5JvSY+0iGReSPrT4EJoQHJbI4
r+juN1Yw7NxYET3ncru7erleHXYJd/tw34EmgYWB02ve/amUvyXxVYgspjkjEuFvaD3jNbYKUV+w
Ihs2mjqQ43mp8epCQ8ZzbEiUb4p5VT74U2CUmGm/ZvnhlXMQItPJ/taqweoMCse/f10S0xGsPiyg
VC4f/whX/zfMB1fm83tg5G3sVO0DvGrWAag4UHESwAhdOXnKby9+VhuL+o4pBpFX2WxtrRMsSRhX
2exB78F1JGQbQGz+RAYpvY8X9Ib8/5DJykzWncxxqbwvLMahFw38IkDOdw1RMWJcd5LQc2VAgQQk
38n42Yg0WDueXh4V2PDIlzMVXBLvXXpNI8Sx5yABMVSD/4Nt2mc21HbDFVTQ+s8FLT4NMs6Z88mc
ApHtniBXAwASDomGaKN+b4yLyPCp3bZvaDaM6fCFOZ1DxG0QvSP675TU/jOwhqF0O/QjNLxZYJAH
go7hvIaDfrbjeYvWQGDczMfVEYUfe7cEq9BpO6k0ugyx+22U+d38gLGqPBWsARU1CcA1FlRTafQO
nAcXkn98vhBTNcCEUx0BYI5UstXL/pTCISvP+rGLwFsAY2Xv61o7wq+csYjfLuafF0dQDNGH4Yas
oUAc4TVHIitikBejFzvnQOvBfN2SXiA16sg6i88Xvg8K+8C7zmm3DTzQO3cGqJuXIZc78YdgJ77s
Gsj9Quy0BiLvyYCQQDrKNctvHg25ZIZeQK9FUIG0/bZuW7ZR/PJA0TcmfEGcHsjs+wLY2jzFB8MN
QBdS3+azrGDlpkFe6o1FmoOPfqV+WkNOoYJEhJ33g7BK9dAUk0g2U6iYGjzO2K/ZlITDwnoHy8IW
luxo+Lsfly2yB8VFsV6mUL7E60jHzqR1gj4VGPGvtdGMusd3ZyzLaLi6kd5DtGmKO4XgGcZh0JyE
OoUMVa2Q0e9t9xsI9r21aqjt8g4hUGtCMEkgve42EmfZIcV3FF+xGTGVW+yvseQDV+hxOM/MYFtH
BKs5FE5odCDDZxtoWsSMOsThSTvhs2ruFfx1IoFRrhK16WS+2700kou5XML2wJB0+WFmgYk9P00u
WaEFCGAW9LDdWHXpST8yU3MOEiWoQOTAjElweuByNy5Vuw1TwnWS2ImagwWWfrHN/pIsHwYfuGyG
W9rDHaGuUKtRToX5NQTpFmuwMiClmyame3cdWjDEg/A7E8ypV9iyqpUqhK5fyVEPPvKbEx+G287q
Kh0OfZ5Nl4wErVuW3j2BMR94KIrCIQHWa6jQdLZuCVIIF1YStBHWpaZjvLTXUzcFT3juZRoNpNrg
BgQRLY4+mdiCBV8fxWS74rQTYb4+gbVV3MNNy7GVyzylVBv0RFCD8Ay50LaIVmcu6jYnmSjNb74X
W+BEku7M7erI3V8KhheAxiCY4NRJgZTyUNtd5iCwM6UGlw6JquhnhLWdr3E+bfjONNvmLwYl8LaR
s2e2Wzl3+QbEnHILxQm1G/5Ph91bL6PTsvqHyzYfi8b81DyQqm6RcsIktiAFFKn7Pa6r9Ud1GxRg
3NUElArFRXZiAgPyxMgDdjjgP7NwpV8hXDc6ik7NhB8cGikg8teNFjynSyMK1pjCNbataLsM9Hjg
qdMsnjoEqjh7W2+wYpuxCshArPwV8zfmx0oTl/LR8nqHQ3CV1cx8JHRcprs8gRS5ilYL5DrVGM5/
11Yq2trFL8M55Iua93CIbbOFYE24e4gX6P7knqqC7UA3dGHDDt/A64vdExuJnjOeyzXjZC2zUFeh
p7ovHgPi/cTgChTg1vGcGdyCFLDxMyQPEdsfs4jG8b9LgQAOmbRqcFzerfnTZa9b7wp5KV/vUIXx
JvFa+i6p37F7aNXqkmCSSjJF5fx3/U4uSmWultSaVneM4SYw8aQ8+y214Rup+JxS5eqB+TOKSSb+
W9GOH9JLb9Qa+Aqw493AdtLgBHAdpudVQhhmJLYUM2PTrZBKBrI+1GbAQksdLX2RHC5yCAcGbuy0
UfwX4GZPsIzlDlPtCEUOUW2EwrA7CPtRPLSP5cc1NKUeGOzU01b1Dw8UIrwzlHcJXA+V75zsEz7R
OBzm4FBMjlspedKY9z3Uq9I/Rt22O0wNuozS2GcBGP2esesBl29IXQotsTBWXHixhd6VRivZTs+d
1HBp3Lu9JwVbPZfkoxCuHuK6b2mjdnygB/kG2PteFij3DgC9BRRcP+NGEW6xd8CbtMXoz0kK6yzJ
DnNQq2e6WzgdA4zXfn+qqRrkCeVfxx2hpxgritYv+luHzB0ffT8w/mgfWhxVFpPYhg0EkBvt2StZ
vHoaUxlvmfsWXgmY402xG8SNO0UeuAjcPA/2sHPPiwO+KhirIAn3kRZ4fh1PVmhNRm77GblCnl0I
Yc0cRqjSPAGvG5FdKNQLFmuwKP8D1lygvIRye+cXzqhqgjCHKQjL4aydtkHDWEryoI/badPgyVH3
gTNpddaz670ztMXP4jheUfOl7uijzVDf3es8RDFIvKN8EVKZStsRxc5gFaUQUNkDqG6SBF+efXfa
MmwSgN7ZvDZrlKLEdNQjQMUwd2/7V/sAFaSIbWqkORM9210+vOp1bH920pAmBKOeCGLbOAxRq1qP
9mD713Gqp9L1Nk3r2vmvczp6z9zpJUPjRmxkoHph6t/rTOD47/nB+YMwIhYnYxoQTj4Ag4UgmQqW
OEEVjbEC58mRBLrFv/9pL3CGAmPKnncMide+dHaS5dLwDMu9dT21T9rxx7V0WC737UgEzBCIcUz8
mdH84JTq4ZLAiD+SD6+iG/1pgzyLBo9Cvpfv4MESuOuWoO7eiIRas/7M7NC9JJ3w2fgL6+X4KOTi
d03LreyLFGoXJ2qezPthz1UUPonkZd2MiB9eAI4p/UNJokUoj08IywHAntsvWuCIHhMoPwgv6Fiv
ZE1YRu/Oi/x6ftFuTW696tvol/JPaxy+oLMuLvs4OhfD/o6wk1/FAZzIlo3Ye55ayiyDN+jhZ/MX
tHhiUnCIPG763N1E3kBPIPLDbjliu1B3cW7G3oRpr/mNjANKKY+7S+x/cpK/6XCQ7MRF29CHcQ10
6i8qBAoi4DZWhZxe4vA91jq9DhtYTawA9ezq8BB9AIHxioMwcx9U68ODW3BKS++yKhlRX2EFpPQ2
HichXgjOWMkYFiS5VePLQjcjKXic57eFDtNNbIXJAnnYQ1l8zqkGQS/I8KTYRIYmVtNhDlAG2qNU
GPO0SvsWGRmoFLeqdt6qVRcj3UWT+D3l2ovUhuLVyYoHlKgo05/J9imTugGoVybnUU4kMyYJygUG
xh2kXkB2gtYnElpk19VYE2yeypkk6x/AiI4WeBV//kLXjjJ+3A/kOxie4024udXcX5l7vXAfHkeR
f8BjLUUThX3FKES71jq01SdCmmlURj+WGAt0D+xCuT374ZYoHQDHnJZjkxq1dYKl2j44cQN9+wNQ
Rx3KHeLaT+4jGdYzv3aKBT3WUyf5ENWeLyNnKdIR++RW/kLufmTaoiizOTZ3B2pOyRLVPMjFkWkV
oJZQKl3A4ILy8CzGwATmowMgKUdS+CnnLiGlEDUeOaEdQgibcbLBIvCeFCUGMAn+Ji2+78B5d5VL
/MSl8+NxBKO5qAT8MNlZWd6jDvYFUFxnvgft0nhGGpuhLshJpE8qPuZx/1QhJYX19JsnSnHobbXQ
g8w3//MoyNFD/b92tLaN8nCh5X17WLZF/w0zGMhCiCTtixJmxxj/NgUucSJrv2nffl18xF7d8eGw
XkAETmMRIdxQYkgQ+IkdqDLGRBqz1UHqwJ5xYhxoF5HK3N291Lgc3+5hJdJLl0N1Z35hExzbfWK8
pRvVphgOsip37abalgQSL+VhX4Mf+sIgH0Dyd+viHd+TzNaLJJR1JkUsa0MmIdTwvsX9CpmVmg6a
fKFhnqCJ56fO22PRjNj7WrJO3p8kbzf20KOlEO6vujxaiO5twNIAJ/HP+Fq7byDqNNm6OHUE+vao
2NSm8kfsGHr61MzPod5XNFZEjxWvFuMc2v178W58waNhP752FuXEM8WFQkzhVmov3qLxTSdVz0Lo
KKNqTRzl6M9yKqtmjZDoQAcp+ORwrgjmQaN/GYNpb9VOqAK1JlVOiUlv6Bf6H7hcr77bCa137S/I
xKXj9QypI6f4hmExzfQaJ+oODiutWDUM7uM3i9SiaXmjnYlUNvq7WA+71NL4scA3zP7RNAi6R8Rk
sfzBRXrfXVJf8z2wRo0umUpBuyBfEZ7HQjTvMz07RL8eEueS/ANDQ32+shiH66ZyMC0FbM0xtW/D
1e5oCyQNF0qYclVYdoS7r4Myj4ZuBpJCmhdL3btQEjHZ0+YTpmuNbXz8bs5hZ/RA0J/cShpmE7z7
3kkkZApbNx+Lfn2Y7YX+l58/HzlUgGOTN1akphVx/FSPMV/kevN+isJ5TvKPJezJ2V2pQzucJhvC
IIas8IB/n8FpTwzd7owisfHko0l+LAUNz6DKT478CeXfU/oaGSxMNHjK0ytEaDN0oFXsy/oMNEbp
CVUu5Rx+NymjNNdr820ESTMbMpnB+K701N4dY1yJmm/b8MRonjSD5D0fU52Rz/Ka/XMOm0DHM/bg
yMavZowwWIezm9GOZhvNe+lwG6+gM0dhnpXUbkNihKFbNPXsu7jEb9QbrVCLOsVbPdtK6Gsh9R+H
F8wjQOioARBcZZU6RVAry1/sAKvQn6fZcz4dB2wEPB/4cNZKe/PMZiXNKfekubAiZZXxLin4+/xp
Wq8FVPhyQ/HDqwyM0mLOWkNHUByKEsUH1O4PB5XOSUBWP9k+piw24Ha+hAehqiJQXwD3WDLQoFLm
rK2WcxI+BBPCkeNEEr/Ph+jGX4MAgPELGB19a+GGUDdWeLsnRSPmEnI0VNtzChz6D+McNQXMY2V6
PNaEsY1OzDwCat4RREI244F5lnUVUpUuiQ5kruMSbeQck3Iioal0NXP+Ctus0yPEd23QSjKjJLCv
pnltnDk35xftVINYTJm3w3dTCJcQHYbJwtZGmMgBv73P2tXTvijnGk1u1HxvseLetmJMysVB6N6T
BZRxUS1GRCmZMYVb+Co3e0v/t6OocfqyfIawJnv+lyjAhn3kT8CZhCPvoJE7qr3yzc2Oh+ZmSFaO
/aB7706ZnBLm1R619zWoHyVXIO/FLLAnolAIFRm5n4/KTeWH4B2HE0Dgl2/gLqT3ujJbEzUUG/GT
lDSCkApWGubHPUsuAZ3QWmvGnnK0uCMF0KSTD0USbsa5FbaLyBahVL06jtwwA1atzggfpBYrdd6h
6V3L9pGRf6Ln2L1+pruJICO1A0HajOlD/t5jPTHp7I2cQm2kjLtwSJosZPlzBcG6a1o6EVB7hKE4
e1t09fUFNGhLwC7eBmIRMstatKkj1DwNqruHErs8JHgybKLTesqieJkv6UYlPl85iYXXUJLN0wC4
ob765mT8X3ekevacgjDbf2u1hUtA+aKqcQhbDD7aRYcTPTV0TPymLZbBUxM1hXamTgMS8iMULMGD
p2zpm/D+KJC9ahjkGwcZ1GNxj3H/Ati2CydxMgXNsa9cGMZ58dUjNIMHJzS5UZr1iOutlgZV/mfS
bKlqfUApUi9A0+F2C36uv52+1WS8tamtfboKDe+g1e8OgFEtvKawpMaqSpEMXlTWM9ZYEMROj1zv
4nQiG9/mXs5qf6Cfu1pqea26KzGwwWXWt7oia3mnRmxDxQ78wjegiGjQLIR3FC7KxCMX7WTuUD13
S8ZMQTzOGDdeizVD3XLx0SD7jpnF81gREymUU+TJAqX9U7gcflVz13HaPyjfhHBI+TQ3LlUlYBAI
247kNoqqXIWolCXWV3znSOdxzU2CtY3AWRULij1R9CSVT4ehwyeHyhvgNBHVXSFw12co+IH/lshn
qXaxN8pbO1qEoR4Gr26/kKZ9qHHVmJKxBAHeoiB0h7a5OV61wUZoedMZHFirvL4sESYQNW5sN3fN
poMgsFtm16ZOd2uEMv/2ZWzHr0MsmqEYOnK7XTWACEc8xl2tAMRy6iO058d83kZhdQlGeONceuXp
9QgeaG4bM8cXbqk4n1RwBu7rfST+B+7LHg9CNrcKpABSNDAYPJ3uvrrpaZJCHudstuR8ic3db5DZ
ZdOuBuHnrfRoQjdmZfNOaAHuaL0Q5DisQFokRl/UX6Egmp4DTZeSJTlJRXBzDerUxSKk+l15nG5Z
5/62KOvhhw==

`protect end_protected

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinx_2016_05", key_method="rsa"
`protect key_block
muLdAs+6DLCdYRSINX4VOA1B5H9iTi5SETE+T/1nVkohmwnwUHbTwwbczcmYlFDHY/h+ekTQO8Up
qF1cwbq4Y+XNHdI1uossYmLDqgVDZuWb840UndgZbrmOC70HzURFtmRdyOMJ6IaEGNy5aVBXdAH7
8I8hYSFPihrUgfc4zgFzigzP32GaUgf6ZpUabaj/matQmeEYfo0HGrzIOeRbqoxwSctvM4oRoB7T
L8x0APebhZaAkP56JheZfz1DSIXYogyyV/J3nFvNrtHywYoRfx0bYP11R+/eAGZcP2BolRQBlCZM
umFb6QhlQeI/BmoBc1erjbG7ITYV18yggYfucA==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
TeclWLoUVF6I5YBon5mC1tOobFp31aMBjdm23z3eReaqI4qiI/Nh4chYN6KSTBd24o4C0RHqxr7z
sKYAaaEnV5GfHalE+4Xg0eoxhOiiyQZcEWm5suB4S+sLx/Fmx7guJTRzBM0N6WrzaNO2uPHVlMRu
eCQQYRKNbUNdEd0T0C/VyHxASPMcVv89d/LM9as6Fsp5Wkbe4kg6s0P5+lTdS3a+G5RLrU3gpOs1
yL7sA1hD87JuZfy89Pr44DG0fdEEU/Kj6if2QP1FNhyXcMfpgbEodJzQG2pI5B35dAfE4wBApwkY
op+OsqGCSfn5KoTXqtvZSVB121HVbRsuvj371A==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2019_02", key_method="rsa"
`protect key_block
S2j2uvys1VHxCDwtsOd+w1ovrekX6JpH8dymleLN11qQPDGZRSkAn0TBfgaYR3gssdCK7BEsO968
CJ9y/78lYH6TDN518uNcw6v/RlCI6Ynz4wsPnbgqtmGhI2R8VQXo5GHwpvzSzuG8M45TvtxDdfPU
6IoEvaVUQwru04JZJYbIN4FfTl5OVuvvi12D3i8zs5y0XWHee31ojkpU4R7a2RBJA9bOodgP4jSn
7303kgZvQTQjDgaCficFZUqO2n45ScIJ1lbPrXV64jKqaeBwSo6DrPyEMVN3rYTEP74OjDldsyPM
QfqOwz1Nz2eK1VC32/JCjQIAsL1rEPw6d/S0EA==

`protect encoding=(enctype="base64", line_length=76, bytes=1488)
`protect data_method="aes256-cbc"
`protect data_block
3kWvzlZp2S3JWsE2VXAYFDj8g3y5GnEmWSX10qLHjs49e78fG3ax7g74QydJxI1u8NRGmlLGxnPq
Yo+2IQRk3jXQpOo+MCDErnxsX/7p4+uU0DFE5qRxjTeagyvLNHiriHUSf9chW7FagP65y1W9PNIR
+527LwJy1dEG41pQoboFLCwhBOel2pNm9gMwPF/7taaubzv1eHVz8r95Y216SDyNEihx5Xgq1nnO
19PMD8r9KcIAIqTB2FvKYIqs+y9QpyZRFwLqC/bnsFgNOyzhyZG5EyfpZgaJpWtg+k+LFj6d8K/b
HfrGot22FITyl56QEp4+OS7txjrMlht0+RsdcxtBdDp8GgAKFJYABBlyhVKd5jkpLqgl0qhrajqF
4IYbrRoyVnqQu3jhrcfzhBuAvNz6vsxB9o60ycdOXQ5NMYdeLci7LoS8EVUvju9XrkTg0afikGCt
ndZSLacbLHx86IfPeuwVXX6lIIb73TwJgwgmpmXsFV9Tjmy7VB7T/aRBCNcX2O+fz7P5M/RbbPjC
DVJc5+7Fj/NpKS4zH0Bq+H1I+cTEQcQzQLTYuoBxpREYsFJF9JCuyPle5KYYLiAeHhVntDoiTxrR
LQ9pvKrVug85veLkGmGfyaOVAEVdGJSTNgwlCm2U1HJJVRLBigYSbCW725BzWOkY1RluKScEDuwl
fQCXBoj7DreC9QTrUIEGOgYkv8jLY2vAX5UC4H0Bu8t7FUzxQxVs4r+Vw9Qnxj0uh3kSFDrtZHUK
pDJ9pfhVzYn5cHsz4vMk9uwKwSbyHR8FaglpgxtKl5BK42AiEZsoADz2Jd0+UrADqoenxTpnrTwE
Y/cMJdW82VV2qQzywDg/g3KIcn29DVUeNEyrVVEcn7EVODpzXgolDlnA0Yoa001jQtx1Msq39zSY
sQ2+Wmf44bSMcNQB2b9/l6E2H/pyXHx1wokaaiUXNoEhUXHksgv4T2L3BBhSc90KtRmNrHb46qGq
2K9+FU/iOZxlentZ0ijQOiUAb+ViHQYoNP/nx6+3iJclHceoUgSabWJuHpcU23dxmY3Sa+MruUfS
/XWlsFD1seQrJ+xexqjy5Xo27za1GhxvN3s+d1Jo0w8yPaRIJ4AW+LCIQilhvk200e/2QNqRR/7D
ETCSuyaKlQRfKfUGZ6fimzHEALv1BMYu2hl3gZOAtmEwhIOPPvDSLPga0DR5D4EV9sqtPxuAWqjc
sFhAL4WlNceVJVDoCEueUd2yBRlEV81s9zJtWWxEZpIH/8OTwLUNfaX+FvcRUr/eyOLszNVMOROv
FQQxA7euitTDsjghZeLIQ7YVJMq11RFlqFqnklBhwvBuGegK1pcUfrHj7UalZiXxGwbNWf4getlN
tZnyVvnf1Y2gmirdNpNYWu1SdI5AvOXIuz2sRlI7MztyJCHqQo8/0g3QEHTNiNM/9+ALjTOp84A0
Slyzak294INa8yClUPOAKWv0pgMgkRA6IRDTURKJ3GgMRZkEy+q+fg5CAsw+qQ+W45thB939fqkh
m9Cyn7HXY0v0wvqyZdzH8SAXRwL/5W6VgFxQAr4JLqQLtunAKSt7giy451KPKYZQnCkeYVY+ijYC
vGbWtPLUNvW58NDJ7l5RVHibkl1wAGBjIQ5Ms46KnTWwNvccdr6i7jth4vt5OMAkDp5v9e8Q6825
bP7A5pF2zL/RdZtnCMiwUCfTKyXpU7YCAZjyspkVfQ/nyFBOXl4+DMmQUECkOPwxqsfnrqRDJHfA
4iNdCSuxiKzjbdXNmSXOe3MH2NpFs3O3FUljJ68ROftP6IBLBJxsOVe6WzkMe2xAwZaUG4gBEvy7
QH8lyD6wF8/e+adtcX7w55ey8u+k9VQO3B2Ej4TSwcSEBQ2DKSGY2cTaE06f6SepbZWGBhY1jhlE
XA9w+u84Pm819I3XihJZgAhP1H85TYciapQmmwyxzVRs1iixGgEphDlgZfFXm48ERV4V1N/y/KTo
OzzRo0Sk

`protect end_protected
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.1"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa", key_block
T5QXILUACuu2UjL6QNhsDsHPwSO8IBDd5vD7SmlO2zY415BDaXPrb39mNXMTBLECKIjiam1QQ/eJ
VmcDsvb4KFUb9TOoywk0xAWyiU+H/sL18oPS2X8TziBe62W+yEKPzttA5IdwjYlPeRmQHVxUn1wu
iPsr9L3KRpwtiNJUiOL1JVlY2lvGe6yGWhEEQ3EakQGO2g8whqKK4UNjVjIKylEcWpvNlAPGfBk4
SIqr3S+uCHS26FQMHdIIFdLHvPEDZKhDvZBKDNXKm2nxs1gy104NmEJnWlXKM1BQ+D/lxZCIosof
Ip9Vv7uXAtirtPtcoRIqk3+drHbr0k2Ma1D4bg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control xilinx_schematic_visibility="false"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="qVYNmErgXmT1rj+EOC18AcExJqJb4K5PZDMPvVr90d0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 284512)
`protect data_block
01UWoqZ6fPM5rtkE/sH9oxGiW5On+4VZeKy0TXq7vTsDI60zDprKknObfk/EkZa8+JO9oY2I+XAv
j/6bLyJUt6wPlIVpwhUCqgrElf7rDHIa53VcOtzuo6PeSSPGfBYNK85xpX5CWsRFlOcPQx+0Sum2
El2mIdFQxGqWMsFbqriWi6YaDsKNqoR6DcnvGFcIvLa3bzx9crqgKTP8I/bx/rOBZ7nZ8Fq9Q7ra
oEpVpTFJDeuQ7bFTYInjdLmQOaRW5vnn6reYoz4mVbIKfdXUEX9W3vX2+CBj5Zh8zdemKLIl/1eZ
rtzkkQnl219RsDYFQ83XkcSqqWxqY4j9Yx8t/YGC/N/rMTurUxOcdUexk1220eHFXeVicVJ6kyvd
zFp6R6CKWOOmMmSi4+3J0cuv4cSwHqFB5i5pxP7RufHmuoXwWECEWymCpPxwB/vP1u0/0HMj9y8Q
+hB3tWWfbvlrAqCSY/QJH3880STTlkF4PQtLe07TjLgXTreavMwtvGmqTmAyh6AnIcjhKJDu5ElW
8/bewaeFI9ceRCf5cWLatNvY7oT7rVruhOy2hSOmHdc89PKjnM/oZjwboHJ2E1Vru0a9yU3m/GlY
TCHZpRSG8JVTbUaJbOD8DklmGx/I1WK2CH+buRDiN5fqe5ff5w/fJUGwKUF6/+ENP38vWkm8LPBb
JaSsdvQ9ytO3LFazgRQHTFlo2Wb8gjkn4hOB6YlZNcYfxPdOvtjI3h6WaSkDmwU6+hrKtySkHSVW
dnI3xhT42TqVoRtifemiTMCpAivV+br+UiXgvTmKGSfF87mnpxJt7N8jMd+uJHLTGYFEEx9tqTkI
LtkiSJMy2xoatBw3d+h0Im3COJ9P78OoRWdms/dVytKrhB0wL1lyDdzJHdWFjAAq2ZMLXQDSY2gE
Z8AisiPvWskTLQd+4d9gzhHiqvjIosSJuOVF9fYCp6UH49TiIdUJ7bxMRvbWfTpNWpjo5r7fi5YV
Q4R1x0sy2dzwycjUAUk0RPJJMWKGkwKMNup5bA96T6d1E1tpqUp/Nh9ATzwTmM2btnBtHETN5DXX
fVRFVKADxPVVfiv/iZM+t4X1SbCxgmzit91F3KJgRlNbVTpEyXY2PBsO1vE0r0kVh0Q30LbPoasC
Q6+8b5CeJfe4DHw9G8l02vvpc14u4v7SctWnh9FddBZSptmEKw5IYBHDq1JuTs973wy4G59LBUIx
qlgwdOzlVQsCRXa82QGg8aWwxb41fO5xem1AGqv7AIRYJ0cJsSFoVwMF8jMR4lrIzYOvNtPUdwyc
MtMNCJGwwvORLt1BN43bch55cayMu6IgeMjmZhUgHd9BXauPh5R4CPGNYaYITrf0bERktGMgFv/6
d+tmKNm4FIayx0Wi6R5IKyvIzu2zjg/tVpLJkiJKw7J5Q5nmJx6uBzlutYE9u8a2MesBfDTJdqEe
A1xN5FS62e1WdXSJ9BKUtDheqFcOoYeMsS9M6cSyvLQhcLTKBDlju3ZgF+FuLKMVUn0C7TQtfKIv
dH/FDGBQzH8bgENB5h3tkV75WIt2Ts3ySfUg07Kkl4DhPaqJhbeQi74aP5EXjQjYG60N5dzfKTyA
8x+oxf0MFEc7YYQzUph+7wvy/AsXbdJp315T7yzYq03qoLikdplZqsc42dEx49iP6BqhD7oyPSMa
J6+ZYOuwIO6eUcWkUiy8c9PVd6FeBQoVJFlvPVLpqUsiPD5GWVNRgAbuuRNkDwozUVpyrcQXLubd
pJuGI9COzTZTiYA3KpRPT5YMm/pdUsAJ6r7U+QoJyMod1x0g8/JG+fJjI9aoq/wyHxSoq6ATuNmV
hQzffUvlLmvvP3cLcXt/U+7gk2fvmQAx0ANtnXlfrdWuOvsFS/iV8wdUGE2BhC3YyPncGLDFJrjX
Vbtq+M8imiJswSER5W6EVuj6ZYgbkCyQ5QTLr6kj9OuPtIKsYOOQlY70pwkoEs5Icbqw9vYqiYi0
Vpf1sNY23g9g7yFbrBviDc4ocWum+4twMZgXqPwQN18POw72M3QQN4ixpShu8TtY1FDY6gLtpTo3
TvdnVZhAnMDHv89ZsrQ7KO2OgHSfmgAZrfWWDfErC/wEbXbnAsupELCLQ3ZMSnjtYtQL/1Z6cUjm
NSsVl2ADCYABjPCwtkqmwtnV3H8THBBLSlp513F8SsC7MgLps9uD4vUbwGPjma4DERw15qixc9BJ
ECvYw5hLsSU423HPpRH+JLSvWHkIVkxZ7N6DGqLvy7peXkXJ8Ads/hgWx/M85WVgcwNzXpR7wBaV
N+itGVVEkPfLcRJLKYd8pERV7UYRzQQWA3GsaiiEwgQ7570N6nVXPWDdmzU6TX7yiLNL+t9druaG
Xlrm6Duu2jTwQM5IwwvGfvYoNsmLktb+bgqfxUxfuY5PCVvtphc0OwyUbMwJ4hGjVGnTPTZJ2FWS
zN8HiGJ4FHMkEFGc003obeZYcgJJV3DC3F7qIv9PBZnjDEepY+BS4KhTzzF5yYmiegSYoS1GqhTq
I1rkNFwyMATmWQIS/0nkJRxZ3jfZCHRQ8e/7D0K+Swloang43eM6rz81xqdk6UDUnGP7r6DiL/yN
BFYqWbI/S9lmy5IQixgw7oI6jsl+ptFn7dcMWt2wBUbpqqqf2/X4e1+W+NZrBdX/0DVcgBSbOEJQ
I30ATN3kaFfvIhD0tVeojeYORHhITVsW1ZNtebORZkvnoMdlIDUJgOEr8tqVJvivP8LEgIzghYXM
FDopI+rtFNQW7fkrYGduFxmoFfwCvP3NxtVDIhm8jaaI2Ej/7RkQA1pvIk+Dsl+IOKiMBiKtaEwo
yDNTLBpTg52px0OGoTRUsJdCIpLOYefq7U1ghH+FAK7hX8cDztvlojZHheqMH2WzmyU9sRvgsebu
coOVQQLjo6xzpdMnFeDpphv7ThIeo3u2z5Y4pKbBPkcAkqbw6RObxJXMCYQGRnR5r+EyrSi6ZcbB
E/ostvh4rGrW4+hbVsTABOgaD07EAE6lC/y9u8zQ5klJn0jCwnZ0AOWaZVRV0E/DydkbhZUyK/QB
kZUaFkrZ5NZQ0CtAAgrnD7R52ZPcdM/428rvNXaIjRPsd0MIc7JzoVKVOqpiJOz2KYlPlvg+EQnj
enFOCJwpHutAAFD7Vy9iIpnp9LtIgtrdwgjNFNFgNMssfN4g+OGqJ5oP8Dkwi6PhqYuU5HSbSyjZ
GJnQ/2rrJbxfhL49mzv5X797g1wIqu6niVx+Jre+XJs+NtMuaqHhMe9/wym/QRHuKh6f7SLOEXHv
oZEoAARKCv/YS1l3rZTE0QZla4ewKzvniwf7+51E4fck2yeUYuzBKTA+M4qmR4Q7sVGI2u6rMpvk
RWXxJTt9jxxTbtDoI09wBea8fJ7McYrVuAmt0R5LXGOgfCG3PzkZUaRKHw4XtTbAjHSjIPn706ik
PLNJ/IOInEtnO/zSGq2paEkha3v/qMCO/FWka84CTyXJDlt9nh0SgGb68qjvSDHTWN7qQcuDD/s3
MKHuFw81qtS3ZBwwobWE2dTUzFb71UhUHMWhs9+Pe+nsxN6VKvVmqTEga+pi/JKmK+RI4OyDUCSs
vDaNiHhiiKH18KFD4VJ2uAMOP6rr2s8VzetCssaHT43UzSHNZJs4ptdXeEynexvf9eKIhzuLCJSV
rTebQlWmuoZFqVGOglnr5yHLOuVWHeo0I2erzWPMkGvpbaZ70kq2b4vFBbSm7EbdWVkZ4PQoE6NC
N4eICjrmq0AJYqLux8dGUL2a1MPGfbJ+Rv96WXCocT3qx55nIewPxy7LLgtEFYNMbyJEQ18mrRqo
mTkiGuXJLfXy13KzTlZrTo8aNJCDVFiimG1is9UtDSBjwwhOFDmM7PkEtH+bsXqJvzbwCoux0Ym8
g14oif72Sm9RFsJxKhm5YjABtTtg9giIt1C6Omjlwjy3EC69CNf1X22QXsRxEOpNnRirQzLPBARA
sFzCnJkUu3Wkzxc8Tg418FRhzSOXvs840agvmJV1IthY9skBYKJN+4ifiZko0c+cDzeIEsRRDsg4
Gc52htu7lxv5UeJZDPX+ConYW34YuhuGtvGan+PMovDsqE6L2GbaOaJUJm728Fuq5r4NPayNryj7
24KGd2/RhTQ1ewXoW9oNDDBks85VCM0Q580RqKB6Tq+QcEXBAMNeTXVWSR1M3OakMEcotNxTxrhh
5YM4Nqh054lBRrqS3ljRp9fml8ypckUYKpfxqC/Oimn4f9FDZGo3BaQ0xuww4KLYiqM5P0tV1aZz
3Lklc2LZ7LPa/rD7hQtHveNqi03cKp51NUKVcEP0A0Ko/LGhhI7WVpMU98CWX6m3oBsbvdOh12Yj
LtCzMlDKRBuU4DKxxt0erNwH1h24CdR2ObOTtzP+b4alUXEOn6Y+fQKrXPXekbVTCQfa6zP0KTZw
TZ3dTmIxeeJVstw9XqGMPMAjZnhHsJPSBauXvgoVV4NkTTwjOJRTD8MjL/15MeH3/XRXI7jCFHpe
h/Ddk6JnIbdFH0S6FPI4TruCT+yDpBy3EkeUbTBx/k4UXw3I7ouhxwCFdjFn57VoqbGncCWOPCIu
he+hUe5wNQieCEj1LG0Uv4DKM2ey1hE3quPe77M+xmosfHPOVTpfybLnXFddITU2pfVFdftPZQiz
j23yGS1JbsySfPHaXHjd9uVSj8r4VwZWuIZYbJl99qCk/N4TR9Dt/yPyUh6NImT4QKG79nE84ex0
J6FRTJ93Qr2hF1x1dUDjRRvmLBAydGUcEc6s56TnM87TMwZxw+4G+MbdvlyTK7lTBzrlMnCl768r
SIqj7geXGhL750jdZIU8SkmtR9w7MQ6zO6X3bkMVMV0BcTEe2HBVM48WBZyJEiCT+YbDxAsXUmWA
IAAjFAjKkoRhYyUXVyD7zfRgiQMisNCnchcxBqj4QkgYkepTFxqe/G1LTdfQQR3XDiVjIiwsLWq6
g20S6J34DN2CUpBybbwvcJTN9JFSCsmfgp5C1/cwwz4wqCvOp3JXSBbec2tjS40TkyM9yjnRLL8Z
otfcyGQKfu1a2A6HnnaDHr95DuYgASHx19a4xNQ87wVE+HtWz7s3DASb9a/GrOMsDwdh92XS1jK/
fbvhoqU/vuvx+OpjbSCE0VaXnBQSAyRNZ2EMkL2Ffvr9bTX4rg0WcYjeSt8NF79PhARB3uJP4hZZ
qpxsT75Zjq8UCubzyVRX6VP9aHnPGWKxoBnKrZcs/egFfizyC4pIctK4f7CqBqZ6P5c9gOycZtyo
/rKkllFW2SpWXiB1pNqulOdWx3WzOC39FkThok62viIM9MW4f5ljO710s+d9QkM+XIsI5aotSpyw
+mjAE/gYWkTxXN0jhEHLpHrzecgAQ0itZJt9fTLFQJEfQ+3YOVZFVYTnMwrGA3xkjq5z10GOT9HC
mAQ3MZH5+VMpmD6KPAW6TnKeGLWcoLmvG0GaanpOBYpNGHz5JkhS7yJ1mo7aDHe9Fq8Nsv9BliA5
/s24Rdr6zle3szk4VbsdPuad0ZcSHg9Pf/LYEX2vifXcEyXZgu+lec8RAMfwGAoIpWhtJ5vrs/3F
gqlepO3/mH1uFSkQWFLOisZHV6NSqwOR6D2rp0zyFv9nB2/T/HO8yMaoxnxeIfQFrUd6aDwn/jkb
qScpX1UcASoCRhLRRbvW46lN49DYiDejhg/PDX88+PrQaSP5qgmCLOH+zeJxLIdkGEGZf846MlKy
DPihyw29VYAC3cgAQ5GCBBnLVUTbaIc4srYUZxSh9oNSSBo8DvpuInHtvafjLM81zN/gnjO1FS+C
QpIlLbz85OESb5BGBhH7PAfqinJKsmHV2jffUb9tYC2U78HU5i3g/9GAevQLMJkNtmORhawx3m6v
NcuK5g4BzR1iBL1gK+oKlPiEDIq1dp+lBsbC19Lf2n7QEIWhZswdasa7Ha7EHkYAp7mL9rIF3i0F
mjpKvmazP6rWT6MiFMx8MDvwYQaEpxxJfQX3MhbZiruajueb3gEVjfwleX9o5KY2CbK6pjHmQqvv
BKK9OINgEI6ewPRl0mT4moPWyBWlC7SCC72PftpVoh9yh041fpPyuQ+I482pe/p9l3pdDUQHIWsd
1qMJArB3CrIxDZTBALN8P3abhebJnvGPfr9vP9L976USfX68tpZWuEVOzpATJBR6FaqVINjMLIX4
xOVbuG0bDGffoUsDl7ZpiGna2u0u5o4RVUfF2SY7v0VmuoTRQZIiILNHgVn7Ur1VH6SNgA54+JxB
0uxMd2pAeLJsRiF52o7c85J1iYIPMgVufrQsU4O/Vx19j7ffr7KZsQW4sdX4y7iZxX1ROjbqLZXv
iWrZ1Hgd4MzZ1mMxjbOlfcpwgsmwPT0cw/UFZrJ2kjoGHeE5x/wfv87KnZO97DMx5wV7sj15+sHR
2rPh6F2VTMFzkFl4pmZVpZBUca9I4oWqWNflMP4OBgPky6K9VDnrc5NzycNhdK6iVzaZCanpMFKd
xyjPEM7edYEaaDxzwRp6Yk5j3f80HyNaoecCAfyo/Yti9P9T7vlgaLADgHoTGX9vBWRrXtZ1BvOR
7va2A0PL29uwUokmqs2ZhfiKjv+Nw9rgUtG/NOYwhPfgA9WN2AaG9HmAEa6nEOFcfyyKbDbQ4G5g
9bsUKdy0vA18L7Ww8vCYCbRwV+ClnAeDtgY9v1rFYpo+g2Za6f/FqLXycRQp4pUYD9WMKcSMUpZS
8b5M+Cd16VNCXblDNStLbmYjEyG/Z/r5Ubg/vLmlOg1XxvV4ID8IM2fhyLhi0XNBHXGHa1LufJ9f
n6n+7OTWkEEDee2cOqCkDSjKL+Rc2gF8Vh6JL6VUwoWPlGnTTCubRxSnQUEHGR/24djNUaruLzp3
pJTpwyKA++2RonpLNVyXHrUb/2Hte1OVWDALyYS9ngXTePB470NSQyhuIDuvjGBmpIleYfW+d439
IRt+fSsBrHo081tPF1M/8SJU0idXsF7yTiPhqJ14z+IfD/Nl8a+MgCqiVfc4He5DnjgGg3Ob8Mo3
F+MKBYeiFlQalBVeJr1dkC19oa6qViW6movuMLK54hxix/L43uIR5CnOnwTHlrsUl4eXPlSk9rxb
xoLMCmL0h4KgDtD0XGtIbPztBDlWEEAiHB/trBgFuwpiL/jKYyRYPPz5q9uL6GY4fkIUacT3GTif
iYeUgKPM0XyZ2yMHj9TrRg/hxeW0PQob6RVvJRpMpM3GLwBFhPtL3byK3eaz6IA412XX8Eae0TSJ
rkv+MLxVkYweUEmD2DFAwQ/2vis0zBjhOzDMT3POnRh9/evxaRHAxgBw8n/pAqUyPH8Zq0jZO2Ec
f2ZS9XAcT5h6y2rK2gHknWaS2pCsFtgPOhLjzcKJGoYWdmwHFrezmQn5WPsfnvB1uifEV83v45XA
ItumYutq6nOzY3xN1n6aGN5MEi7M0/27gZBU2ll+pRugUrJokbelrmBr8SRQj68UwxozmyPtkFlK
YsS3EEulnsI4hJYBzVOPwbtr0lKPdN43ii48hbW0fI2yBmgetMEETtSv4U9X7unYwWf7RpCGbgU9
wcI1bUBhKewnWqXMbos2NKFY10UoGdlWDwNghMpH6wcUnateaYut9Ioce97MOI+WDeROOCU+Vcgf
ZrzpOrZrUAYgdomeqa37Nw6odgSqG3oGcvkh4ABi0KvQR8VKg6mDEW9kebYVARLo14Q8kUsqURuh
bvnBGrUfZCQFIb/FBK+z9Zt1NOsIsPMl1qnxGXS21r8/tIC6b4mFn0fdMjL9SZENJfI8juAQ+w1a
OxFLgoRCAZdPg6zVVdCDCATj5zynQLNnHrStLFVYMSlM3bN2V8KvyCKaDZo3Z2FC1M10lhnzQ2Eh
5/7c2jKvB4+U9EFZ6wiPiKVvx2CTs9aUJNafV/GRUxfZa1QM2k1viXlDvLVqz01L3KQERgsftSi0
BH9I+OLUfCmHmt+pFN4wi5m/nulc9HfVpnRPwdDJB38DFLijdX4+lLv6RB3YNCcAR/B+zozJVog7
CYnidtpGaknJwdhV7GuDAGHoqxEm4bBkjAcveZ6vwvDC3stpMQNzZC2ZzL4sUdZ19sZuvKOAlJ2R
rVnCedSZ2RqzQ3EC8y7YTP7j/TTTnl/firfRi+hsSVztSoSfQC9Bd0TBTgc1LEq4j6Oba4IoWQTj
dYIz7XETogVal4Oi2rv3/r2AcR00Mb+3I3F/s43EQ/DtiTwaGey9vX9dS3Gi7+wuns3U4gHIkOYP
ibKFjdKAgroWHGfsRNxeaJoUEV3dwz6d+DUMG0TSsrN4oBHNSYDmDQxRmIBhkAGPcxZffXCf13Jp
4FCW0/rrvCZRiEd3rdPGeJRziiE8GcdEeDQF5KqJmih8rOm4k7N9n93GfarWjyNwoEFUpkiqc9Yt
yNIZ9sZLDwhLF20U1PgHxiwSxzCNtXI6CiFivsrPQen9HhRjWwi0kQt+otiAFDPaHSnuT8hXsfKs
TLWAmeB86qRqABOYxZWSIIjUgO0x1RjFNY2Ek4G7O42huoR1OUA+ytC5l0pBMmsbJ/do5EMcnp/m
U1BKM0wAZQ2v3rbJnyNK0CTB8vI7AAiNY7oOaF6GUfqrhwLr7LdZX8TP0VH6vViX68B3Zxakdsic
IaTvYXz/1u6Tm148Oa7oLRLxPzxCBzKvPEYLMdpFjRGdJQRD0Jh9ipdRnhmhERCgKaM+mjwwqr4b
sS5kjOHemT5ZwUgCVVE5p+zwEWAcFWcrtUYpmuT7nJ+Bec7mMypqivePkUpW1wRay1Y5VAJC5AXC
UcAEgqQ0HqVYTh4axOOZA5Dkp1c1Nze1wobqXgXDf7WmmsP9WVkctVTeIOGDNWzYMMbnmxbYct3w
hPhcYQso6AMMpWU9WkkyVFd03JNjzlXe+t6iDuY5X1clJSRvCsUXh5QluwfrO/C6DD+UJ5JV+j20
PCYckWURTnWS+h0gezftTU8JVPdEgnryoICS0rk8CiYFKLypqCY5EEU3NyIVywcDbuaTf2tEftcC
QAwuwUE0ousRSoBTNJhsOS4c1Jv5C3oDaemqawexnMWvCpB7XFjAHqFIy461QIYVydjda/ckocQZ
LzEYN7yGbP4gXD4U1U3SXEx7ir0hHzlhOiwu5DZhXqcYX4rqeVkVymaF0s81L0rVEHkga5RW2Sca
bHoje+9z5CT9JTVq4Qqno8Yb3o0QDtyr1cIwXFgE8Ux0mRLJ/VwRFWwfOBbKkM9qRXdSOcz7quvt
B/h7CAPuKt55GoEcAHEwjsyCTrVYOoW2nHsm3oNc0PWlHgndPkCj6xKGVkt1b+IFCK3wJTJtWEa+
JvgJkPy3K27qI3oam5F5I5QcgzbolF/CuikRzXEq+Uf32Ca/9t6jfnJgUVlH5/erzq3/9ItyRz/6
O7FdsnX0UZQLmmS7/bRg1nijYi2M2FbdXoYXwrkF8a+w6zNGX+JhyrAS0qborIgGcr1t/yDc48XJ
4d0iUkiTD5rZHaHi2lUA6y0/sUGVabZdyAWcqjY+YheILIYaNPz8hDhNSrFg9vBqLotZThgIuobq
56kL+z8mQMbW4yhR7Hemah5Y1NLQcycMV4GQMRsF262HhrxPNVyaTMX6ykMq1AQCzyhnuRCijAYI
r/uy9qUr+iCS7AHtwpM+u/B5+fFSYFD20VcySyn2+39Md7cMemk/fR9ci5FjCrXNkMbJhA+z5Y6H
yPB6Vho9Cc6UDu12vyHWBpjwd9Y6slqgIXzyNalYKA16vT5OtRnz/VKq21WHe0ph/amw8c6TdbFu
lF2s+HfqP4McfoHlh05o7mBQ3vy3so0ClchEEcd9BB9iZbIvBd39Q2f44rfqL7zv/cpocaaLukf6
ZmbOENI/NxQxAQpi6YKTlyZngrYrfFBeTgmTXzXbhbB/OsqSe7oN8hfL2DCNXHI+1bIGzopa7sly
DHc5yQVpto2nbirhzHbleH9D4ZgTI/nF1QkOXB/Rq5nz3VbzVIRVy3HRnkXpjc0uGnpbFAjQjNWn
Dm7hDaAR5k4LCQRxJ7U2ZisT4g9M6crtsHGDBFKPxA7nFYYo8mHErYaF2YXjsKtJhY1roGrglnTZ
KytLlEjnMyJBt9w4ji0uaIq5IZc80/YCjgRmRRv8gS3Hfxvax1Grlu35B+HgGjVj456fqBsoRDjr
HH+O+lQudYQ0hK/XV1wSQvry5DAA2yYY7pPf326iuNXIEe7OSIZtcoIEHJog9HaP7kl27CI42cEk
0Xmv49BRYWA5VBIUK/rFqGncjVNxBOFwkO+ng7qOrzehdX5ZzRVh96rCSTt0qoiAc/p3oEZhicFO
lBdqcW/1Rpq5u3LLMoNi2zP2H1e/THggsRP9X6yGP3IZTNYATh1Jd1JxpPA0kTDrjxRdwl+RWtQU
hV2A7H58zCutOgmMel3wRXavyFF8IwG4ydvm7EsDwzj4l/N/XfFI9GPcsIj0LAf91T7ns3niLkvj
UBttpoQdlRv8dlR6ZygSsJNh2oZXetB/cMLXU+VCdbSs77h+2e4nEgybkpgcW2WWIt+eZqG57ObV
f/vV1Yz4x59S3Cu9fX67jMnDkHgIZ9VpFYUmMxMD6wcmEq3C7NzObe0DNOQMj/aWWuYSMz9xs7A9
gY7c3i9hhifTDy3dknBizw8rMhKG0VYrXBdYh4gi7djrhbHeR+W6n4BVo/107KScfaxl5RZOQQ6e
1mVzXUzZSt/oD2ZpeNagvW41KMqO1jL8bucvPu3TTd5R3p7Whh8LkTrk6C7h7h+u3P4HEEw3xh1C
pHp7BEFf+zo3xao45v/99VP9q4NsRcky69NrtnYU9XlmxmWcNpfcviZDNgWRJxjmonIOWr+J5ytK
uf6Dm8AGwjtujIeB93ZwUcn0zJBhnKPwgZymUNBjhENlNRV5IX3m3swUkkT8sBTxEz3HVG0CQw6F
txn6i+sTwIeOdsCLvV4wo8l8Tg+psKNRdED9GOZYygIkYhzAqCdts3R8qLrBZ+7SIAN7knZE9YQ8
mhnwgbz86MNFGe6WIszBXzEbSWJ+FA/7f3yUfqLpyFcxfFgOLma8lHPGqm6/MzsY0xy3q1MLrCRU
peCoRdSiqeJCcHkQNEzMCPlIzH5YRp+vA4x0iYmeMdwqmVBQbDRwdcdJg/J01WJvTsqbnvE8V9hv
B5ZALRblf8kO1OTw7svpuxTp5ihvWQX5Pc2mqhYSAEO3OoTMlCktVndrjElMRUYWTIS5HAPw4PFT
fAmY8wJZX72WkFCFIx7ea99nSkxbZjT2qcpXhS/AOPTyI5rZ9iVyzzwiUeh/eEhgNvQtdMpFiHNI
BYIGC7YIHrBgYJHCQ7jAfmBNlig0mtHPmHzuqQzXqtvchVgXbuWnGZAKZ34D8IwqciDycU7rQLEy
fuidTJErhOdFrBIcxesYu3Tq2it3oBqKRiA1OzdfD9XftZkwgSdEQlWnoB4qsn0k2kJoKKaZ0XUP
fLEWH9t903KUjalAGsM76X1U8Bic81i08003vxjQ/e+OIRdBvGiTExiDgsQOAV3ZtQQsvSr/aPxx
X6ddVvut9eo60eAyZDtcSf2oSmWCRUSL7qJ6DRB1Qz9FqomlCQpzPe/901uuylx1ehLcyGDZdG5+
0e0wsh4L0prZsZSkfB4aW5dU0qkAetx1NPv8pPAU104Y0cciW6V6isP9gptgM6EQdhjiWmmDZZHJ
Ode0erOMHqMkKdUE1jkBQdxsYUy1OM+i8n1lDvQefJBedIhX4hH+GGKAMEvEDfJY9jaXLq5S5flf
pOq8eg1aNJs5uiYifbs00OYtAMtA/o5/AABDlhD//9cd3hdxNGkTb6Y6/JHgeQxCuw26i8CzXXrB
q5G2vQJHYAHpOuqtA+DVAqn86vjevkNdnE32ZbBogfqlIATbQ0zqjnYVNhuJJ0gQx0SFPyOf+d8H
X7yWEpqcqZrwTW9v0B9xYhgD5l6/xBQvXebViY/EfTW/GKVm10ZpA4DoTYzanWKew8owNrCQAHg9
0B80DUuzQnKejGNT9up+WuKVU8JuFfPH0815MD3dq0EbrmeoaAQWHVfO1p7yFR6Dk8KIGr4Id0AO
CWu8jFELiSbfEIQ1PUT6x7Hud2QXzp+Deu3bEDkxCzGURuL7z0TTcNk56Fed1jmZ1TxFU5/Uav7T
KEhZh246QUnjH5VgQl6jzyW5mMfBdKBKuGn1RWvE1V82hRFeDN/GxoGk9AFRu2b7Y4dPPdA9yMfz
KLeMUsFOWibmcNb1tL55m7jQfaRJeYdAawIO1iAJ/aMphrSf1Zhg0egU8DmqmwMllnCqmYUGv0vM
F9gVak3wrou/BuHk4oLXWsZptclbqjZMCF5rEDXu8CrEwjVp+GN6cPNF7rOcOvZQZE7suzyoIAE9
w+gxZMg0Zy/aS7FLC+XlbBK1j0nCwhzIzTtf7coYN24g5uyvj3PIbI+VAwNZxmSwmE2NzHNQRs8L
r1ag7NAShUYdZarWRIxQR1IJYF8Yu4Lzu5WUYQGj6JRUF0+0mRTPvIc/YsYxDFaA1JAxtIt2Ps1i
cB7Zp1Y0CfiDh1YnTHetQBe55ydmNWrhTHirrat1BVW/kmRSgqzYwMjZrH8ZMqmnCwTlS3antbTU
rPXwPx7d+UJ5RiDjQUs8HwyMeCj0CnchI8IQhdlWCr7+BmufgPU27U0Xi/co/LTYOdiCBGjVfLHK
DUz0AD0bdTS/jXPjZDw3xJYpj7RfOZF40/vkczeHtfG9+g5rKCOktdjr4Ddv+wZVYiILZFPnO0dd
skVFLITYE7bRvQxnBfiCdLYpPVeOWYh71qThCdWtCqHSn2AHqMCIl0g3LDwsUFOxxdo0DyeM4dHn
o0h+QIuXrlk4ZC2+Mmdre7dYKsaeYNFjbMFPpKm8HETkFJ0rQhQv1AlYGyefRacYkSIAMsI3xd5o
sxtTHMfrVPGOulkNdDa6JMM91mSPYlCBUWu5KrFpjNZ7kyeyXRVrFLviSk9rmizJq2Q7hqAvhYfJ
Dgx3T+2ewcdIj9VJQM7Io51Ddm2od9b37vyHBdpJEmvJv2oc5xJmE0kS2PO6sEFcsTQRcZfIz4AU
eftbeYqLl5RsBkmo/7LyYDSSKxdhdgQvgdopEXH9TTLURxcXZ/wZ83Eep+Czy2+9wUCjM7s96nhw
Ismtxj4VWsNyoOmRVw1+wW/SavgX6yYP+d9zoGJZc7SKR/Ifvd7cSj8cApyjDWW9HdK7FysMVIC8
EnmDT6VmFBhHEeOef/PH7Ys3TNQmeJQL4Kw06MAsj3ZvPsA5YWpSl3KPotlFMqiaHihYR9oDp1oL
Q0SlZkE7usneFHEKvVICca/rNmdJnlqqqOHFwa0cXyGGvIiXzt76G9UjIV/hJHg1nFdeuKkkfxrP
C/BfxndFa+48jisbUB4ttnW3k4R/cM8Y3xKabciem968kibNhZeRwJnJEFUC+llTCY9P+M2CyL7s
L8lqEogHXTox/yrxrGcYVL/yfNIWXN9rL1af7L1hUrm+La/TXh3SDTBl0xEE8KCGu4M3jlP2C9UF
j8FDOrjT4GeHfYmpQIWGf2Rfwc1TwDCu8VnCNHPA5Wf82LvSROHtVELwNIfxOPkUawYsUKpfgeP6
DVwF8Psn6JZfsJ3juAu4cAveIuhoYNEO/mUha40pdm7gbvyb8BzTAtPlyzQp6qev36lwvYKKEuWS
Mvv0Ud6LF6jY+PQmdroF4yL212hyKaE6QGDoqmMVpb8c8iF0F2KjtyLw1RHzhTrKncgaRHin4Kac
B5ubKCf54op8FMvLKMAGDoRrUJxqT7m4ilIvalg8QPNbXHQIFv4Q0lxqyogEDam0e0C0d5fCNkbR
MCK938HorkUo1Xr6IEgSXAFEY4e6Ne17AY+g4JsMNZIacHqQa8LV5UdkZbOjDR2HToCvptMbCwck
xy2cQuY3qJ8ypLi4x+PVUBHG/QV1SDJvWrkblIqIq6hO57Xs6WUuPELMtkdDKCeaI56G0gu2xsdU
Gyn/gWHtrGOGMtezXsPqR0hMis9Op7cpYYcTzwnsDNHJp5cd3Z5/l3LCiMcphMNQlMhtGOQP+Na3
qQTCzNPOxmp5GFsoTAxqP9g1yMcTODFZ8Q8+OKgNpnssjH+4TVzrlr/CAd+YqVpasK/C6FCqHBuY
zMVGTdexcT+w6YbB+rgR2AEG8ZcVl2m2tGFJdyeYnQSMvp41hKqQ9KfZ1PhaxMKin0Itmke0Sv1B
L2r3NhRfYzjvxDrf6IgU23YVycKV4tDfURMK3au7GUie+73CVRYHMWwXfhKotorbFh2HKwtIxaKU
6ZV+n4VaLPU8opYaTCz6/ZMhcp+Lvvg6yUgIkdVfyf2kot/ws3QoPSK/0QKJjyzoIMMG/hbL/Mra
xWa7UH23XhZbwUJi/GTPD4OyAvHUnlcD3k3V/Q7MX1p/xGwyOpIX7RCrGC+XaB2Nvre78swe/AF3
dTCZ4v1jZVslfhiGT0sQjaVPn16QBLumvmwbtopWDw05jDV5zf0nR9fD9NFaMsXCiNn8EDPKTQpA
e6lhpRH9OXuwSEQF24sAYnU7NYNLN0ae9kwcA6xIC1/UWfBKiRHQc+2j2Pj1UPx9vPCjf1RDExh4
uMvaNZ1u0uflex+nbJQv/OyjGUIKotCVoH1zQO5N0h/bTsM3yym8gq6uH8Jp3QVHh62Se/c4K/lo
s7KN3PtgTBkzvXlxCNQmebBukKpyLHjy637nropODsM/zE5Md6fmD3HOyPjuvWtXWAAfiOl6XeOn
OhekFjfAqLdEv19dXDj5lAf9leJUWzSmQu/5v9Dd/gVTwiKxoyc8/MvXpOerGbAyRe0WvcYi+Iap
EwPaVevljHs/SnHUI3O+y38kHmFbB57we9F6ipYs7Q+XeBRYg2tP23PWKvsGO+pq1AnadAAuo1dX
oOkFFhzfIyQgjzanV6Im8ktA8u8cHUGkzhhR7QMlOev7npFuGNzlsQWLq05fAaRy1RSap/ngUT6W
cj+aOEmg8+s2blF4mh07Jw6WRwj5lrEY01qhCQ6x+iKfrkBamBjtf4dqX3tw/8Wbvbh0eyzVTUUr
LjrqZPQxxC8NWgvV8OMc1MPSI2mq18MbDL8cc9OHzl0qaAhbzURXFC7mHNE4ketdProLqiGZCEZh
5cTlLqkXEDSESiBrWdEm7gsG8A1Us57zXkm6qbjTb2hZKhOgevOSgDj6RuVX9yezoJ8OugxEdTtk
zBSMHptxMy2LXQothsUYfFCkv93XX6stywxm+bCJqBD7xVJGzQsZPWBhMOoVzt92185PDag/od+I
5kPV2llSqVG9/dSmQfobY618P+Z6BIdd0Jp4k0E4mamoBHvTCPrWkkusSkeyu4QzyTUSMzOvzP40
BGx2ik54m7o6LHN7Bebue93j4vFcTnxuVpJX4siWwgh/O/7cbndEa0AhTPSotf4LaFijLTueYRUA
qEAxQzYslidO+lTD2PkTwMwTtkqjJQRjvtP9VlGhhtrro76Kfkz34fbo0/GDp1F4hhP8wtOyRjgR
JsS2dYnyEPl4ZF60S9G3waRpwXo4P0XEa95x0XqW46kqv0LgQmZWfvgiyT2wIyS2OEuWg4B4CzxN
kfE6GNQhat0WMPhiCDk24JjuONGivRVZ4sM/tnMJjZ1MfhdqrE6HH1WeA7q8LEKaJ3iyE6tUG6l3
V9OBp0h6qd9xiZ3iHT6hw9UYGnueZr5aIR3HdZP1GowpjwTJyIm1r1K4Bb2gMnKj741NHSGapdnz
HJlZS7UXLj1K79eRZdP2iF9TVJ8hukxgMxs+V0jxz2G5PoxJYnhFndiVC/Mxv3k37DsHlGFC+Txx
5ebfflevR3UQB7VhPf+A9THXVpiUo8W3WUNtdxlyNPJH5OAOm5+ef8DmR2TzV4fK2gngAybvC/I1
MKE3yvBOTd3av6DeimSa/RbzYYIJfdqDzjxnamySDD5ITSCBSJ9UOemtandcZ11VyToctQQLGej4
HA6Kr7sxt15SBVV+WPk56H2qrj8B/XtFpQJSairKhOScx60eThi4uoSr63VbwuRAjc4rXivO0k9C
i6QePwh22vPS4c2BFP9niHfrotXLjE3v5Hqox34P1+w/TJ/Vxv2bg1h8mWXqTkcJ4bHNpa9viZ6N
gH24O2n7ksAy+0I8BO4S883jTDrdpZwBmTLoEZSEA+YkGpSzXTVC9awhQpcqn8xMBQ4EFCNocH9R
v518j26v/64f2ivUv92AojmKXsRL4oCwCjDMNkNHyeMMgjb7Tm1cXL0SrrASdRwKXIYkoy7cTm7B
UClkpIyu4TLhhmbZGpNPX3i/8uRR8WkLIgQ6o1BcAIYDq0SWdyug8XnYlAyU+aFrZ12kOBNhPCug
dtxOCLzKER7oESZDo65I3ZBhuV4W3LpUuVHru5zMsKtuIPIfLdDZlWmF1GB0MCsEBw8cHwIbHfpD
tIYnBPKbU0u/7zORiv0WPpsnXlvR4Fp455qioRz9zx586c8yRhMtLtHLEqBoBZBz6pfGT7tVCSZr
ElwJ7xQEq0SFFfQnyJAodkrhUSNS/eoh03TT9AfIZcGyI5QVNjr6YOgC7TD+zH7OY/rSiaUrrd0U
DPrqawqsHitNgKa5HjTxG6GZ9I/Ljzx3yIKqRH5wU2uc63XCNr2jmsy3M8VV0gKycC1F6L0JboTW
cdnr6Trc2OPdhaU/4IyfdrYyT/YFJcmV5ifdhtosESriTqYF435yd7F+gkCn90H5CbGiqO2CqC6E
QNFNUQ7N3uhFjT55tLUvblcd1Ek8Q5gcnKzqjeCYWOJbrqDGnQnZcV9WSElYixe9CtGkb8WpzEhg
1o/bS+lD1f8RQ7ONJkrQ3L0uz1wX4rNnbsODfu/DaGYVVlVuAmjnoMI7HdpZi2FKdH1VkUm9JGzL
6I8mzbeAcfUF9kXNEKOfprHAICCGYG4bxKNi9AqX1d5bE9AQmQokoKiIVr7U1jWPDFsKL1MR+hGX
ouOozAvYzC1Pg2TmVhTTZndX6t5rUOvUcxhIeLnNHhibdrqCDgDHwbuMz8q6FW0FKgtQupT7aOv2
8RdxG4/kZODoZ5u6ykg5TN+kchDjjOZJPX2Y3irmtw/t5Nx10uLxbt5Ewg4zy2mHBiGfyR25QOhf
oFZVng2XdWHnTkPRJSxKX+tR5Di9PjJPjNK7d/mehCT1PQk0BBorfZSIDprI1OMd6fG9q58d6XWt
QSUfcE5S8Hi7VFBA3cElcSQsUu5uLC6g2p8cf7kXUXfElTbDmfxlLV0QrP0BY37E9uUHg5Hug845
klGJCXT1OfCGs2EGn8Eyehmpja5Keom6VIa5NkO/SVQSgmuximnc79Fhmwbd38RxEwSG9nXklM2V
pe+7XJ64da+VV03GurwbFJ+gbP35c9VpJyoNkKJzABXI1opqc5750KVcKhplpkGFB5y3F5EHj5F9
+cdMb8aFwydsVctWFbvfbBV2aWzQqDfytcen8rVHXUaJYP5f8G0DuJogHlEEztXK9CJPbSf9i49i
svJ/XxvEBisJTeMp84T9ZqVwfpSHKGvZ/Z3Y0nE/T8HinvtqVqfCYjv2GBgWjv/9skYIAL1SqPbG
BT0EFM3b2CbMc7u9AySfexjeIGj/yYdcgKcaMHpge9go70LoR6VQAF1pD6/pQ2au8puoWBh15ITD
Lm86gzI9PvmQ6XBMB6QGNZd59t5pVx0phd7/2ev5Yea4rCfjPJYhD+dvJg0170OBxWYJlz5T1hio
hb2SJFvK+R1nM2O1hAhp5/9Ft9/durn/UvH/uBr+LwGFq9s1ueXmnGRMC25/lTXiTDqqFTiIPYei
kPLNf3AFkdm2G1SnTbZlsH7SF/CQy75JIsOBFhn0ek6NSRxTy1+tBTVvAp5ry49mtv0AcJvwtTsu
8Q2BlUTlP32PAo98edU+cAWfg8pjXfDsyZJk0MsjTTPF+5iYtUcU4iU9vjJBYDlsS1JzQb4D67CN
uSxLp2Mb58uWghDUJeUc6pKFHK51OMugLywvH2zDcZnp74GUsFfh2BKA42/jXajz1cRpSs95IX8v
TlNEw8hCrrdF3MXglH87nTxrclqViqi2NjMJl7VdZcQGtkVMnfd70dKaaCA5DFuaf+7TI5hkK22/
srY4Q6wLKdaw2J2p7iEJjz6K3haUDngQmts3Sn0FYhCDizUncvj01FoWNG3Ff0HjWrbHU/0liscj
H/jfIgCV6txUwS5wKLqZOGGBXQKqsnjdwYKem4knGTtz2jb6YjkWGabZWXySCPeGAudE24R3moiI
MT9/gE9kflujfAQwfSrtSPPAaRJBPxhudPsVDsLreUi3DBzpQrYPIWAK4tpKTRbxfJifZqEF+vZn
x/SKDCRNMlazTKbYjpwolnRuqhE3PL+ixl+Ej2304Lz49CfTNKVzG1LZ5P5Osy68vzKbIKmktGfp
MaOAt7KNCi7PG2w3FQzjxqqNY5q4ztbXSB98iXo4mshKAmYWMi1tk9OBhFJwOmpq7jDBa0nFZjgA
ovDg44nCDkz3Jlyp8digGrtyoDKI8+gPCwOz+Huc3Cn4PijtWxMa9ubXNA3R1oTePeEJ+hvAsOXY
S3neSRasCdiPQt6zlkqkWOW/lQ/3Sop7CHXxX8A/oE+qydvVIXytmPTvdOEqlMCPfaMEHD46pHZC
KzzTMz4BP6Nnkbk1XGqaPlUzxqE8Xflpj1/lczh5nbUMc9QwUqcy2dJaBMkeYvk1j4SlcIxFqb6o
ms/XJfLVTYXA4yfoo1lEjJizFYbCfmN1WHNx78hrjhS2Lh2S5LjWCuQklBnZ/CrjAyljB8khmjl3
c4mn/QXaDr1LrUhzTA9pg58VO8H6q4foYiYzD8Fx2KYGUSlZLwxUl2WfKfrlnuDzr2ZxCYgI9KWB
59853MaJkGw9Zq61GnsEWGg7n42gQt8U+xI5EDoRMSyGvmrvRwF9jXNgGhLFj7Im656Vd1GHuWQU
yRmh7zISzWZceAuMWgRa7Imz+8uqI3tPN1hUo1C5yG9jGjLGo5Dsfg6helC/3EmCkXF3roAWAWqY
L61hd1skGdfHnqgo14cf+14QLGZnTNoUSZbswCHNDjy0fTY1Vu1IDqCjPH+j5PztL0n9gUXcQc8U
/weqFZNm/22iwLKqzraMRsutRM6fw0hN+aSsKR4ScbtL2Vh+cE7EOhGzVD3vBF2B85nEAjfuy3rz
6ses4kf68OQs7fTgS3qmjPa67MVV1hxaLv+Bs5tm2K70o/s5JjA2UZaSgOh+rqM/UJ1w5lgC3mio
MGTT+GrsHk/GOL6IRBBFH+Sxz2mtUD2eltr/WwbshOHZ6E49R66wu4foLCE5kx60tB4nY5GKr4Zk
vry+EobZokowFwAIdMXoABPVEMJ2vtqCo40yl4U5AJK9ZFWRPL5UvcMH3DicUH0djtiyUqb9Y95P
T+bsyzLPnwNrqljYR+2xRzFjx5qjDew7G666ZzeExlij1hnva7dka+x3CHBrjfRITqjqy3pqxvx8
VY9PFHaS8AXZMWqELXH8k+nq6O7MnTIMV02uz3fXV0fBdCtrvwcf5UjEx9IBlNhm40S6lM7dO8H2
DK/IdH2oj5+4vaDEYcasUeqaH/XAuvkrT4nImrNo0p6UvHKnF2D5mPv9wmDkLfgb6nkmnHfsLA6r
evabgpyXxJ9s58QXVDX77Fwn0usc5yRIbd5yGfGDo9NHq95SQgDT1Xu2UTLoempspyHQoniVNSwv
vFw/9c9j1v6preG6mo2aKSPI7JuLqOjspMxKKuCngCB+nHfFzqR4d4Sto5N5XyPhN0WzFfysYbPS
bHQk5AFzsnSVnEyY/KDnKBJDII9xavIUm0dtao1HWQJ2Pn7dIeH09Os0eBW41OixuEm43L+poZRe
Mvdsy6fFQjxAxSgDsow35M3X8jxIDXOwaRTRv8W98OMJgXXiZPfhzVNkxPe5SYnU6oG9z0Ik4liJ
uYXbfmAl+pQbKC4NKC9hkXDXLmHLbnf51o9qh+FHONHJFsF1ucShaf/Xr48XMvf3B300c3avccO5
S+m9cWYzL09Y2s3pGhIHdWFU+pIXLfsrhLncAaeEmEz8ag7t2Ju/GN7EE1DOVN40Mca5iXBxK1+r
CqTaM84gN1n6M7/E6ALw9Z0SsBJI8s85sQV65aYbVnpr/vb43HK/WISdYwE1ilCnj6TNqitSudFC
ielZiB1nR6rOWAy5ZK/na2Oby9yVMU7jsgNoNJvmcNiM+ocB1Jsv1kcK8QUwjwI7sL40r8xENHDs
JKRy4wXvfX/cpf23xVBwBVGpv5MhSEQ2aVZh2qcNCO5yUdJnXyHFJzvO5FVTfI/hX3lzD0gno2IQ
Ak12ni8/MM1dEh9Y80pUdR7QObkJWVih91spP9xzgt4mV76tmq/J5TEWgsIdzCQbM5LD+BjU5J5r
rNTNoa+ym/Y7CSgTgzAyon6LKGV2CueO4U61sPpSS2uoJPQf2cgNh3nddd8Z5797IfgxQZrKLgIe
UPU+GV9UKUFjDge5nsCy8R/s7xASJxfOo1k4lYzM3JPysETqYRihfvqSDZkb94lih1lxLjS5a3Jy
LCYhoSd5frHEEmmOr5SkmmTC8T22uWvttHktRTAkfOCQ/zZeygg5ndrQT8DTWqn6JdE7fVCyS2Rz
dO+FLHOSe7LFvzAxezGV9T0VI0PH8iPsziprlChXndlDwsftoiJdOSu64pomVH5hTmO0O7k6fRLI
J3Q/BNl6Vz4UIF0v9XGGW9zp171uHuFsULmq2hXeJFUZIRbz+4mRmrrRDAXj0S+lO/JkbYftJk6E
zlGRLDGInFRdNHOIDoiINVImrq///oCUIn4p7BesjKfT+huLCoy5EN7EJUoqZhSuEY5/BYi+uzW2
2ZzvgMNvoMaXIwwg7UDoI067/MQ+7XKAj1joGmnZUH4RHdVpQbNPArwXDs7ARr2Kp4v/pdx4m/X9
YBySfovnI3F4VM5I4XZdYyJrZU0rLWooAk/zpziEJu6Qs8ELr3/acMguJUv63z0lcsEhAOjidf3n
+wmd3eX4ieNK73vqcaGe9enhzPE/VMWKKX8kxpdyo3UoJN6H9Mam4mzDq75FN0DmnRO9UaNVU8s0
+0iAVjt2/3oR2j+L4FG/iArJjGY4hxpEEPBbHttT0x7lM8X4WzaCeQ4pEJF24HuMrFcaPMHxSlLf
+IIfMsXsncd9XupSiZNDKd2MfTcBwFCZTTjV6GZmrrl6cIolFbBFc0eB57qdf8RTOhvY4SZf5hu7
iVbw3y2PZQE6LxFw0kfQ57blnRqi5ZXmu1/iab3RzFU6hAHlyL00TihrkDaERMdhHhw3EPtYnZgX
FvCHedmYOhJDQxi+V7HMxsdcwbDqK3tKmoTZQo8E1iIsRAs7QJ/G0ymVGzjo3WAtTvu5vVBjl+0t
YPcoPOuJMLD56/OaokiHsc3aOM0Mr8yngkdCVic/P8MleqE6Pbfk65k+6iZYIFvhgoizglBygAm9
0C4oW+/BUjAjQPjy64a+eXiDeOq6RBX+Ek2LLX+Ernp4WYH4fIsuHntuOSaKUM09B3VFnonWyPlv
cZ3XRVHz2cwwzqaofWnB/RBfa2S20CmfpLVzz/9UqsL5PdiO+gpRqaO07s+VtfeikPId1wC6b9T3
QPE13GIWPr0VYkmUzf3OQhL6+MfDFNQngKkk4WNNTlogsGMdYrjNMKOpmzHOhJVClMb9JPBZDuxV
m67uTRsLtCTPufaaW0WUzvBucTiGNOU5NRgjjQDb0n9bwF1og0pe7uecyCngnC8tj/yUBfPCIBds
ZDUI6OebrCEOo+ti4DN6+E7g6HtdRTbDlW8p4mecdLSYXNFoQppfh+kHqcWrtpULf2asKyjhT4E7
n4TXG4p3bytoktwAiCkwt9Rr0zjl8g7CVYO6uhQjy2gRVBvA06voWNSm41CHlRkc4QJU8wR8i7ou
M0YZNdfSnOsRsB6FIilPK3kuJjTylFFFG6BnOqsrWtjiWhVPs71AwctiypVlp8fT/ZsekT241vKL
MLrsRn5Ik/SdvKoQfG9CrNWBxUKIeILxlFhIrq5IeWXw3UpBzEpHOHPUa6z7PsYyzIcNgZMo6pHd
DHnKrBRcUjdulxsIUDKjeKccc01NwE/l908swWPJYn2GAN9SlMA4q1V4WLjbLY4NItmXQfF5PS7a
oU92bP44wAiL8TGVXYha+wazzutValrCRR9WQkXdwFUBGgDx4YsNZ46UyYssxfddLyjW9vXCcA+W
Qid7QnDc7Xpi+O8Aqyvj5pHzojDMi+IivX6gVKA1R/MlbZoc7MHhOdb2IeXMV573chxC2SaM6W6O
ulFzZtnP63ssDO7xoKeNJQ5JirK7Sr+QdQyaHzuGdBiJRY5TMoL1KYtU4IFKAaBrYDtLEbysT1Hh
3dX2+yrtQziT4pGIdbTfLPbo3mIeB5PdVz/NE/DhuSOr6kXv54jKSYdGYQJd4m1tSCHmrTC+5eMV
iTGTjjHpZLRuv31Z8i+l8M1wydYWJrKBWNrg84neHBaDUoVJ0yM9reuLO3YuNCuERb8Wej1o4pAB
dEzgqLMu8eYdHjmhndrA5INZkluS2oaGgPJa7L68s846T96drBQLL/IOvUDQU/QKVqkCdy/IBb/T
XVGjz7lTbOC0nKeLPAO+GYntbzBEPIuaQO7wCAy/VZqbimbsi3B3A9IuLfWWEu8tKSROPjeCB2Iu
0f9c/wRAPAbA94hJh23JuWY9lfpZeQWPzMDv/W5EmbjOmS8WPaI4muFXDlxB+D4+6b5Fxd6dH6a1
Q0RNyE0NDzcIPi4p2R7N1e01xFDDMvWIlESUIHX7s82YTDWuSTfc/T3Xb44Z0cUIposezf7g7mU7
NgB9mT8Wx4NvoY8/WQrs2TQXjKnTD8wjM0MFDBQY3/jmj5U3y/JkfPAce2uXpHhvguo2TKao70yz
PMghs773T5zok+owAvpGuk0X1S1P38KIAtEUeU082CjukD3LIMSqbsXUytQqmbjN1vJqsMZk0qaI
4Gst7i0+iu4xXZ8lKeZGIfCPqEOUWWwSIGf5aJX2VrImskv++oMTvuSUkANOVeDjMZY0Dzin+Gey
Yn2Xvu8r+w095k/h2zeIyojGN9SyTbyG5YvBq7w3zBHhh0jEgKY7FZksLfMWdQl1mGlKSmgrA6By
FCSHcamMd/UaICRVHlMnPLscCVYlijnH8Uofey6QX60ViglJf2mWfYQnafJxkJfJAnG9U6HX/wZ4
MIRnJh19a2pgxkIQw0aQZ5e2ixrDHhHgnqUruPUQp8GJSbC7zIdphtj4GAHkAey63s8AmNqcGeTD
eAtk2eFCu1+/SbJ+1ftY18koZS57IcUjai1nJsnOKVhUlM3YMrE74a6MuLutDEDPNF/7cD0F8XyN
FUw6CiV6Jl1a9lh5v/Vq5RwmFDUlHDEOfcLTOcQ6gZQ5BZ2hjJeiqKGpLtQT5C8h7Z0K1V3p/S9l
bHXD+TB33wwbrIoWNDfCZcwrCUO6N122idrFmeMSo+WLYyuP6q9vY+Eb8yVBGPALDJEwgoKlqg9Q
fDnsvbWSA0xXjhgRh1MPZQmzGekt7bGntNQQPYgszQcE+YxhZFEByz539NCPkvalTPVoTlecl96v
fbiJwTuLjH+89TEj1f2o29lJciipFbYAj0r1fBzmwnRDuFISCvjL1v8Qzi1DAg9y+vo6dzk4IO0l
5x8lQkOsu2QEoo+k84EIx1y74No3DiJZfsX6hKU5em4CVEeaDeU0pkbgd46V6J1Qh74CyX/WN4P3
WwLoFbx7lL+CqMNnpHmXi/7b5HloaBFhjWnFG33d2Ql9YQo35oE+7QwbnJquFW9sPO+kTTnv/BZg
I6iWSuxHjruR8nGw+sm6B1986D3EGaQvQtXbkUErjFtbeaTgZ2shiW8E2o5mgXXgEW2rWqeFUOa1
OEju0letYCKYuyj2oUtj3O9HnRXf6OY+ds+a2WvlaGt7e/1u6V+WmcOKuhxVyHbct65poAXM8BsG
EU54I+uUmEfrwXcaJWlm6+pRYKw/Fyu7exllcv/UXj3ONqCes3UBoAcFi7nmdUB68R1CyQkpKYcN
E+RjAdpFXUMyLCGKNStgYFFT2gDJC2PC/NwpSahEe6+7T/WFB16K3DzMgeozVigJDgW6dSLai7N0
g+j8qjvqh3y3CBV9H6mJ3SOOzWmN6Vzq5eN3AwAbHZVNSERQHNMWy+tqNzYnhh0Vk2awqdXNBz0w
0NXaCDDv/TcKUGis7GYHoBIeHWsfUuCnsG7HQhDmUiLAgk2wC20evvO9JP1n0p/tFq93XMXRmCCF
Y04fk39ZFE9pGZhg7qHDrDNxhhycsGpFiFv8114CtHsGD8FfsjnCn1OjpUj8Qc087IaXrXNEM/Pp
1W1kOdqjWZdoSA4nx08RZeMkKxvt6DjrDs9eyh9QmOLAd/ck5SMrpZHVIkB1cGJqPLzVi5MTQTJr
NkA6xPso9+o6U8LeelX3W3TTFou7lVNXDpKDAy8mjfHTvceMt/hq5PkMkYBNXBx9K4v3c1vUlXsu
jCiD4OduDVE4pD2m+S1P6Enig6TT0Xa4YOsObfMos+Fole5fctY4IuYlBBrQlsrrZaW8NV8txvfs
+/IxYi2DOOAbKUuxWSgr0w4LMnOWiQ+QUmAtZadhcqNPwejVNul3DPlidd0byxJCI+xa6PaTBZQH
ca0DkTsalGfPs+xlf7xdiboAW5+qdWDErVAN9YP84c4CtUniKw2lpGVGMm6lhGpOhpcNSf/NS+o1
j4vnFMKbGc9HitL93bFNX3Rze7oO9RhNo4nawvpccxuso/0b++zcCLKocpA8Mjwze8tue83Jl8sz
vqwimRiglX55reAIUx9pu2R5KiATmpIbK6RVSjtD23QMxVMJ0yFp34YW4+yMkcdp3PzwbuygeRXY
G13GCagINjbjhG4zz6+MNXipezUSumsMmZffbto75+XG03k1daVAJLVnGCMNSOFkuZ3zyFeNNxN4
RTHkyrKkIeZFHCZwaLrD9tCTIqXJIX9BRLDj9Omap1GBGTftw2aI4boH3OORDVMLeHpDXgRUhh3G
WRv/pDaLmpjgBQOqfX0/rSLAFCUwStr1GUiPHcIpAejCLaBLRo5rBN2UN7eBH8drQ5DNmpM6Lgrr
1SpC3WqdgH4wMgEm91PQLQl3BDkUKZcGPgq99gMFDVNEYvmGGt8rnfo1DiRSnI/wBmRynP/1NQeE
ujNg/sNVjyUZ1bna2r+AP2Olk5b8eZC6xGQb8l1yIp8MYS2GThJHjmL+ymjWBkwp0T5DuDbISSPZ
+xc1xj+WteOo1Jl9IFVzXvQppm9pfbkk9Qh08orflMkbY4j2X/gDTLN5oTHSHPBXIevKd496ypuk
x2W4iIMInAkQWWtn3TMQcFxwGjZcyPZEcL5/Hw7wBI90zO96G8Lkers3qnSI2S52pdXlEoep96zE
2sPr9p7mNY0x5E04g99ihK8I03rsOlFWp7VF+Iz8klAEEohO8nse1XahzMRWr2RoPGcdJW/4X6iJ
jVAQUYr/bdZtsais+o6WY/WxeKp1IW3ZtHEWsYs1gWvFUroxROmVHwWiZvyrp43OpPRTXNsH33bA
2tK1pCX7w4VwTjWc+21cYJxNn7Tls5DmN4NaC8U7xFKTIKrj7ToZC81iQ7TmGuV603HAELtfpQ5W
8fK52n3GmE3BNaNWJdpbaA7kyh43Toxdl6RGGJd1lKSurw5YAL9toFbKFCnNPB5LVUome7BuqRbt
7qAQ9KqiaU/srdoGGNn4dJIDarEHzry5xwdGcrF6cCsZZ344rvfUnKxNQgzLQB9e9/VCjgK4WatF
STX5oybv5jN82iZZU4aJpjJHEL6uOt6N8QsVNNKQDGcGVDwlPVD1tu33D8BIaKoVi9hDktlKmxNP
zs7c2wsocLShL1DS0f26amnsDJSaXBXnmlgnxhnlC28o4lgoZWKASsrXpahXKrlSnpiqfBfE6pbp
osHwR1vgencMRttxk0hRk0JJDMWwWa9FffaW0/LexwV47Pp5yrh+0NXek2hNMSsoKaFGSuL5efL3
ijpJw8LccQ+/aHu6/QE8hpiYgqB3LeVARdUFDb+uDIjHe1B88hnNfoGbCAtdif5fX2YHCBya8xa5
tV8hS4lPmfblqMY/YarfUu2W/t65enS4l09bsB+HkZYBmvBGlHOpgx+yiiCg07hBG/vUu3GdzREG
8PtiqioJCAdJdHrtKxv/nPcnpCUwk7u1aKP0e3baNq39Lf7H9Yoa5DhoQkmMYBIo+nqeo7Gb4tz9
quPvjSJKubCDYxbx+ShiFMO49WF2WLDAhLJopMoEScUPi7rwX3G15b6NsHdkjgKl1ALxiMhVrTVD
gm6D0qFtJbmJqnDw+jnhCEZTVvJhEE+fhjbP7gVziwSS/6aO7CnxJscRa8/ENOolDMU5l8dfFP6/
KxlTs80NCT89l1waTT7/aiyr0dA034UEFVixhMRI2LQ2xDcpxLgHXXb6aViXKFypEJAxgMt41fQj
rRVA9d5ko6ynGKSNPMDUldDXNtrI89u9JAP0YowsfvlfDnHEVxDQX6sBf0KNPhUOX9eV52Hm0e/n
87a3VeRh4O8eYi1Sgv/6CjsnaBHMIYhTpGR9wgMhylLD0yvl9x7+9/vnfr5cefgx/+PISAv24TNb
/CZi6RbcTKNZ7ywu9Zti1QKzb4s6EEkhMARpblu71WsQxutQPsyXrVuxBBrH7fq1t99f+ho8+61z
PbM6j5xKkXXmnMU7h1KU/4mjtPuf+iPry2KAP5ogzMRKzok0Xb2JxR4pGaiO9UGjckbwVqeAKu5d
XImOC9uwJArB0oN+M2NtH1UGeuTffhSpWO2teNw78S8Zv2uow97/bRRZfGdOHJq4J44gV/NVFkY8
3uwjeIy0+R950+gIZJB5IiBhwK/LPSFUMm4OVgdxhtZcFfVoPI+nrttLsZgmB3bl6QB8fkr9HaD9
/dDlJ6YXW4Y1cV34or/63X5+cSpd2zNlQ0mJJ5hhST2IkaR36wA8W4e7ox9nMUcqmvMZ8zFgnUPM
LuYvaat4hpT+GMfmGxE2s47QADMYa09GKUV+FPlDDXjbeBbbWltYNzshJGnzbM8kR73xBTDPc4M7
ja3YgZy9lFRznJAPmzISOamS7qjF5OKkzO7UVEWjFSgv/V4ozFoxslNDR/aKCAp0DU2qy2UDWhEM
idy6OnIBFtRiW1ENdgsWT5v6fNwmaVhhIFLdcg2Q+onD3r+J72jmoWxiPkuzBgn+RraP0K4xAdAA
VKIsnYgTaDqZF4NH4YDSNVSb0mrpZYcywgD91tbC+OoRyq4BXjFUEODeAfL912VS+l/Xpg1gGbTo
v+2ddESNkiFbINKbTY8k6BOR5ldHwFO42y0MleXCABWK22nSoftLfeN0wXYf5v62r0OE+DiIeXhT
GEh8UepD6qywQjocy/VPBbnztD95icsV3Du+6wPaBnXNID5nzJOsmbrUZ+8OdJEYHP/TeDEMwcwu
DGdvZS9K46gdRN+Cg5HSGkgU76X5cH/VBoMKmU+8ga55iPn2GwPb3ZqyruRFQgSYSGObEZKztvgG
ZRyApSgjBZ/bWyl6fRLHzqMoLctKlYHUVvot3v7ca6sqniGgaW4/dDyuswcOjqbZmLNXCUNh9wk2
f/1iT0s6k4VchtyiHuf31sSN9M4bbRq95Mh4yvU2dU2iPsS0j4Yof4ikWy+jNLPvoKw+582zTBO8
eKLOH2MtV2NdueyL0pHgv7iHbc6IG/MNZ+2+nnuqKaIgx/gSIi1S+I2VKLrBrzbIQQUrLHS8H+Ok
8A+Z0jUxsCTJRVUuHfx3AG0VXgOlvqsnCrpAuV1lv6u4wFuz9ZIapXJZ7FWz7XLCYUZLckKQLldM
OMCn6NX6DIKAQLDcVYnjmDilWY0hUr9Wdzd0ByW/8UCLZXfNuS5D6Gw5kwts+oKsMnnYZM9z3M02
mYhBgbRJ8ogd7fLyYN59ZydXsW833dd0IrT0aV1vyIseqGSofHZeI1Bv7WV4km7wMLmuSV6u73NH
thIkmmnOzmRcCoCMwUWgx8Vwa3Pvk/TrFJ/Jmz++QiMW1pwGcICsqViTsavcYmdCcfEuFJZmyBRq
Ia6Y+Mr/O2uijVctfGrwK928ZE/WmKCkP56CTZlszohr7KtQKiBJVHkMzBkpJbO17915hKTZlkSk
2dJN6wL0DhXWWko7+0t+Yen0pyuKlpJLIjk2qNS3TFyXbe2+vTZb/Ud0dnFbQWlFr+owIMreFb3N
Sy7JK4cOoeZed6EVWth5vfUUPaxWU6EWSgVVR2L4NWImZKIEHNUTuWUtjQKMFRtylx7PVbfBNRrX
TW7gxNVBMc5SBEljHclPhLwJYFi5qvFSHyFe2H2kO8s9F4ADSIVwn359RoBGoZthq3xIqOJ7eCLS
bq3jT71oDzXZYcdfE0AFnIjLwwIW+xh00rZQd3MXkW7hYMrsAYJzYNiTYrrDnRRfWThBdyfdhYIh
H+KthuUoktySnNKuHfm2Ey6Fm4GP0f6kX9ccz+rKNqJV8EOggy0a6LKUrdB8S5RuIQ5ouq9OC17o
ypt+X65LP6Wqa6yldm/ic/7etFDPDPtH6DLeZPRwYAMJH9ADxfL6q8W+PeGwNAVFfbvcHNL5hYG9
q4ksC7efRixlZAdEZYkDP85llCIbVNhaINpB7es1sUe0n48rvJrecv76dvtHj7y8nsZNdccn1V23
e5dJcFZIuyHi6BcsO129sBWqe9yjPNFks9yGQGZOvRJivSACtei+T3Dl5vCXx5AiyHW4SYz/Le2Q
0DWNVPJwt4zfao2Mp8L9iJnXkylT+LvxE4oKDmfvfpQWY1m95JXnQTIqS6sWnOuK8R67D+qGaE0F
lPXSuprLvjCFKtrI62KsquQtwQuOTdGKzoYwA7DdhJZTsbS/+ldSrWR1+CeBtGIEBfH36Jfdso9s
7jILI1W0xrtznyRIw+4niRePz/QJbntaHBtx+kD+DaDRDbFYQQhO9sVOLUkUU9GAsHrJv83QMNIT
otqZj6MPHHsDFNXGW11wqr5lL46mWld1WSQHLkGV0u4gwHXEY+0SlV4uuqtJr1edeWCV0OSEqDe9
JLNWm3tlmvkpyxh5Tt/1PnYvPtb++v2niYfz2akoDgYFA4C5aKG4MzRYf7197tPIYNwfYhfrfRTs
ioLI2TlXbw6GENLcfAqf63hKeUZfJ6JX7uZL7F61G7Z+BqeetaIX7+sphY363MU8fwDvAgsdW3QF
nYp97ziecFGbrp8EDTARifrNWPqaviFvwAddc8K3USQnsjCla52UYvZv2skITZojz4A7d6BfNIKv
JjwStGRlD6VlAV0BCvdNyjTTKsoffe/fZTJJ2Mas3KKxDraNswi4puzReBuI4aByUE8aK6nPKbWb
Rv6zsAUn4Qn8RLnZ2pa1OhZ1gbl7tfREbfLLQRnpYUPPHMxCzRNhyIoCB8QCoMzqGHCZRm3UN2ZV
4dueb0zcx1aYXN3b1cqwlaNaCE1jykE+K7a/Q0RdkUjIi+ZGMLZk+LLsU2YA5dd6YHGACOTeN0v6
Lzv77s1nG11RqPh9sqCTfnvBNsQ2WSLpkVAUVOTw60FUwC9jocR2BHzfVylAmWBpj+uptsLyLv6E
y7C+i9uSvauNJCeM4KK67F80GfJFt2wEYw9hvlXcBUjrPLScuhW8l/54V5AmU7Dw+YkbNAT7B7iv
9mLdnFDrrbpGVishcQ4ENuJUiru2jfMl5UNX03SN5xopBKlrTzjzbsi0Jht6UNDU4q2ZeN7v48tX
6aowJldfiCiEbuKE3FRmZ3qJljhV/NSMKOUTgyYE2OyRqCzhk4Qhjp535V+8bVUVC//Mxdi5N0ru
0a86M5gNxVM2uhcZXPiSM3FycT1YcPibQqV5QfCSD77jcN3TzoC11S3041yfrqcQ6L30wTBHPqQt
WFpx1OREMbK3kNAnas2wbis49kStx4ISGWCbquv1jE3ZNgM8hFbn/CjQtwp70bRb6YGUTcgFgCmT
tuE0kAufV6mqTFTv414w1I+pooG9t4CavZVqvipJLaLyyaG19o/ljArm//2ajfX8Vs2NGRO1IMNV
jV81viO4lL6wsLM33iwijlam8obX1Jg6Uy7rZzWUycbhyDq6INBuRvh6lYqnmyLKKHRB1jUsquKY
jkaAmOYg3FKrlTs4BTNQMwHm7YU07/EJexU2r53tuqTrwSAOA4ZvyWmuRDTU2YzkNHC6CC4SxiXt
KamVt8wh9wHyd+7ERvmQYFGPiEDLKYcyhfWS2+ppqaOsWBUGo2QZ1lZFA3ZZS5ijMEvAXtIcj744
k/6i7OK/A8qt/KJD2Rp9G/nueTKj50gIUndGcMJ+To5hXekzy5V0c6D7ibXYIp5DKWQCjjfidt8y
tOVF9aCn3rPa5kv+d+vODhTsURmgxWwMpUd6zEyAMTur0GFdRm4Hs1IV4H1LtryNpUoLZ9MVh+0x
rUOrLdTnWEVDU5qc/E1rOzAmWnUAPeAEeM1ZS7P9Y/TPmMrpAIo42D25YF7WgVWb68u5uvWtAVvR
6Ple7I+K3RyO7wZuP7kv2WA0AzB1LvuvW03SFOicpGhQrpvwXO93RwsqHc9YiuK+O0oeNWLxfbrL
/ADuqdxi3ovBPKovWCQQSfKNeLdxesDwMQIOz3sfTKEpEX7yUys6X938IctdtYdDnipVMvt7hwBv
KFjhB7P2UxYwDpltEC6cyjhzKSfFTfdceeBFyqZEQmsZYF922X54S1Ehl90yV0aOIiNIug0rwIYm
7xBfx5ciYUucV0LNGHNoQiPcbxxrHg/k6gI9KOEbENgccwzwySecn9hCgpuaIxtaJl6QKVS74vmr
C+6rAPuZx90r58Ilw+TRKTTQBcjfDtkd2xLFv5urT9Wy4wO3UDuzQLR8Nhzl5J4tmiIGv2pVic7x
00fW1SPNPvZqisPiQ+bHphLVotjBvSfm9kG9tQtAcmqir9omiEE98tWaojTW2+jUg0pCnI0rcmiy
+y4Sk9hQFoZL66DQvRLcRXwNBOvQMRaxlRNBsRhi4aVbToxYDivKuneN/XExbXDf/OjeU/FWozNU
hG+O72YIdGPyqTgFEWZiKbJByAdlZkddZbdZHkG9PEnz5ej0miHmwRLkvd+hu1FWxAS+1UZ0emaz
62hCZmUxYhYktRWXvGyKLqVfC+I4fPfrhxXmT+EK63HSoHbcZ9SYBop46JRh5fiK95ospJQSgsT9
fT3tB5NIA/bGysL8u1G5lixz9MppY1XbjJMRKEjdHm3rRsPduF/GVEgJ/uEYj1xbpGW78vgLj95N
23BUEZvSCYveNlX78D5V2Tt2R0kEVXc7ZzWYl/xdawzs1f53s0Nnerz5+SqVfZ8wXjdPueIUiGM2
UMqMtZFctXR+8Xt2cJZy/LYMkxGNFx31ddpHOsijbbNwRLV+uJQBEhV5PYIDn9bW7NSQ73PNitl4
LzWwb/k12wlQV9Iop2OQ+EcqJB8/rkRX1DOx1ebclR4Gj0aS4fHzyWQrrdnyyJg20V/lJBrWw6US
8XXfHU3K+Z75nD8EHWBA72io4QQm8YdO19tKjJJMfqCnfJk5sH0bm+B9HuXuFOhPatoVtZxxFJoU
NAcoxJp3qFjf1bX+JCp16GxYBCin++qKKiFtjvVJjZ8Ty+VjK00M5bLUZDYlhv5dAJqHmdrk7pUt
p+zO8w5rZA5Fmg/imncpnJw3YmdVhYEAFRzZZHz3fSz9jCFZBVsNa38PBzHiwM4S1HctUlUviYJp
l8bqa0vmWiUYYVItsWeakXAQmxBiKqHK1Db32yId+8dVF/VpusruOQ8+TlZqsW2hvrm78BGH4HMR
nneS7NLzy7K+Dyt74SrOOgmegZTTqZAaZpyL9Crkc6vPQkXMExu2DvFqMZvctE7V2BUG/tQhWyf8
Rp1lUTHskngqoMlKvRGJ1Ma5kLIstkvT2NYN64OaP21uuS1VQIWyjoj+u0eB4SjIiYhBGODkMUho
/77T34X3X+xZqFOsuiSSgAzrGbc2UkEZh0U2lKZTVHkNw7qJcAveFelQKg1V9PqK1FjiYibFwH2H
SsgmBpe+8AqbbNq1DZH1BMRg9gzj2NdGCiYGfL5dzW9+rVhZshbpaBeI6Fu8XCFdJ9G81N8olaeU
sqgOI7GESL+AVRohyR7yNH6ikJaHEY/6kw2wzrWRxHlHRBob37IvjnV6liSYz8U20B0pWowN5bh+
VpaK2ryJj/WP3c4HHWL2wyYaknKZd4X2nFvHzCSImMqluKUhuIqOoCps3SPrlW5s0DIxEH4ENr8S
liMXvikajQNvzdnQ6F86Dr/k0DZ1x0Cgn2J3xBgCil0BmXIaE8e9QcpxiSIWzphPWL+2GzHBPtDz
zpMrbD/yVYoZYDCJhe0FVZHQCfj5R5BNzcm/yrvWkn8h4PSBUduU5vUS2szzGVFSJqZE7EWlrD4x
IibroUSRsHYa83PqxDo0izzBBsMg7Wpq4qD0MdZ9+hnj3eCwUVotk/9Lb6+95eRB8Lh3N27mhS3s
ei4WizbO8HhURt+IrZhoq/3X0AZsjbT66IBPkus/8aEVdwJ18o5M9Osj5RmxwD6jH7PiArqiFFEH
0VeDNxjo2YPO048zWhj5rUQQmLPHzdwmSIqhwUpwT3v8M0vXKrs4EUGSbM46mmvufzIM3xxfN2IR
sA+LMVXI8GcvgaQK7fhjT22YNHIWZXOi0W4a7+lIC4UNiuoB7CrHAmfjWtbYm4/rDgXptcMJIq0X
2p0n4ouGTp9uOaeTdKYG/xWRISoDOqC2TpDKdicM90z2CQg1mfSKzuZIFwWZ4KeKmBGmn3WBg8mX
8zLZmqk5PKAGsm9HWW7DW2H7uwV/jHUL54N+YkQVQR4gEvmGLcJLnu1yApKU6ZF6FCGRw0aSGZV1
zzd7Y0sSlb2RGpqrnxJp5BVdRWkjjL/Zkc9uwsKHJ5n/xjvkOSKdN4OKqbunaQb0p1Cz25S/AABs
P/kiln/jq2kyyWoXiQPTn60L4DSFfLVGO/9mvtnqwDGOe3xhZI+IfQsWEoKXR2iAX92TuAt6NX7s
8GHEjbxyVDcXIa0rJWozP5e6jpVsA0Ra2y4LZhMUpIbniOOSrOJ7JDvpPt9budj01KSbAN0oP3p7
jZQF3XENJuVEF4NICr6IiheHPg/Qs7vH9DKu/EhUqbfopyCNAYn6+CgrCP3ua6xxixXXa+m1LgE2
QBu17/DDYswNoT2vU7zv5E8qqbIvOSCLl5FWB5AqXFjaZHcL/dTW/MiqNCvmToqpVz17oLSwPMBQ
Cqie0zX2BOtfoSquxKutuqMTdMIBmIERmst46B9j52Qgn6kbsqZkG4W6xccXyrjpDFAgY86AUFnF
JO1ruSBh8f0WjBREppv7wiefFMJ+n/aHgmX1NpJ9OPyIfUoGq5PbXJ1zB15c4VbwXsHrcL/SxcA2
MfNz/eV5EalEBfodajfHm5M2F08z1GqxTGpG2VaaqJkRNHGF6XNcIMTVlYumM/eaqaATSrrkkWMZ
0nnD07Dkhx5jl+alNS/G6d3SyIF7BBZL0nYbFqpGbN+S5W9PCOcLRgwmqKM95fehJlg2TAAfRdXp
8rdhkDy5LJvIiGv0aM0iOOtrmhOtxz/AcJk/YRlFHAzBQPQjZ8OxrF2EKQJb6dE7S1gTTmCTIcPc
uyChJzFXvuByt/2zLMwfAcIWwhdUJeii7OZwjvU5cAMzWE6RiK0z6sjVL6kURw3wLjUa6hvYmiTd
va66P+I5btuXPNmaJuGxTCwzBIiEQDsi54DYRPLM8923ExxKfF47JKroK0vx5Q2PfUEMiNC6F9Ei
xxuANXFOKRmrEy7Y0kmtDddRB4djsqm5+DmvM1xYSVKIAJs8ytBxhVLJGkP55nJLORDtrNVSP688
R7l9SJlFkbE8ywgoGrREtTBzNuC3u8o8JFEfpds2wA89fayjheUaozl2/h/XrjX/hjv3Phsh0wZe
/1vW+YM7anYvLUp3xRbuMB4JWogt/JBOFQpP26pDeIDd4h57WgsEdbP/jaTkxYrLcCNhq8JHk94E
n9IfO25kj9xks3VZujJE8gDoD1HKGKloB9GU9a49lhZyqcD92RAnMdNTWNKTg61WP51W++eOiYUe
VsvHj+dlpxhtqaCrSUhPtBN9SbPWce6cqDtKkMGoGXXDF9tl+/iaxbeg2v2cHfJ+UgGubke22xZt
s5blFVI3yItPq9b1i4uyl8zd8RjiMUkZjFE4wTuK/La8waKzp+4pG+tpfMHbG67CB52/CcUk0dJR
iaXiGO/gx/5cXKF5pS+HRJ4O7+CwXxh8P9NiiQ5BfkT7S1ermJ1ilV4kgYj63vzRpyNK/Y4ajLtH
sYQq7KqG6Tbe60si2R0WBaN+Rwi7Nm/83Qptb2qj4jOGdSJ2LOugI88/EWaiFXMj1PUa4pm8951m
TTZ7z8hL65VyfjleWYQGoOJx5LVZvFdoPWFtT69wTD62KzQUNAa3G8b2eoY8yVsDPRRT1sNuzf3O
Fmy3GRtRTP06rwGk9xNAK+GcbKMvfga6Xl00k+M5PTevzlO3/ohOV4MAEWvQyoJQ0BNwp9mvv/76
1jauRhTCXCg34h79BeSBKof9LTb8nGxKA8tNMEMQ+EakVukBBn5iEmYQRvMzTrCHLPihF1wpil1e
TMBoRj54foiSCFcPD+lM77IFQsGDNMmKVbllZgkW3xRraTSmg1TQ8teCIXot79PvxLRJYE53ZVf9
S779TWuiXuVy9CbYHpXXPA522r/hQhdaIpHCRjt5YJwjUazQ/KKT2t9ZVq79BiwECQvBqxNBFckQ
+lDi0DDSlcvAYV5PMe0PVROFmAJJdUfl2Q2REVLKM/aGUMsbPr9Sjsf9LZZiHTRaVdIiRUPaoRpo
rs2GLMX+qmjx9VCAMIEvmhAiZfK1KBrU0xR9O+3+S4i2SWxKp2JCcVU0j6CZt0o7sCAwwSb/+jgr
aBr2QGf0Vf6/xcPpmbpVxeP0DXcoobL3DYmb6gTD81WyFCLRzpzL6xrB4MIWng9WM4fu2+03vVLt
EXy3UY4vOf+y9T6TabxZtfcNFMyHdhLiY4eKiBUTuHQodSRSWHTu17YFUXh86LvUg/yZZTp+a06z
PB6arwDlUJyTvhMQE5V/0APJnQkrbT082taTM5lfv+J32Y0pUZiS3Ln3p3qirvHXLT5lzKBvAA8P
cF9qktzDZ4bn0n/h5LyUMXbaZDvU+Iqz7zz7e0H2I0WhA5KgA3nImZToLN8e+08evXLQGnNVXUQ+
Wf8G1t6OwjJrAYjvtch75Nft8WcVbPLBJw2lnHSPKrs9++aM8TPEVXowF8H02+3Y0l1h9q5ayn9V
iWpV5rIR8C7PBdtJ2G838/tz8NgCkpW1MD6P+N3HQFvc5cAdIv2BagxTHLWzPSz0eiuUahZTVM4B
0bbB/NhhLWl0JaNPlYbkzgihzp+RyvDaWR9IfzSnX4aTMgPZJ8Xd0eGoyREqzczAVMFk+Ym5Wuey
9d3zfpqgPy92Z79xBUBLkp/5HOR94nOim69n5vEWK/Ebh/x2TNr6TTENoXVLk4sQB2g1AEPQ28mC
1CN5GQp/a05+qfNEYdnIHcAR3sIJGL87cOe4FDtWrhxvFwS1ueb8CYyQIR1La1DJ75YjvoMDIvyB
hvXmBBbYhWWdz1rxA05YH2aUQXaUbA+PPo4ftvc38yenmbOuDo7UQvGJR9Nv3DilWqEPHX0DP0tB
wpy1muBRyreBQqEIVaBfzffmeI8KXTpncHQA+ZUc26X0Ce+s+FEVanguuM4HBchyeRtile/s3WAC
ElA51j1C01p5st6DUTfLADXBt9r2RITMsEdA7N+0x+s1qSsW3zN6vbXqNwF3d5z4tN/Y11YZ/e/i
bsdy+5UbVDRGKOQVGLyr1QS0WgigTbwuGQ5Zit/i26qr1p1q+nYhzqf8c73QYa2jqx/kBOavmhSB
d3WN3ncc4itEaJhN+0GL2XyJPYGzWineYbPicVcFdU2zGIRTF7Pl2HywNtlU/2DqJEIZNLR6Qnp5
ZTQEbttZuOqONWDtPZp3CYdOWziYK74xNKj9q9EXUcdDBUQJDBpDfXAQFca7lnVYRTmODHSQST5h
qQgtmXQBCt8bqcLXsSKJBPwQ/6d5/Uuhf8LD5HT5QtfYLtl3RP4tfWVK/fVJzI/Gif3SqxlrIDlW
ljciGRaSkdWuAQUcn8tlCmXCTWgVQJDU15G7o8LnR4k4PHe9ikKg3CRRQX/Bs/6GECHwc0e9CZL6
/dIX0RHWl3wNVoWFBQfYatVFCOjRBwfTdQbsQV8wVJVGVSPavqfYtw0JR99JWJonaOyMNaBJAZxB
+jzMG6UglY+cutKJiE9RajJY1Am+sFF8KN2C4GtZ/IrTzz5uGdj7zKZMn/bJEbpNwjRX6PIOUJV1
XHQVC2hp93HPnwEhjPMVh9uiRTbfa9uNL+wzxwUevFDbfVZ/7XznHSTKy+1CERCdn3rLZ742rmtc
RE30YzCcCuuHmHO4SxmDx3CHlayFZhHi0c8iUxutUi1eER5fpX3ineLhMrIntoZBJaj1oW7M7Eim
jOKMiYttLXmMYtyk7jmpOnTDHIPWf8IRlC+L4PuGhbK8k7gI44vwnlJ4t7p0kPjPppZKmC7BoN02
wDxDtG0lzL2ig67zpCbJgyRGhYfmy/5LY+O4Rqxmb0gdVdfrXl82DZUb8uzKp6JqVhNP6NzAbTKo
zJwvSocThSNjwZxuWqNDHjdyiQr3P1Hw8Y2i9pUMY0vRNKzoIbiD8RqSIPoy+FOhUsNiYhj5Ye2J
l5j68TKEfg5rvQ4hB6Ssmwnrsnc9n/ZEMW48/eoE6Q6hAjXMhuPwcrDcigtBqdXXSPt3f7LdFDVm
mnY1a8Hipofy6yPhpPtL+mbtxhednz1f9z0DNAyudlgwI/o5oPN9EHhTeCtsyLXEH3PezryD8b3y
EjilWz6h1PV4sMeVvI8MwSnIUlqsBEsuWx+2N4Q8VX3Nn3iAiAUbF+ORVWPWt2AHYwBjyquUVgt5
mcjLu3FyZAZc4Rjq+5DRXz/FrACyIg4O7ZbfNcXTp4HVXcDuNGLjfp1HpswB4sv/jzipvrn+jSFl
MBZF74zTK0i0Wzvr2CmIMzijx82rRHxNN216Kdn2JvJP302/M0EIX4/iNaNnTFc6zwsxMyrDDC1P
WPigeh9AM4VJieGkmuHDca2ShNhyxgdSRduuIF7udpe29VEmCL8FhFJnxjK+Di0BHx2ZaPnGhl9P
UXaP0LB35V+6YHR+nCHTMDInr+TqCVe7/Cq16L9Jvl+Z0k0FkhQQ5wXdazwtokQi8r+oy8dcMkfs
TClYfeYIdPh9KSNLshVA49LX9yfIAVH5EEGOcpiVF7ZPD2i2rc08A/lqBATOfmYpd/BdSs1CDqk3
MLlFoEJwVUin6w9lxOCXf5wMhg+3oAbwI+G4rTP+IlMkT60Ss1hoqePMHoGG1DCODdznkYRs3F5N
Dj2oXVYq7UIycQXxDtA2aT9aMCdvMH5YL1xeYNwBMZ/5ez9DvQSKADPqJp1VlDQwaOyrmE9LIpjZ
6LKryVRItWkJVObZl3DO0YyEP993fyM1ynZ87EXgYvQOYxFebL3OhpNp+E66esJ9PEtS32LPhvvp
MLzxD/J7JiQr5BpbMMzbKGArTwtnUcBupSRLR4oELDSUbs/1OAsKuSY6r06hikRdvlPqebDBgAN+
RJUJsW2JWG6srU3IbzGAMWuMP9SaITwdj3NDpTXcKg37AQe5cgfIFL3tsVXKDKK0iEt9BRsHL8Ka
anu+ssAsM78NF3EIEb4SyiKC/+Z1Vmsl84cV6NSeW57oElD3n1AcrPH1ngnYdS8K+xw/uX5+Qpdh
yl3+ypTeMdiElzpHTjcQ3oKVGC1eb8/811oDb1z2eTZ0+3AeuvCOllZj11fA29D3fIjXIGr+6oIB
NlrOwapHkd89WN7mLV/DxdMFjz8jQOK7XQhL/4p6XIMN9u3PtiJmPD2TDe8KT1T0IB9BVPO46IjN
VtznRPpwBNkzuC6x1X/vM3xjzwL5fGwJbCalinTy2ZyqHctM9M9BG3hafnQVJ7kKSl7R90Q0zM0V
utAULlgU4FfnaixOksJW6guIjYFOQ0K38UoeBLB9803f6CMdTvJXfh8TPbqKxkmKCvVSNBt1TMTl
P5akvPm/f2n/Daio6Xt0ADo6S5pheEs5hz/mKS6Okcg07a8IgICj2Klpnvuxnp+6NFgbAX06wTfi
SmgLIkc77apvq12EDnhs4Xuvy4B1aX72m7/A43d8kpgMcLsYgXVSbKR+wb4kAYBfE9mnjGgXR/M4
MFvB0bvmwwj1855Y+PVPW3zVelCHrP6ocefOF4kZsxn4dvkhIVV3vKaxUdA/FWRevT/LG/BPs/NH
nU52TYwU3amigEnG6N0CabjVKtCveh5fIt3MlS5sbf80tQdrnNrLTeTuhqYshts9opnmKSq1FNyH
J27AH3vpFBQHDwXSYhBxD9hawyhLgbxwVMcqgZNDeDc9XlUnnBddNSHu39d9eB1q+EwZ8GtKlwPy
3z+Vl97rDTJdp98ezcUCqhoTA65xp0n/+YLdAkLzMJRQtRtcYeSzgzWyaHsGFQdNBYNxf2elX2fE
1sFunaDldwGW+PNEUQAgWsH3y/DJ1MNlxP9NMagF1xX+qEFzPEfvLhqFKDPt/fAEUEDYzSS8QHoV
8YevBg26h6P1fLdBKrv6zylsNBmPAi+b5U92oBX14NRQ+kbhLjCSlucUYfARyGmfp+kT30035tpP
e1qSgTl9l46Y8XTBrsP57mP2JJsexm3WcoytLsmWFmkeRzFFYdaCpc1s/ymgs3QFs3ILglaBdEph
DOlvrZFh3f1ZxaEYHMAsAoPfNwZVXeY6OSQlKO4OPEiPzJIlxx2Hdo92y1id95l+xnXhjShNtXeT
EDsDbhUnLKbs358Q7/jhq+CuhXD476rcwtTcRIp3Vfr8dGqabUN3S+PAZzhyQbisqOL6KaNmNHC7
jswaSxM6Wvf0F7ujJ/E430XScZVl/CHebwZjbtfaool8ei0f/Zf3RvKcuhPpvdR6Wmfe9obtBvMH
elJvITJTzIo76SER7Q62QJfXmvUYkTFkI5K44DPeFDxcNWNPCEdkIH2/g0WYGBEq308Tip3eW3Qb
Q8vVGVYfS4z9YFV3fEvfr3xCMHmcA8pJC887j3jaLUfQlmdvSHWFKUUmzWg3mvwBemZSoG1JucTE
xls0pnDIrDq/Q+UJizrncEDQy+XAmB7kSSl+yjRRPy/5VJZh0cb3ZrwKJdKHzxmSYkc5ApF0rKHi
3mT3FbsVlcwVWL/BnX+Ut2ebZ74GYJNZHUZFlTkUMSPjkLNDnB8j62XRR31fF6brVOt6SWDEdRe3
6wFOZUZNQGXatsCkzVd78kmJp5bv4NeKck2nLP1heiUQiMUtpcc1DOrK1VpEwo+XRZZcXYIWfwTg
g+hG2cFHPTYWdOZckNyWuvX/wr+J2tVC41JQwwbTiVIOS8UQ6hZDywH++uUUBZLNI2Ld1y60jV0o
MoAz4d1eJCTkT5+LuwWMcn/s+Wl7MU7ML+E9TTf/af9rRPLuxQNX0i57keUQgwT0QXUrAAS3iRyg
88339MonGWZuI0eOm9+Zdk5AQKwAEHs4R/LFNP3e5Ve5ob/usXpaZX87VoXOp/cqkvwLwwyLlzRu
VgGc9IPBmn3v4T6QKxsbPMGDzHLdl4ol1JwBbRgWdLh6hA/nVx2qXC5YYX32kShceGOkMlQSlnsQ
yAOF+Sj4eV2VngT5tr1BzyYYAG1BnIeCHWiiVDU7NHQFgQwFNvqsu4b4epn/RGK1e03cqm0JgyJS
34E9H0V2KqrNAvhcgvJeedoP2tzFj6HLRf9W3D0MYHYvnRDsARbhkM2U1U624P+IT9ne8vbbAMeh
8rxlmrgkvJGQoh0uwcNeV7pi0ay5fmb4x/XMcswpqCdCl8xsjUwtp6HSdDWcgtw7DCK0ns9UC5Y4
vmdL3XF66WM4+acMNbF6CAfC2cbLNgaUHxYp2VyEUyJs5NE0KbcEMaY9Vf6N2Mr/cwIKQYTxooji
nLGnFUNAZM5j4wwL3Q9dYH0byLVGCI7NL166opFzvKhuSRYuG0MAvs6Wm/N197/EMMhpezk+duWn
8E913SQO05dPMQOlHfba1sOUUjc19IgPg5420IeEzjVomUte/cr3kqLjgq77p7HdyqdYtbhB+LPA
o05HakqmAfd8yYhbrVuNHWG5rkTmTQGvLnQtw1ru+NdeK1qRcAPN7xIL5LpNaE94mWJyDspnpjlB
/oanIGJMhh+Z3jjvfGMA0qacGMoJhZpJPkC4N5pQmyFecJT/WC6Za1aHKjjf+n8wiw3fkOcdmqH/
xFKTZ8rHV17Y3n761m8lOgzuP5dRzoEBqrgHL2xQ6V7iIJoOKvwLjuTf/ZFDvyfBs79K0x7U6BTu
jEzc9fYVO/aFzbvip+dU7Eqw/PIofaq2wJSRNtB0PbAVDmLFioXSsyPkIaUa/2kg2GHQEP03wgXH
gOp2DWFFVUyMiA+0VCHC39fiK3OOwiPZqyduo+lyWMqHLDUwDDPeZV+PLKZT+voK3IYXg7/F48Xr
2QrOUNREPfEbYyuJ2szpwxKEkVNvD2jsUFrNWFsuiYrfEf85kWBzfDm4kq0Tplvktm1jFheFco2y
FEo8FsmYvetO2j+Rm6YMXDCL6TnjSKbWCe5Lk+JBn0YII8xf0as2B5TB1Zu/OSk3qOSqpCbx9TzA
dQCJxHkaciF5gwLtUxdQS2A70ePN85aMuAJ0HPnxLFTorL/PPSctKUXGWXZKdsXb+mArAjlu7hPK
5Uj1PGCCo9UJqMjqJLc5GNVHuJZhBqKmR+4wwZ+5eqz5ieblDP6jR9ckwVyO7wcpTCsGmSqfOobX
vxTr4GcXpS83BjXIhcjRGnCHT2yQ7HHc74KdhF25LhUlGFlhMAS8xaVx8E7wdevgHPpl4HPSCaDX
Y2tG8lAd9tu5tY7lx/A7zYyNkCcW10HJ4+jYO7UXvlpNQYOcEkENwuP0HM9IsKCekBAyvU62WxOS
UyVDPBrC/bRhOvbnd9t5XdHdYVVQuyHOfgIoazuLZFh4f8KBK2crEewfefsyYQJ+RRvK+HXhpulU
4P22c46tB1RWYh6isBYniTRMcCCvHmfZDu057NClrQkHl2/MNvu3iYgCMFLs3rk77wrFf/RqIZea
WSzBhVdZgZEaqoYvi4SmSPSlf1gvY5MWXM6WLD9FdKuvOuY+rBRjD9BllcBxJMMJK+SD4djtOedy
653BHoGxcdo3H3UIX93+LzKX9wlf2wicZb/OQZFfTRVAzAkbwOw6LCKU9g87/qlneCgQFCrHYEjf
ZoWQWx0BsoPJsOiRajYkJeGy+BEAy2huYsOXLYnf4urDDaRQ81CIQ2K0LwMWKztEOv8ALyY+W0+e
2LpMhxfMx80oNUGy6KZ57WJHWv0Y8N/OonafHaHrK12QHAc5k9zOlBrgcregRXbnMWMUpZRDLaLq
4/wW7NJdxdKGYXgfW4EEadXdIrPWqkZtqNN5MSVmSot7qEwcFTRd/UkUHDV5iQ/DaqwNswprOoVP
L/n0e83FCQeIWWhhs/ogvKU71oHYn4Xq4n1MF2xeyaznoD4KeVHKwlMwryIWWmDNkbvhJQXyOw64
jF6tWrVzquPXv2iZcjqUIIqeZ88Xl37xkXDowaYwZr13/utbVaTRc2RNd4T1JjETulsnif6kDymV
ZRyIXWc4EC650LCMbICRnqpMilJsmI0KdWSURlvePcfBcbmM7TCrj80+/Kj0PKXxqZQeDbJY/VCz
TvUTmqyBAMoL6bcwEr5SpnaxWWM7cve7gmfwNqtfE2DhsGC98S9NzfOysAv53hN1vQ2YZzRHlgMx
pGHFkjz2SVe5Qtef7hB6AVselQXQTanEO7fAGL7k7luBLSmSpMgdKR7rb3b66hK5BuJzgPkfSjf3
I+YhgtxN7KuePUltuWMHKFOfPNeWYJwdiSwHAY8uUTjnUASnA5QlXzZt8WCWlwgTwzYCEaF/+gqx
wWy/xCV6GCxTnA8DebjFg8/oePEUBzcgqfMe0UhapzDq07gYq3MYnkA5GC1jfriuSlxeZmHGd+Sc
5C9c67ZdfFSPmsE7Bz9zwNr5cLs1PRqIkOq4oFE1/vt+7LsrWjzVc9vyPB4+tzhIQzSIKZOFWpgi
GjvSvF21JN60zvTEoDnQ/DxzqmjK8kUrTUy+aveQS0rUtGXNzXEXe+HcDc96accNFVyLF/VqLWYi
p8mM0LEUIRlP2JYCSpCEUtn6o9vXyDpCgVGjnEXZH92ZAoumFr7eOioh3xlvz8NUpTUuQB8uG3uO
gOu1GQOq7ryo7nb9vbtVSKCFZLi/4ZVpTRcd9SSOYNKlxhFOuqAk9oJmEVfln8zbs4ccB0H8dstU
ljF9cFR1B8aOVhmxX+o77Ca6Ieykj+Wz2OXo3kdWmVBOHisdl6oL8b0hiGWOvT3en019I+RdQq8P
FbdVJLCF+H5IJrwNq281q45AbtFbbKB31maj2UNF9mKRatoAMlEv7ykY7SoIz2uDWjG/2evFcfzd
mREFzG4Vwkiv6/jtyvQL3rMVfx9Yc8q7QbQxBGHgH5kz4hCgPylOZJx6lNoEygOQIQ95KxfE7mwP
SMf1WOyfDIy62O10Q6v85G/yhyc7r5UwSXwJ0BJqqxrR25EkNOoUY9ykVmEWD5rYo2k5IMEtWG61
mgf550mHfu/1UN1QW2BVcg/grVw7BCS7/heDfzTQXLlfsn4dJMv6Xk/1dUI8mcUOc2ja7Q3wubNg
wxG/GUQBp2CqcFdzjgMsUza5HBBMefWwfzE7F7T411Kt02LsASdI3E2doS3911KNLqkw9zjIBq1c
NZrzKYw+vRVkDloZHzxTH0l+UCkPhcc476THWaZtWVgWDon9meNvgiYCU8hxSb7MBwdiUAUh2r1q
jQVc6RwmqJ613RPdMqmxD4jO80gRTizqViXSgoGiAzXPEZ07YOWqP5PTUELd5up1PFT0w8k3dRBK
iDs2R0owZ4V8paxPF20Y/ifxoXKhCIsAJJWQ5YR2TjkwjyXrS1uVy2R2Zxjna0LCrm4IXUs5lW88
Xm48h50vzWn0DhLXVjR9RDhFjY1sNlYCkEDXjam//RmREu+yV3bJGj+v6xks2ht3g7Tcy6jQp8zq
S0o6ybqAl+A+Atmf0326RkTzQ/zTvZULgxrlKYYXs+GexFqONIeHfHBWIAglfjkZLpoYeNq9MfHX
jb4MxMO/jzR0W1xq4dcUPwS1NMxJPhj7Mi/bSGvF/D7NJ+Jc5ar+gMmiHCqEjO/ydEH8Ujs6iHql
Rgc6WB7GtIlQ4Etu2O9sI3h0tI1bpsbG3nxjz962KvJHALi+4L3hXMk4T4kcn3LX2c2W2mioco4Y
/iP8cgqa7yKC0C6HslwQUvYuS7qXHAA1ysD4H4Id1V34B5zhhelelrIFcNfzhswKehijAzYOP+55
8szZvwOahBVPPMxQfZqyuR5Xs7+8zIy9pkqelJjxeFibVuH6UvpnEwy07qUf4GD53gpViWEfgbYF
iRbGUTByoKifccc4QRiJytb7bKONmeqcIUJ69Ow0wlkTc3jIdf6SaiN2A3ngC8Y5TasaCocJRiqY
9ghsY0HjFrBDAaOefPIR0115D53kBb9cdMkfJ6ItjKiHEbGWmsbsiXOI4sbWOiMNnRe3V9lb+YdK
dldGsPAgyw+lLG3/errSZ2EnQa35OpM1eEBYBUx5ZlLTZdcHIn9LWqRpNzwL8mlB3jrIFkJ+Pw1t
IEInNGNFhik9v6jWJmQWjTu1YiwXEYJClppiAlOgsB9JWUTR0gOBZsAJGzZD3W9ST5oGdBeaQWXn
noaxE4MTmtTkpxEHrxPG5aYKIRXI0xw10G0eUkrzIf9/CSnOkihUZEsBcH0//PtpU4+Ui6WQ+Z45
UTACsT9VtXGwwaRRZM3WYfDafuAz7bVAlbZkOMWse86oyVnWUX51qr/vjEGjYH1gGEePStGQ5MXq
p2rc2GeO2AsHeJe+bb3QUVVpiE9ZSffq4DOCOJ6ffVTln3Ecpl60LNNWANHT/s9ySuZB97oOIT2B
llVT7MyLbCBRpW4X2rQBEIp+KrFiLsX665nuWmD5iUlblWY9i0Pqixq1iwrh71ddbYlmBBiEiDQI
/HMFSOrZ/nxQYa0583rif+E+TXMZwl3OuXmKAOi8yvbvJ7v6o2OrJBQtTb0BPB479ZzbCxHi0x2f
9/Nme+q5kgjoAS2/edXGUf6IqdmJBFjYTUtEdXrJOBCFgfvl8X8ebd31LKEVS7c2kxKtM/ddbA0S
9Kr5m1GETIYnFEREhylqMTZyWbuqQ1WUHQ7ri8C6FAWM7YQgbB/ONOyKGMr2T0Ddl6RKMjhTDM+u
3loT1h8zMMkPHHGG65C22a4ZviCY+XHPy6StpNbZtiofyFRmpYQI/aRAoBWZvrdrt5JpCypsqRT/
1jc7/x+tTVFVyL+47Q6m1vwzTzv6o4TZBnI6AzFhU5kaNlK2tzMD7p4asHNmwF0eVscNhcDhF2Km
+4XhmCXSnc5iMWHtYeOStM3QErTB6z2ixgOrsCg5nH+t3H9aiGlQ/aGRBFdqPyWAQnmNmR1vxqWJ
uWhcze5Avj4Odn0UOEkjCb01gSbvgx5UwZbwxXYomvvDqqT0urVH9Oq86o3HX94i5HggpZxR24Vi
CSuYf8uO1bhxLAoEY9rllmWNn4yQ1M06HhnNMZnmqaGq7xz7l0vFGweHFrz26Oh8cHXJIZf4S1OV
dgghy2qEnBHEVrIoLZm/vJLdarJsZGZYszOku9alIJay3k+kmwXQdWE6ncSP5NSp29OUdImZe17v
dQtyHTGItkxA8ww5v8Rpp+ldcFVQhT7iJUCRKQvwgUOm3Nb7+IaDW4bDRkQx6AAiWp5/oMnGWfBK
bM/sYC36Pozt/tKK4UxYg8PQWo38PYmWg/0HyE31tsXgGRGlgSc8UdCSLmYZfIsrK4k54VzzvZNp
P6l57neTylrM/r5/f8liFsI7qAI0IbUvFZXYisiG+gbFpHLKnQJVL6wx+xwIO9qrqEPrQHgl9jk7
Opy3kEy3NlFC4hag/B0/OEdrQIQAXT1/P/2KC2FDE0BfXIN+0A284WPhJoFwZsvvE+r6XJN1W4de
d3gM1Sp5upWk1M7Q+2vTmLsbc44ITXqdXRZAd7uCuDc+01l5yjiNl3oT22MUjYYJV879WAJq5Ds8
YgjcBf01C4N+h1LUZaK50qcQzq/XyVHpAGpvCRqsbXMkxiAXfxZkSkSwgLrnqdWmsWHos/cgD6nK
5OY6y5BDsKCCo8XSCCQdBhwGkgazNiMGenEVnJ0JpGSE4rQ4bDWDEgwLscrmwOFA7AarBBCe3Fsz
xDCfjpW18eNuQey70xkOlug/Mrv0wmiANgrqAfF7g98lzCnWwNlKBxOA3d1IJfnbq+uzdPco8gbi
H3+JetH9rt0f37BWxYBsxixudztJmXQWH/3fgzAxnujnR7Bff/nH2mClrv8wFHSRnq2Obc+jp1+1
SBQBkkhsS06beK7AL5rRPXIPIxvtZos4ImyM9ev8MNvkge1pVnTrHeA1y8Xn8Zg2eOZCcfmsdv4R
j6NGRZ2BNXQotsQ+Lt/GwTxlDJdhpctY81tEoWzeBQGoUk4jHSZl6DL8MItshMFC3MmI1N43ELsx
29lmSLyNvysOVSfllmg+qVCLCId1+cUMuyobTpm+HiMKP2HF4L4KcM7+SNvBXGVgM6gW2KdcOiSu
VZAPUQjifYx+Rr6z8mkxSjhPidM10MbGqVav9Y18VbIpGkxNg/badCYw2ar/aqS+e8S3Npf8FwEa
vtRnMSlOTy4aKqqX/O2+Nbs+aw7Sx4pTtFEVTFAQiUW7Fi6MEEx8dkTAZBdDu9urj9ipCn644jog
bztzYIg1HLUf/kjo1YSVC5yv6W1UKw9zdXjiaRIom2cRzeDs5EaguQVeg5+vdwufsqP/jzCln3Hu
pN4Udj+fax89FhxNpT/iNIeA33oT9qgt6udBZcUoqv0Gv5Z446cfCJ74YJYOzvK9+BD5AbDibYuu
euO/TYzMtRbRYLlksK+Htpssm24Cvx49StCy+qMOQBeHFBkNAOS7FqpFPZEaHe34bX3Ewwhh7grd
U64OlBPXwQt7gUo2kKvZGFGW0DbPaLwttC9bNm5028jdKKzFdMduszuiJa41C+L4uSA1A0fUf/Ro
yH93iIZsiXzM3aejfVVUyAEGbs/Y5yZnDWTfhs6EoJZ62Ytvq0n0wiH0K8tuD6Q8chSYCZyifbZr
XzXYBZl6OwIfaEK8qQYfS4+fEA/HMfyypPHh635Rlore27+GeBDPBp2MbxeMa/9i88LXvWTZzC9V
vKritHz3w9fQRmD27TF/qrHwfJ/jfQccnc8GcGClu2qSQqMhu6/N4egMqf7v2rDU3dahXe/Vmbgt
gAiA9NTlvgE5+mud6hx8TtJx0jx0399i8/dUNLIopckNb2hGt4PX3nK2f3jo2pz78U515op+O4OF
krhgfs+h57IGbLEdB6i+9WD8reWN5T+ScSEBQGS/WGmG6zIE19sewWVm7y17kO478Ce+FQIRqYCz
lny2UyYMoUndBkVTgFT+4xBEV3N20TsoVojwl0jjCkAd/Obke0Cfi4nsP9K0BtyIJ+w7U5N5lVNo
tU/DZwkYdDTFP1f9kFJSG09GbQ3CoUcOSD8ez12KRer8nNxeTuv3gAYyzPkn/xCHC32d434bVG1/
td7ooOb0HFlh2GTZr2RQNk6zVy6OsXzYSmJPvUQfT09LaIKAYV3wjHH3iP+mD/6HaYm285hYufxH
mkwA7ywCXUQSQ3Lf0kCs93mu4Vqmq1y5qTGGAnrb+9ufnBr8li8VTlvntKjB9eGCqKFryuo9TJMY
8K4ChnfQuA1o9ET4LBLw07o9FDoh4Nd8RhlbyQkHoQ4Yt/pFxzZyf9nbSrbqVPpK/HH7ZkrGm6Rp
WRuCSeG6tFDX7ZiWxw1U70+KVf9kbzk4/bNICpjoCo85uR3ieM8eWlTnLDI8LghYDeipkmQ52S+g
RBi+byPNU4kY7Gjuh1GQQieJTO036KuLb/17ihO3jeUMc5Z+BZ6W+igmw2ntajTWMy3NbNO7fe6O
8LfuUmPnVz2VUjIF3cK+tK0sP+AIWI4OP9PTxQysMwWY5wSbb6nY1SRzAqgU9Veu8OdFTirJRe2N
SqfF9bkeGrnZ/1QqU4rPl6Myk/hMSGmWZm8FSoklVqLZIwPMvlsTlroIyOQer24K5ZxpLgto2Bh4
JeSF3EzmG08ZQ/J1TVnTjwrXGqdev5F6hDXAMvlH7QDqpcERH2yUptALwhErJtv7Loza+0McSz4b
I2FG8HpjZLBVWVdepqMt2iKfli9PAaE4Cfx02jmvGvln3y/zW6QrDCdwRcon2lz/WxAeOWRrOgFI
72zJmMGJ3LoKMfXnqnAFbh1Ot2/kdmLIlLsBdmA4TkQ3Y6xVwhpmXYUfszPC4eRZUbSsAd9RXb8j
DBPX3pi+TLj9if857z2WGTFiChvOGHppMo4nMyItrhqgYpOxMRPEaEX/eFUndL7xyxgGGByAou+7
j3wbzJRZ0t/CmkgY20AOozesDyaj6uqWoKozVrrU+PRa/HI2ZFsbQEYX/RCTzvBQ0R/IY9Y0nO6p
YbBXzZO5KpjFD4Dn23BENxFTqBIJMesaRwq1h1fAJVoE4vzu9j4MN9DBH/M1bWD1WmkhW6+KZPvY
O6Z/cTWAmArcVWuzvib5EEJqiVy2jigiA9pObqd1i1mQIP/EnSnm+eQqj3YlJKt2vykZBSz121xw
ULMca2BoC39IpHDOjknBMR0YOT5UYSH1bxlHoUh/HCynzWRbGejzNqs7uMZKy03+vVScP6QxamAX
jfN600FO7WJ39AXL5mIU2sUasb5C4L3jOpUkEDUsDZsf7N13xbcAurrCWtxI7d6FAauqL9q83iLs
bNiM96BNZwzfvHVJHLY9cyMZp2lMaJjk/JDjDj7KsyCTqpJAeXei/Lm0nlxCVa8P8vfa0XcqfUd1
FBw4F6dxe5D4TWC8P19r0PeHjN0i0Y5r+fvbhbgCFCoEMKR3lfS/dXsExAWTFhojP0fef3x9a7cM
arpo61U/tq9nc0ZmZRaN55vPGC3tBWB5VJlet1DxhtZ7ZR1A14DhJFLRUKtIF1h0O3XfZSaK6GZe
GO3FG4/eehVIi+fGqKR9jBientFjJlw6bXRUsfZHCSNEk8laSBFAMWqzAz1GLHol7kjeHyN3LM9J
0zIEuhfEuicle9knXxwMCcCRiZN0aPcG3rpjW1Ok4Jwt9jRBABIWxpKADLexhYbxjkVujvwzy4pa
eDdXsBmEzCUXtwnpNfn2EwmAhwyw7aXvfydI7j6HFRpdkU8bxVTOqXUlRAF8AFkployguUf+A5ew
pqnNsnz6YbA9NU/PAjCdW7GxMqpOGfxbuhBcrsyKV39UNhOtL4KJqCoGRZ2wn/omKUIXmsTTyldE
HgRoW0CIuYlZg5KYmp8GMtK1KmgtiYEG2FWeI2naZM3ZfnQ1aX5gJG6SQmrbU/uAF0SubrbhCysD
wY/YmuRlNK4FAwZK8uRorrNshISkdKQ52IhiyIK4F56Q8+RuG3l8Q6/TPXBsBAFAHaq/d1voJ0UK
iAv5IWLx4Hwqqd/SXOzTvuWn1ijm3tCExo5CAenGL5U+7Uy+fPwJ3ybm8qWkI07X1tkmR75AtyWp
c/koYaYLPKuDnNS7xCVPZ7lMqmnoTI7veOy1aTBWUqDQbW1vc/Poafv5bkL/hnjhPo12K0w/lA+s
1zGZ6dmUzXlHzDdmCsVUjg+Z6dKrJUcvNcNcG0DfJB/bWNRqh0uWrOC5FnCPpTAnAFa94SH7PC2u
l/cK75sLrBxrSv9i0vwmgvX/lx1JUv2397GyD8vK2m9y6ffy9XBUDjMDC5RyxxNE5TGg3ELgx1Wy
2oHIt0mRneGROPB85BXLYIxhAN19net8CnotPn/o42wU8YTogcsSl26APkB+D1xXyyrCnzvtyMx3
kz+UE26ve+mWR3UdXEmylz+eg2HpyS+D9g7m9aXEf1PqWQvpUEX8PwHwVvUxdmbhDTR8AWg2yb+6
iyV0rf6Gsez45Z/fdMzd4cxivrfie/dVIS6zmxXfzHR99T7SD/NLP5+/T3rx6hSket77eM0KKurv
+TZJDNbrE20wir+6agEY0rHI3HbBVvdD24nCWqx5DRn14hyacX6YBCns7foJVq6ioojritTab5sH
ribgC/1GEMPLK2JgKUaU22m0F1ENBNx8LNb7AvUCcF3ZvdP/1tKPqGhF/VqcFmFx7QcC21A/q3je
lenhEvGy0Ptm0lbHLkyPAqxfoycW+7TkyMfyVl8+nDl0mvD4CvW9SQM8np6rUT58eE1nS2xUSZCQ
L9Fn4Kftt3E0aGoEy/JG8yujdiRXTWcaYTu/j4yurUnd+8emCDANpXN5i+Ucjb474jcFb9toGRDb
NXMNxhO+PeNjjTfWTR91zG7MOEFyXcHEDW6yuE/SRF6oME+QhyPf6TQgdQPE/3t7l4yXnvfa2ppX
9A4pBEwKpCwqiKIokWjDV+3gBTJQEitoA/7DnCJ7gCkh0Mura4XEu1acarCNmpAD2wRbv4DFoht2
KmJ48wmrIqAZHFgc3QQb5RHJpTlY7Ozr83S5gjQHptz26pFqCIxXgBXLlE17npydn+X+IzOlXA6Z
TOT72axF6M3TLtn6tQxWGmSTaXEDSvSdsr+QQGCNz7njv3E+3RDJG7UalEXpP6jbMey9ngxkoXpC
ReYro2pZP/VQ7Q5N6Lb6p++U7lAwjarFUw5T/VaFBkRN4FBoH7dLIyO5BZGQxWK64pBlzbS9UI/v
sV0ULpyJHxYutvEe+kFMVLe6W9MgXb3g0JjEzaedzz15s+PhQUBrh3hG0Iic7s0Wu9Lwmd1oTOxe
t6AofV3IxTQBoX+t6IKAmSOIXsYFG0m8j4WCp6vEcgV23b4JZDFK9HCZmgIPONU+pr+wgTP472K0
LsFAqfVmuvzJPWdYMz7Ub/hd1EsxiQLSBSTQrNW6KMTjQiS4v7PGkAsSrRAOd3krZkfUKor4ggK/
OKvTzXKhDPqw8AasmXPTcjIro5DTOdRQBvumh1UaZ3ld2Sc1D5qN+jzkp4kk+1gpyaTztVd9GRCE
v0U8E2LOhdgkdNrELxpO4EO6ZMvpXo4Efmjwr10hL44G1y95vg0sLp67wW8Gv7biy/CY80Tibf5l
A5rXP3z99YMnYV7xbPKJiS8JsyL2jz4HwETehbPXwMhScd9zJ9bQs3izxibGJBp8sB2L78Uxy+n0
nRrF3z+PXIkhedO54eOVGfz3nqASl5IIXtnMqO4KDHe/oDR8eYi5SEueCn8hS2bbwjmGZy12/3K3
SLzMM6Zqw/Gb/n8JBat0/e7netUTsQsRiPXMA+WoXdErSEhGdRVm/XfkgyTM9E+MWTD7qt+FXkcc
SxkOEkMt4/HGKe7xRlWQEG+sX2/4rfK1IuPSdZQZRgqTkgYfc37CcIiR/Cimh5MnNtSYh+yxOoFL
4OSfimyXhiJAAFE6PNU2Txrun68LPUZ10gqfq+WDFo+WWcgPsF5DraAsvD+v1U/IHnV1OvEVUNN9
hI5n939/UUX/bkC+GtmiJPxIjpw0mm8g3XuSnYe5YMJ5KMCPS7JQO4wiQxE6Xzgc3NemP+s1cB6I
JJ/dynCmht2v5HzyxuBfuijctFRdehVWlHetjqZlj4AtWqufMFm+AYcnVeLfxnHPdRqSvX+gUMC+
+KQhwHBmz0IyxAVXX3xHJHo1Nun9K+AwpF4edRgp2BDFUiade9MOh8Miz1JqIZMvV5L0L5+NzHv9
zzUtiarf5jxL89Q7bVHoehlx2sAiBlSLI94MKu/ZWCXI/QII4RDTGlKJ9zDxBj0gbqdVeQqNEhL8
jG186bXM1gOumKkhzfiYRsgb20srEnhtT7losMrKXoSPPOL0mtFzpOtNCCQbDXC519777nRzRdSj
en6xxsvsMDnJburN2Vis4IrPJkiUMxfu4pU2+A7O4xObxlbiu54PLKttcZqeDTCtVZKMfxnQE0rY
yrIMfnw7h7i4m69fY0yHRDdB5nrruIl2PwZLUaO/Y4kCNhyP2Lh0ypFhA7Ew02/kCOkiJaGurcdQ
8TR1+PARNh5zKCminOlnmwU08ttAcse93ADisnpjYfWNWvZJ8EgiHpmYSZcPgaFVWm0Ja4UH4MHY
qscEa4N5GKmgUbW6eWuXBVpURrE8WuaDVeovn4MtrCrsXO6US/RDQm8mqpYkD1QPbyQsXW3hhQ9v
BVm7KEXbuHQ1+NAC7kKwTNud66yu5uNrhAR8tg4RP1vYpa5bSF4WboeaQEP94u0VPH9UdCr+lWNI
eQBMDyG2D6Bs95k1375xF5hRTtjLi040xVDog0jtqqBVwe2o7i8/nxzJ6iuxPfLLq9ushwMFr1ox
SzL6FB0COKJIANpTEfYy0ku/KMe3Flgng07TpGy0HEah4kv6xJezvE/8IXO6beoajAQC1gWLOKUR
rYe3/E5FthQ0BC2TFM8XnUia8EALipSE6cYJqCBPHl2YR0L03Mf1RSA6qL8k8S5QXPrEgN0o4Am8
7m9dVkAEM/2LjOZb8Sn9Twx4EZSYT9hBv4FWSLT1Gq/BiE6KvoTBktnjW3A1wZkiyBIJHGgFse7K
1uxL7qVhJEaFy5Na7DjaNTi4kW8Z9OFKM8bnxW76holmkVP2xZcYR1NwwcX/S5pqD9F31warvGuW
pdpBMuSi/svI9iI5PAeaNNNlrqXnTttj4B7p9zp2oyiW8dEtIjDFxyoS3mLESHk0ESA8c4ZgVH4I
N+ar/V6WJN+bOReD4RwpCzGtekgySI78IWfumBlFp2qzeKlAI5fFZoxukZdasaopUwE3pqzyApMV
XBkxJts5VEVi04JucxRDYM0xOrOdQHcsgCuHZe0LWn707QWeXWBOME2/myqyFiJ8N5j7ext1lQBU
N1ph+6C6ommei1bsD/M5IT5dMBPfvzoAGi52cij22UJaxrKNVHqY+NMdolmxnMcJKXP9HUTtGxzM
mqGIHE/ojnR+oOWKBW4LdEK9wpm0j5uyPp0Beb/6e51jAw6YrDX6kQO+VVGIPwANV8qkgEPWVeN3
l4TXYhE/BUdp9nqYFW2b6ogYolQmYBRuaC/35sWrXjBCshHweqXadwmYk8lDcqO4qF4aX0hXOSVX
CJTd9FgYRCXifjSXdTCz0mtqTp9sEFSMYm/Vo7ZjgPNwHITRXa2hx4G6P/7gGy7H4GMhqKZi5VNg
+f4JQbL+X8dJR1sECrjt7zwRTfZ7DNE3ONF6/BBW1VZpCkc/7MuLprcbgjYGJVq69w0WRPJnAukk
CeI/YUwhCrIxWRhEl+MkV3VgWbf5qqAgvWIigyYbHPmhXJe4F00a4i2xlPX7ygI8Au2X7TQBwB2V
DLHmQ3GavrunCiQY4OgmNqwq8QQ32Plahh6hKw4xlfSGhRzllzSWVQOVbfW5LJJd2c77Papm7WzA
Pph4ZnNYeVRTXOwbyMTZgtsl1439/EFgglPkoNk/Lc499bT14ug9MKpgv+cyG84gPtQk30ENbtvK
bupr9AbdLOBx2gJ3cz27cf135J34hMjZ8TFXVha+FP+XEFOFa91pJ7Hyr1fnFTNtlhMGI06LTHx8
y+DEUDLksk9l+CTRt0OTjuB/kKx4Lf9SOyHsi4oe2QW2bStIbxSFUZbHZShkyaKaptE1hJxH68kr
++q4O+DpQSHlDCbNPXi9fDAS4abtjORTBDCtPpOycdODGIzVbHwxh9fJV3MCz2W2axXZsY+Cl6VH
y3hed7WsXdQw6KiiAwzUCwdFQE+iB7ECROORJffGFZ7OLq6Ks5j92OZOLpOLB/HW4S8VaGXLRCQN
zY+we23wrwIxmI6wTWtzM3bNX16S/3EYKAs3d1rKqQPkSYPRHW+WbNAa8oZvvjC+7oK3ZLpzlm4A
CJ6CXNT1AJ4jKhNxpEEvAtTFzry5aXbTFi9ACKkpFKYRDBm9vL8/VWdxzGpJnd9PHnW7N2kb9/PH
hYZYfMMp0WyHP7S9y9BUJZuWjlWtewvjcQgOcZim0bOCSRO+4VUR0EXzl1SkDs1lP69qQSGC8b4R
6JE4/qx+VfaChC4pc+/ySTkYvlWLJD/Clb3MJduE+oja90ZWAku4OsYN2yTaje8H0vh4Qe+2RtZF
3RD9C27o4PlxjTFJxCXkggLg/m/dvmt7UhFxSeNZze4T4PNSqUnzi6adMpTCxAHLjX8F7C8jvpgY
nm+TxsKIhHBZgVxRxhTJcjdwO36XUKrSAVeAtc1aPQkJbXzJNA11AUmuN3qfvADK9yRjr9FB+e5O
Scitf48P1YtheZWZDPKEUnJX77aLBwXGq/1Dr0dhP5JpcZP1jvwP/DK2lYcVVQvKYr0029+Kf4Dc
XpdsT6OKgsuB21065vjKg70FFFjB+8szpxPGR5hhYHYtZr9poz0je5+RCJj+Ib/THzjtYv++BndL
5h94Pd8z3sRThWyPZJUWLkpodDbtQrfMD5Yd79r/I6a/dUq3hJ5x5Kbw11OLVC8xdNIvQliVciQg
KyG0UtNoBS/1bLc7VH96wpIkgpu/qqSwHsVSFhcxe/5wiJUTYy0GTX9iZkSoEd6GISg7v78UJWYg
e6sYfzqtAi24qiN7dySy86jXlkLwwFUw2UtjX7LMt+ZtnxQQPCZIGeJNm/m3ImPzNwQmgAbMIEV4
fDTI45fBwc3/MqcH7yDXUVv9lEThCmsgicDqx5qfDqH5wiQrwuoDmVXc4JJEeROGZBSDQxZNJZbo
oYlBVlEKa/8xn2QS1UMFQ1NscXV57ZcAT0iQBFbwySiG3zOC+P29LIpWSMu5fmhBqEO+zVXIC8od
BcdDvOifz7sGcGa/J20eFia2ETnCsQSwaYG1DmBurtWVyyPgMoyOpYz0wTIlDAEM/M6DKV2s/NVA
wyDowdG5lKbiMAcnCKymL1CfJXc3pPP//7r0l7nwygpi2JRVWrd5KuEsVc3/DDbjmfYd52CxcUWB
QMj0H6qE4I8oZ9r4zVKR4tB1SQ1MZgljsYI9i2pPzlHxquxrEi6YN5CYWvt09+kJpH8FccvRCn25
O9ePgaTVN+RwBuJjNK58mHZjRQA7K5FSMTXAT2aVL1ma02cJCphXCH/rI0rgVTRvSTigUpS1IZgE
A+uV/DGs0R2loXtYhYZk8gO7Ytq5SKuwu47tZoOIpyPem92x8K8RoeV3hSMIP8KouvUs7BVcBbLZ
ycFa+HhAL810FCRHEdM8utp3sRdFDqHRFbKaJyFwI9B27ghwHVjlkQ/8qUT09ReTQKaMC4QlyVyG
6c69yw1bNWKyitTbB1hzzL3NLG5VPiijLfffzTcsSKamQVuqhINjIkKu4/ewXLwnya/SYnpIDqF2
XV7fD3iZmatSxJya1vpmRn8dIQKUak1B2HUBaWyDPuAoIw5RPhD4lZJ5J7OE/MG6TdeI8UKUQvm5
0JbHIWv60/x5P/JDX7bpGfmk069NUknCo63/VjsepMjpIrnYwf21RaaFwrM2Jpl2K7W657HvPGwS
DgYZjP3Z1r3/a0KIna5DyQSleuqnn1xXPG9swFTACGfR6lthKlOa8vF/EMtLYS6fTvrG8TkIrnEI
vzdajB3gsX1rvIbtPvUAofsPFy5yoW9FQwk2+MDVBtyVe5vC5nW9LALkzlqRioQ9n3O/fTlZJH/l
eLDpE8FuN7jLqk66R45yv6Fy3D+QRofFqPRe1wAEBiMze5njraw1vW2+z/M3Qz04XSR0KOoHWrYQ
LughhstJeMSLueaLCmiQ3LvKDE0Kis5PF/690Y9RLAexw8pn5XLj4R+PzPbSCf5YcqabDvRCQVs8
0BXVhA9HuJITyft3y0P8Jg1NhG5IZJjfmmW4Ek3MWaDCxi6uUruaGPz0yW5Z4PyHhcpM4CQHDzVY
w0v0An23TqSWny57auh2sSNGNp9CwTIXOs9jawe7seyCqxx4E9dotC9wcUOwXPHmwj7fdacUyy2p
An95SnHXObl18SPUj25nEogIgqufmzLJq7LtvYqppdykkzIuahZRDMlmiO+affoNJz8E3a6v6KQh
SymmTARuNYQbcFBKKUxg1DyfrotUFrfuzavT1cfpdRD/UkqUGAoNvce8AbZI17O6DoB2UWDNgaAT
fhtETGMB160eGlesOtla03fCi+q9emqkQKOKUuZwg8L4x+J+5/cbH9nJk1e4B2lyaY66xGYzbYYf
z7HzzmNOsPcu+9mx/01Qd5GvZYW7cw58eq8hZbu5ZCEXhsDtBIyY8LSO+FAHx3JCs1SGJ12RC69W
EOf1vTkR/quYHgZEOZvT+gcRJ92Qjg0nuzrwjhVgkc2HUhfYGNZD+kGtneqmOFLJvZVtjZ8D32z9
YSIR1rahtwefnUPRvDxOb21bNoJ6S/ESKApYKR8H7yWA91gBKrD5PEljtjpbpbhpHYLy7o0Ck9O/
EDiIm9LGgtBRwPLes89Dgwz+0OuDanc6V8armCa+IDPGB+4GeTCpX3rF45dxTCY6MF5T4MB7BxqC
v2hmuSkwWiAwRJINDzoCoTiwKyVSKSVS3n+yoq8N3cPR2iKf3RrGdN2/m0THJ9RhH1pJiXk3goBT
m5lvj4sgOcp9R6XUKv1p7YFi6L/a7SvL87r2UHOAVqhU9oY62UpWBnX8LRFI2AjRUhwmfzr3JAQt
mvEBxz3+AbO0+fSUbnbr6N1lY8HOW0rXsanme9kTIwwC1rajLUpi6i85jFGhFwXPMZUUPAakLnYL
ZSMQ66bJpaP0dg8bXKSamaafF8cLg+qY/6JFCjMWCPHJ/aypskzFssG2+XeH/4oLlZ9tCaeb6TTl
vXhsEZfcWz05+q28uuaT254kJ+h2YPuUEl9RDNDvoVpklzjo6h1W/mLTsdGaJmzvzAQYdzh2cMLy
Ld6ojsomcvyEYwf+m/tnaNIPZ+5RTETW+T7YE8cl7GLfP5bATP2+RgyJYD7a6tUsLZMxXaCZJmUb
5/US6W7IUmBAONmUYp0mMSnwoSaqX6qT/WWEKq63e3mZpMvVWK1dieLSNRlSffFd1D7MV0wU9ugc
DA8CuvfyI89HfwmVZAj0BioSuQ7UdIn7EG2j7DLBBaK5dDY+k4Hc+MTI2wcAKsIwPlVOaklz5NTU
irYBfx4gY+F5Y4CfQfAprnMEmH7xpb1y8W40PASmHDoqaioQpLCJ+70RgmeVLZoQECpgRtM0BjbP
tmzU8XxUXQa9KxlQnzEprnkJwu4PWQLaNLE/CO8guqIF6lPvI5W21a6TrppjdyxNkxhnpda6Af7U
Pgxl+Uhjx/fdtEAiSrk/AprexzVCTmkW/2VPDNvg9xqAOhIwEUK71HXLvNgtP3Q54DvOyFfNQzPQ
Z/DzOeTLg5iBlCQlrYO6tZCCp/uk7xBzglbD06YY7RR02AN2NCQfq3A4SMDV+2A2LPG91KbQYIDZ
CvaMArCuO8pZzGk19MY8pDTFwILSYe8HDNw2MnntFddtWsKrztVZOIY3XIAAEvBY882G/8o918F5
uOD2l0RotH6W7b0Im1UvIfHBBT9xHgHAckTTnWB8vJECBaq7HRfJuhAONd0llIbNth3yQT0MAhln
nSHTSeCbY9PUsYtRhxC4paBgJuOkaS+CGxZJfHq3TDe+XbsKWJbJ0Z+vAqXZWRSGahmuqZOvXMA+
pK8yhwhOtTSmUyaTrgcZhb4tYTUJrnEbVOdOL/2jK89fQp2Y8RBI8mjMioU4NoVsiByoxWKh726w
BHmJFwUzvF4xQJ0ICiEaQha3DYIShvqWSTmXtm1QbxyfJxbht9p36mc6PZguxaMbcuIeBlRzJtar
Cn+9YqJC/6JUcV97+U8BX/IQtvoS/jiFTa3uqnsi2rWO+8OeW6XRDlArcNcp5gNv3IdjGZDPw/23
WG/EAB32FMGDHTkJiuqdw6782wLBgd0wcNJNfOSXTzGxO6CkIepnbDazIhm/4U0M4ap44Nx4zTTE
XjwjKceSTtem9Wym5sV/Ht81vNuT73GS8s1nC3flBdLvkCG/2+B7SGlBGyOW6n24+7GpVapHyPXq
JG1fSVNrisT5IzBMneYg5iApUyM40IqQWoWsBR+4y9OAKboRlywVef3LxGka/qmIzXMY3VKQYaq2
0JmgJeWu9ODaAhfD03vFIIhOjIGpgs1lMbrN6KQ5vBcpR2qSPUxv+dh+Acbb10LqOELIRNYQE7/9
c8Dt+0i/sNwNm1pdW6Dum5mepK1CAEKkDHE3rW84kyVKYBjcTFWBFvNcnQT0IqszrhwQMKUzD9xy
n20Xdo2siJa2ZhqWgWoTqz/9KL6t+PSq9jKbnqopMeVIsBgZbbDayYOY0qtFpcYsmeESyT2FL7+Y
CKT2jpi26qR2dbroVu+/Nvo8RVd7JSzBIx5I60lIVchXJzU8aEtOGoUH8EGVM6mNP30JQbGEid4O
XBJdM8i9bkJ2C5Vy83LUEb4SLx30f4HXVR7zIhujSqOaLfQ8ujLoLEVrcHqJYcrNYJBCnzP4ZanF
DJ2Z3m4kd3Ym7VwC0Mv5Qjr3qBRred9a46QB4XufobcIpvaW2Xgoq9c1KT+EBItyTfcQ35fncXQx
gHwwMtH7/jIDo4fw1Ff2sEflgy3+dpri2K+2QCL1FElnLhyCzDX6HdjCB7wFOq8qBKw/ZfLrdCfM
VR6u+LFmLHGF4+jJldF3patwJYFi08rmaJci28slTcdV1k6FLxL0yameGMb8bUhjOY4Ub/gyyWWA
vlVx4nTNb+qleRpBpczgfiCB2b56hbdLZiqXqVINU+l8A9XWQkMS9tKUdsFXjlJTObsEWaleEgzP
qMZZTNEjRVCwy6RhcRiQXslSXDrJpRrOMkQLvh0caYixUMS/vixrBvZ8pSMFw0nhJ+YcwZAuBeVW
sRqBXsNHfz5+O+KcXsUXufidO1Sck36J07CK97gC3m0SWpuqpMv1bVMfapFdDxJUNKQyNCIc+kmz
MWp2LufB44oCfpH/YaL0r7Vl7dz5BwjZdYAJu6DXS0GtD4K/F3E+gzmXnMPuAJVSPhrCSJAdIpsr
ut7g9tj8dDn+E9oV2Q4g31kw3z2QBUD9J1lfDt3SAIG2o6MBg5H2jAwDsCUrxWvnWDpnBsZgEyOD
b/FEfWoWEw5ioLHG3KT5LSR1iZiGpPyxtFHyDUATekfSPb3vEASM+zfGX0XmvUfd0spYDmJ1SBnh
J9fqs7LEXJ1GWGIDy2VOS8J0Ml+1ws2LkZSXlUzsvQLuIxBgQdOe2A2zcqNJgdYiEKc5T8HOgIEE
Ur58HhRt1X0Ijd00JuYeFnxUQN4F9I8Vjgz2WLnba5NZ7AKKHQN/hLiSP+vsZbaJEwMSK9XrVPXJ
Gb+UhzM8rP69F7MZzlreLw+sTnu0CZSmSyivLotCoyHeMRPEngq80fYGzpWDpu+reFicap7ZZQmx
st1tlC22//r4hDg1H0a/TjDF0A2v4/DQyNf9HdvvPnlRjzCO1uUXQxO4QGqhXZV6tFwiEWJhZM7X
fsQ1tws4lr7j3qdoSdIFGIOn7eWNPqaJuHcr679UfU4SA/N9xKQzUVckA1nSrsRuHjQYxm/7eGpZ
xt3kU+hPl+ItF2CRQmM0wApt/s6QyoKPpUz9hqVl+puH+zPcKmZ3ekngDerLzhqL+j24BKzDBVtA
9DND6YmjFyoAHh861r9n/HQmdWHeLS65Aeji7e9D6t1poxr/aDD01O3XMtFAs6f9Hv60dsLKa1zy
E76lQ+ezmpJZJC5TAvnC3FPZxpHsU3RZZfRG9CnARvIytZUGpe1ZixzDSB2QKIN0Kwg5psGnLHM1
Ngg3HhEV+Zgf5OzRCiIniXigIsGMKVMAnP6yurmXjBXcSMIbMR3irISl4yMEJYkXGfHGHJ0b/uvy
Pi+1W2uOL5PZU3dxWYEg35OtVSH3rE38lddzTouyqciwM94GuAvCr8BU9SJzhQOvRVocTLhn5kE4
pSd440lUfG7vc5MxYdPAkf9+VCRK/41rdRySpuIwYbunl8VVGrWMrZcmaZ143R1/6tcC+zNh8QXk
EcM0ermb5Lm8shX/qIIZlupZcOgSisVS5SV2pQ/i/TQio6Z836JUo85WEmVJcLbKiw6qZw3EwVN1
UB2mu7PN0cRmo6PCMT0RCiAxb4WVHG+Nr+s347lKRWXKADMQ1FXTKs+XEjA91iyr96KLc9jkJRlT
RtLCqq0tHTIm3qigxCdrjy8h/WR7ccOlnqn47qtRl0HM7jzIdFlkstnybjKF7Ztv+EMb/tecVKpb
f8TGL/8aNtP5BxNe/0YoMdir3FGpyIgQecKeJhQYoO/tppgSOG0AJGbNpd43zVAqWunrd5OuZN4u
hKRXhIPLftb7XWrQTKfG23KA8Jlp2eXm+F+0MV2/fdcmt7+jlE85HQuDZrd4Tbmt33uAv+Bs0ghI
0s3XGEmo2qEIkkx7sCLmFzUwcBSJFWVL9LVFnmlKug2LePEZAwqJO6LvxFcUSUTuU78DnitWtNrM
KLJ92vKFk98jaYGe+GmwN1/IssK6MH4ALtfgyGPxzcTPnZGQ/d2kDifwJVlKlmUa4frTH0d7geXy
Y/G/KJ2lcgjlAI3hfcCzqJEpAux8cpl59U5g0zMczPlx8KsNf0X+Rw7iSLHTh2svLzoQFw/5Zrfy
bw+hnlwSFth/2K2GoHih5Hw4hiJlCHAfa3C23SLwG7Ml8PgypOlKK5wODLdLvSmNI2Tnon9AWMw2
4/9eZZb3oM10Vn/WIv9HlUwjYBJuJAbsDI/c3+bFshP6KImQVgB+2FsDEW5lP/x14fH3iVOhLuS2
EPT7eQ+0wA2TK+8sqfm+T4twFZ/FJ1YWKwxMwPIdLKeWDCInYKEuBjzQVbnGDLHzdwN8Su7lNrhl
kFbDtMpDatmrUs6aPP/1pPl4NcRXs8ru4RY1VpCE8j0CKilN4XkC+FwbPAXroJq5m8usQORoLoBf
VaDbFPZ82isucz/fwBBVxl0HCK7IDLPc3Exqop6+ZmfcaugakJpyWpjbj1ExVBozzLJMSq3/VAkv
B8K4c/3pbdnnRJ4/e1a1BWVVJ4j91jnO87reYkptum0noTmk1W0mlSOoP3hX87CYMhrk/lrT+mB0
HLb3J1fY7AaYdAas/Y9N18wzd4CFIsz6NUlJFA4Mpn9TmjJwAcOreGkQaFbFdp2iXA1gAvGZTG2K
5ZKhbKBeIifYAK9nWtc2vCIHU7pgptZHntb1T1Hiw9I/kHCmDaPzxPuyHoN+1ImqyN8gUlkxfe6s
gueYRCmRRkfLwk9XbTDkRlLUXZruZsyObql8bngp+J7CgXTy/npDs80hR18M46dmSxmNazLj3xlT
MNd2t/RLqzoLKxvAJWn3ymvvgQEi8zVzMA/hMbh8HTWNt2VFvnduwek2C+0uQ8FNef/WU45Rb9e0
IwdYhAH4HcydJG9vGJHqP+NSX0J+KF1dNlk0uxJS4suZypRcX6j/hmqqT3KNq/b2xj5uc8GQ7mS3
Uu93+iJliNkr1kHmQeaLl1sQCf2al1kCBoxB65HX1+bvxAzwMx6lOSpoMWK5MsDf6cdBfJleMF57
YpsabjdFd6GpXCFVG7ajrgUbzeEdMfFyduJKMXql8rpAyrrQkS6BnmYrrUwS9b0cAQKWMhVAu7+/
/HGEncQPD81BZNzlgZuVYQr4mWgsFx8lgrPNUsXboAKKyR76D1sEFd5mdnX69sp+zw4Lp/In58wb
v7EFIjyVmD/J6/cYnD1c2nQNzQ4+ix0DwypQQTQmBe62No9w9xh1KyuyE25ndvJE4Q9xBsqyDFsC
CRfGPW5Qc9HIxM6KDJR2Icx3smM6nS34QAY+xwHnCKQY1xvYdoh4r3Lz5oleZ2K0yzvuZdNzi3ZI
+aabgwdxgMR1U+XdcDeihEH5FDI5NFpeGMulA+2jMfNErVEDuNa2A6VnkhBWlD45FVx4uOf8SHwn
AqQoN5I3wpiBD+Un6a4ZZF3lSyGTgP+pCTtN5CsE6Yn18MLmEx4N5wwabei24fgEgpw1HIXTB9HQ
lxfLuFhGrxE5lJfgs9Fl/aoouZaVirtSGW0918i/5DgS7GPVHZQOObQDwyr4WlIcDvKkRYEGduVp
op2LtSflzpJebivhHUVfTmfSsuy3kH55NqMBBMwbGL+6vlcMeCEpWMsD60p+T2SZXkWMsNF3RlQY
cq1grIW6UWRuj2KbQD6VSLSON/ULZHsWrFrkpLaSeTRmRw0Vn9jOs7ZBr/u9BLQJGR7fQyI9kiV9
bLcKcOB7iz5GZFic3tOq0/lGsncmmlUYP6GVPisur45UW98ZYapk+jc7qgPNt/nBFYwKi2NIkAnq
Wv51aGEH51rrYJKaBOvPL2O2Vlmv1CffIDC9Hh5gXxldFBdvRLnEey7ybwXj+/wn5MEjZzkhrc71
Kg4fFQQ28UZp1E+3tPeXPYItIl46W+sFv0x9GHMGGLaiuccv66PIlYItSKphs1/S0K7kZd40Eiui
hUbPqvYMXdbTPpfoWIcgY0riPZaaPW87Md62nN+rsi+VvgoqKsiYGltaiwJfVDgZlc6OqZJLtXlh
EXO5X/+cAQpzlP7iHVVXUcklCkr00B7e4vLCTrLwfBx5t9ZJtyo0GDVTTF+J74coYvrgwPq/Yiar
T7Gonqyvai/NlTw59xYx2iLsVpBmx0YNcTWx7TkKZrIoUDrml85hGDC4vALdWEhYV5xgxtq6s3rn
X/8XkiuBeZ9hlaU2wKelWjq2PYKVb2QGPOel3QOCmT8961y1RwRBaGw8GmUEaryLI4/8dbz44Fpn
5PWov/7gjPaEe48O6qxcX0dITmeGo5DOGmanTUuatbWyrxzOLPnzhHY0PbREpvWs0b/hdjtecqeZ
zN8/c6rEtlk9zh845ppQkWcxjpLgwhqZPyHPUgTHfmpnvuCAI+ck3YNMth3NnwIQL8xp/8TN8RF2
J6U5k1r8OG1aS1g1NtND3ZuuREUFJEYqnFnKlbBn0/xnvQ6Le4aPliVD023POLXDlkfgZmNOqV7H
6AjAfYzY7uBFDAxMNek1ke7nS5ZnWLdf4Reqye5s8uw6aIEbm8/Su1++OLCVhc+hE2K9s41BOpCJ
/Yvbh0kh82IdbVk8jExyE2lEia5p4fy2qqyKbZjMt8nyQzqUpviGzctomu/y6u9Ve1InhJRVyq+3
mWgPHrDBTSOuwNVRm23+/3nuadry2E1TWiyPyMuPSBp8yX80yAmd5rIILIUAnwvD/skbkh8uTApq
p06+HEb9uYeCYWuUr+Ch4lob9ju3DhThV1UAqbmHGzGu+hpeUvrNhQLxdKuiCdmbZg8JXoT3EWTK
8+84J5MnfBxuO30yH6eCFBCTkNlfBAi5HGg8CPIQtuFOwMY+3/Jh7hRMd6B95aXZm6Dej975D2Rj
Cdlrxh2JnDRw4hSBld/6FVp6MgTYcEIh5ST1dZRhKFh0QnFyh867qypeXjQeBKH5tq6TiclZZsFC
L+yZaGvEG+sJgt6tWpQ3xV9FGgs5gIT0d4ke3auk4O4y0lU/fJI1cG3bFae81HoP15XvBEMXMK7H
NQna7d8sT6DzBMaYhyZmJZ38G5cmpgBPyVFXLIHfIS3fN24AqvVE8ntSkg8P4D0gXAy/KyZFW2Qh
49M7cAHDJSrdAyt1QDM6dz/+SNjT3+ENU5iGqwbeIdIaOvV9bK25hEVxl6teh7jT4fSIrTpZ1Bss
8RXQLGuSFKua/Rt+EuogScivjJaYn2XbPNUV5qmNbUaeBihA/NA2lo7JriQfnVXA1lN/whDwgDXv
4apdkAvd7/iIaQWr6fp73pLTvxd35TveOg2YA1SeAbQ7OpRirLrmzfznrOnle4ReOKNQaE90ojhe
gcTTpiXcIvyYvrYOvC59xM1N5kthROocGlgZ7RLCMcHmtVpm2/tEnA9wz4i/sAsHxKlVC9W0Km3s
aqVfc+XheVjKhLgBjb+wuM9H5NVKGtdXiDO9QsFW3awvBLgJ7TBS5CFAFpchi/CVOaSnNnOOkqX4
QTFErq/zWBKfs+H3O3O8SV6uYrB7q1mC4DSiSVtiajUwr9zhAKzPix7NpbA7swUjWXmm8nR+suJJ
caAxuIPTcB4LkuEi0vjEkQBmbWyLhYtXY1PrqIq/1TJ2RZ3ao/rsulX7ZsFcLeNY97Tfzy61j2ps
BhqYHB8YqrJpvrXbsbUfjNWsFjbUNbjEFULdBleu9EAr4v3UFDG4mjhstQoBE8b/nGiQ8caOFJAM
gjPzbco1+WfDn5gsgEUhs6iKTiZXy3NwyH6qU/33E/QBYDAh5Xfw1WN1hnSLQxEo4FDRnXwS50zs
f36uxojbcLwpaEcxZqPQJVl90DSIY+2Nsj9MuPaLJ1WfpbzES7s8bONzxvZIOlHJThdaOfgIyrzk
wPcrIhQRER1TIL1wnC6I98lreuvyd9g2F1SDwKg+tdvH8w0eoCzbRO0ssN1tRao/CI66FGdCiguE
azq2fSHEVOoxPZetr1gXLdL7cu8ZtTR4FVAMNGXXUhWycoSqe+3XMuO+BTqHHgShzTO/TNvV9fQj
ZpIki5EyzSpCFNetaKvpENFo+gf5Y+//TbkejQy5Mei1S+CV+9FloOeyE8lSn9jpKg+D8Q8fox9L
FFC1ZpAZXZn5NfFwrME6Z3+wvghQB0V9fMsx4zDsWKkZDLPMBk1rQXOf4I1ygHmNNhho9VCOFNTs
QWgv4SVIgCLFV5JBELabvWw7BLTfL2rLfjG5TKBDnluqm6MmBd4EG1CKU7eUJvDKL0GW3RwptHEO
vV7rPWQsM6e6vAiYkw2bBNuiuicYe6xcEStSd/zCOKWX2LcHoP0UWLJjTcUWyGiIRqf1sh/+vUUI
N1R13EHNmDId0XDKGBv/X+qgVI8XWME2uM3+Q44Spk3ZYeqJCukYafd08kK3en4BLu3QyccFT8oq
TTeRISa4pi+Pf2l56+74pm8fFvAlwQvUzGYCwVkiXgK7Y2eLl1832R5CFzCxQBPT+6LZbePili3/
CCUkAVqnzUVCQjZ6eFKruruCwwCTLev94qVM6TC7EKmXmuZQLvwHAEGUhA4yzB8OgPLVG6mB1lNT
7XmRoP5fgJGy6orLIz4RZwU0BKkWms2qRX8l8yCgVbwOqvYVVUWfvhfM7IFlL/KBLhYjwY0+pRH6
xRiMXyZZ4IPLZCLYZR4tGfZd0pY3H43iWfA4hlpXLev24LswYx2zyvlJ1hRsDm1nxuzYaqvIQoL4
ixsvmYV724L+RgdG0idlVSVHOVWLsUEe4jMbXmj8RsGhkjoO06QNp2IknZZkxWbXRxJG7Aiid5l7
R14kwrFqpYPX1BMrI+/v5I2pnTNxIUApv56HUzJZydNpa3SSn+Hz2qEt5iA9XJoUAKrRJTrsSLzN
FDcm85ozPK8y/nPPSjV2jPja04DYCFEC956JIGbB368Fdn8YVBNLHOkD1ffVnCfgX/UsCYigvHC4
LHOXHbOhbXC9NIauFn0Yu1YaRoeCuIomBIhWc4nAxIVWBc2AeYgVMkyYlq8rf2NZNYYg3CxDfvoW
0zjda7ug2tWTKylKGHRc2YhOi/3XfAwLBtOKJr8N1MmRujD/nVry0KBArdyx/UzK1Xd2q5JqCLhZ
7ePIJKVxw4VlmcP8QNMiZM+Z9PrrdOIhpwrYTQA70+D47eeVPUkXB/ImJ1IidNVvpvumFb76/bo/
3VNCSnQPLZSTmYi2Y0/7cByfqF+/FnhpkveAzJizoWEGQCiY4OXGLbif1DUNa07bZJ/axwu0iwB6
cDg4lyOFgVt5pBE/zwhgXwoACiQoDx22S52lCSU1EZr2Ef4pI0CUvXi+dcOUINqg9UVzYNgwOkvC
YxSk2L3quczZbYKzkHOypGPlnFPFVTY9TsSEM9D/HWeSSRUw0Vb/sAlov4ZgHZ4ftzctKRY89gJw
QT3+MjEd3QZBa1XLp67aT9wuzIi8XuOOGARJzBfsy01/0oZBeQMSs3/tTi2NcjOYiuCSYrYtMasB
qi8gRDeejaEVi5GUiF1v6/XJM/zA7/lxE+5RcgXtjg4Azx5lKMwvdzxhthnEltXZbTVtcRDhm4wG
0hD2CzVqmufGtn7omJ3N0zRrcJAQvnlpLMYyMo+WVHZxeUYRRSdq6hoJgZ7UHwLBKUJHdFEsahgc
fkcpAps8bsDq+bNN8wIZwTxX8O9otb/vhfTVh2iJqsAiFFG3IbFMvsgxBu+nI2DKSEuVDfIgtiCz
RIBKxXc1WFp/W0cj+Q5MI3mzc3v1scY3hKl66Q9tEW3L0qffQStFvCAQvlW9DxMX0KABVHgjLiXQ
H+IgrbgLZDRStOZbEzh5rUR7CdhI4l0Icn2KBkCU3Kqcbb4J9YJfwFNmMJZLXsJDcW2cSZi24t9u
FfBSF1zptN6JrBUSeZoRqBAD1k+qMHb724Jy/bs3i4UtaumQf5pP7DEFGchIHAB3C1ylPlxNPWAA
CKkZs4GWdYcpevmqkK2Jujwl60N2C5An+W0X9gEhKV2WrJp60oF2lqc+5+zs9YePBr/9iqHYWOCv
SAgY59/LnkLp2rqCfAu0yt8R9TH9hdc+BZtKT/8Pu7+KE3ulI1WCq62l3mOBeT2RcEBEVeQNnYYE
cmtisg0e+7Cl6CEImWpPMOPDySYI9W2KwCvgV9MlSq/56X8K3EpB5Kj9Y6pEhka+Yy1670CRM+aE
xH2BlTJQJPOXSQfaRo1GuOzSsdMYEZ6D/f8od45FUAKBSzFs5ofAri6V+iLcKZbjFWRtZIV0jBi2
eWFXGNx1e6BDyohNbfjIzvMizohen1QjGLf1OS7lLzBO7DIHXg0vaZllkTg6g86P4HZQMKxB4pbN
4rbn8b6mFYT4T7sySTLCDKtIG/X+9zMuaBKYmD3uVZoLedT2LUUyS/gnfQiPdY6dwEk/q7McUuWu
WkCDRVfX2HjjTay5S3CFMm/p2AiGdzIMveg/0UuM5UDb83o7jqv0mp7N80EzahV16iUHcnhCImff
95juJ+zRrxgR6NuiHWvYXfjrrIzLocsEYOllkFhzi/wAKzunKoAtKXFb7JS1P4ZzU1pLzg4cxdVS
hlnGSFoHWmleEhFRqqqJ03Vb5bxT9miIL/+kY0w6GBGZv2djoSK8cWkQ6KyGbXmJ1UYcgjWSpTFZ
H4tWh/o+c9y+7+2S06SyyPUq8mHvGghS2/qXt7mx0SJKLBAG/Gzt4bcLvebEqMRbrGOWrBoy6+pJ
5x1Q1NqKbrIZxm16aRVqqBe8zRido7KVlo/bTOvW8NcagHSHd7NK0XYOjDNwG8A8FqlBoO4koiDc
dXQIDXibGN1wlXqr9EwEP7h5Kj+1fHr8TJcSYxJs3F+KTS/yk/3uX3LSeYvQL9me7ayEmbskT6Ur
FKtYNmf+3PSViGWWIwEl3kVTHc/uDgEMxbDESLy2P9MPC8fxXTy0eUMrJktNEemTU//5J8S5yM5Y
DGHL/PGAFB1wRPNC/IE2t/gFOaPc+ywlMg6ArC6eTUfCYedDLYh9BOSExalgjdXcHf0/ud+2FBoQ
oDtq5mxnkK7bGqqnMlpTRHfnEBHaN0HOuA+1lTBq9jVrj19MXRNBTXC1Hpa1Ge/CTLJlf2MAkp2b
BZKIMjAjLpc5BFdp5uI/wzByT3EYn+ZxOXy7njTJ4t8AOLwU8+FGVF3pCx7kDOACOpD3TaPTfxBV
DSrW8H+bK0bDO9skJ5R9pubDeLRb4BW8XYxMny1+ysFv9exrBZXww3VSVb4egrzv1Mdt6iNCKRJ8
PQRLWuhZZa/LV+xDBwHOFcb7+z5Oe91h6gl3ggCmTSTj1CPYOP9bSwpGKX6bgmQ87h11yajczx71
9axPmlV2lt9RjpB4S4zam3qtVm9YYfKbSb0toS2N9Jj5HgV+tNqw+2p5evNZjJNxZM4uC45+J4mC
jyNgptMsxjGut/GXLdohrv/ykmKiNL18CkhCqeHyZekgTbjpTsXb95lDHK61M9DNIbnjPQu7/k3J
sJpcrN8WNWN37XWZvKAuhTjDgIb7iPmXzMl7ef8MkwHWPuTq5AwFQu5nUt2rZJWVTsmFfvOBiHnw
eZcMmBvXFrQUW6xhRfsZmfLQCJGJdVv7TIslrXvv07pc7+Q/ybzSESfu4DeyaX+tsWBwVDi7zaES
v7dQrdWnrb3XRn5Jas10Frspzh+2qJfFpd3doGsUt10cD3fJHx/Ju9mx/8VNo0MVVPj77s4WbzE+
qbxK8nSCC70msimjFqVV1bcaoK5kwxdQu68pfYoOGv7WvE9ZOHY3iEBisgBpL1JCh0sV+WJklM73
bIHqVygpnoYBo+rWwVMFp1OLkKgwa7N99iYgp6qhK00ZznItm0GjL6bRE7NOhmiQ3iEIu7fGXu+x
hFF2mM5SujTwRPmP+GNDi8W6ZseFfeDkpMdviSOps7GyLDRQmQ/nYw04QjswanIQdnodABYZYXDa
cnu3TLhJMFgAxVIIa+oeGpE5SFcm9siVisjJQRYHimXryyBXcwlpIBmhlovhTPXpOKfC9Tu0DQ7q
ZY82T8TKY2YK+eGWTXfN3DBrE+Br4bM1SQx1ry2kHjExnojflBVTxqxT+fuNd8YkzDKL4TA75lcI
A1jrFkQBixEZVpnt1DggPVMptyzU2k1LdxvXlSzM60kaSyWKBph3+SlpOvKU4dO2j+xuIxWcV83A
fijxkFWDJSBuIoLxAHcVsNbkn5dkKxNs8ByJMWEZi969CSdBoBNEopJEOU2dQYazGsFxneEyvWAS
LNmS6VeVuAROZtaS02hY811ZMVeBnwYOmzrlhVC2TGMPDaYimCnPx2R4cYgqmmJZvvsSbKAJldwQ
IZShAFj/fcFO6IZ+/RPtY0Pj05l157S+nKFHDRAwsf3avtzt8eNrVjBXQWc85xTnp5j4o/cQiMCc
wshusejjXmmcmJh87Vfho2/4nQ1aZesRFx30LpfpnErxM1cQdqAH+V41AdCp3bajXAzWZcQb+mjJ
s6AYOENq8OOVj1f3emoQIKk5QohChma+kI5F21mWCNxinJbXhS/XSQqJkzbmuXHYlh7/kaKNOLFb
1YmP7U0vlkYNObAcHZzaaWqRTTuxPT2N1tqZW6Jyzjbq1xTE8SPEHMQLDMFlg1ZBQFnc0xWpWKDm
oT4iUYNu3WyNUctnFjE8gPIm4PXeW6OBJbPL1txtC9FlgyJ/5P644zpKafkZGuQMW5ATMW8vEm6K
0ILFbOQ9pq4E69uTelOA1qEPgaKR8bV7Fzx8LPFQ15PAwZSr1PI7mp7ER1NLep325da2s/+AlaoR
aJ4qHP+/+4xUwLFDhAwtzUMd8rOSJw1wqJzvgkPe/rbZDB+bC3cPCHUCjQa1ibg9QyOCPWz/zeqb
kvr/dj0utdaw3MCJj9qZo/wuU8N5Ed6RWUJj0wN7nTEE8fmV7B/VGY2JfbOKPos54LaILFlC0No7
ESIBY8QHoxFJLXZOcRsTf8fE3ba7t/2VHQHLddIfymRnYyGEfZ/aXNRkzka15riXhjGPj6XCC2EB
czhVqLumIraP2rXTTJ8EyNpOARzm6DMT2iVBv/x6k6L/GnVAccx01YoYIo914U/Ukb/I/jLsR4Tr
gKertyCrU3zNuWBMGPgkdJtwaxzNdmOcSF9mN4ACVhDWXCwHqFppyioUYtlZ+GpnIlVjmVwBJWoG
zzmrYO0+qP2t459hoNanhekBBNkvqNLWoVSwxX14JVKwI4E5yhIJpcikpnTFFUTn0phERPlZAsov
7UbfgWpA0I4eHfBLmpFQ8YJqmUdRYcXI6mshBSpFUmekQsAI1iegG8fH6ilO0H6SJ21EgygFiJnb
s3C3FFEM9rvhuUg+sDDcVnBs6hoOIyigztSupXnQuKVoQ/Cz6gZK7rxXhLfdowZ/SzmhyWtFmQD9
ycoSaVI0h2bmQsYqac+z1Suq+UY5moXdu4hglly2DRv2cM76EsDIcDC6Wu98rdLo5Hnde5sQQIHm
sJBJThxa5HrOhd2tK+gXDkBfeKs0tXIUsRI062Ni4ljP8Mjkzw0y00aQLER3T7Gb3/ub7PNym8Et
O9B51BNWe6lPUj5X0UFW7XgutV3erhi7TbdTyVVPO474hkWlEyXsQufIpXwHpQyt+pG0Gt5VvIjj
dDg6oerpmuY3gdlK2KEn/IxHffxqpcP4jans/5/hXW7GfTvmzqi0iSy8ULA5pVUXl9kdgL0+/eds
sU2duA4PZy157RpfWtPtEt4QRrl2GYvQiqVaTEuE4Dwb0dqGn6lvayAoM+QLtpQXGBDgjIb6YTK4
i0/jOqKJBJ5dmCpzi6gK32sYZT04DTVG7kjYNP2ws8JeRKBQt2rT4OTPf1T82VddN2unbWAJesLe
hWNj2vBxKQoit9B/FxhEmGKHIW4WlwAaPo7+7obaziPafo4BtHUVYku8ZSLpRJk8ynjeOQCuhzNU
pGsQcjGU402wpywKnOUR4E2w20GCR4g6xfCMoaR/DMkWBg1rUJW9El643ADBX94Y9H5H3hcmbPE0
1F+cBerN9uN6DOm08tgY7xk1pSSANFNKRHfxFm9FOzjeaVA/1jUgCf4ukSF7q6GbVukd+dBkkV9n
oorW3t4lhp20Y6WrasUXB2sXXBMfvsXypEtEsOVfvk21+dZX2Vvk3f28KC7ENAVvMLFQPF0Pmd8O
oS2x30QeiRYrBu/e37x6TrkwuLzzL+9yS7M6soMkTEufx77mDS4ElV/0lGrJa88wTFL8Nt+8cLcX
tMU04j30NrcTiT0NL9cvcOgLzJ/Pz/7q+s+eUIgnmCIGjzDDGrxjre+ZjIqi/E7mMNpQuSNdK87I
8Kia81QFSkRmUZxN98hVttSG72F78Gz5PTA4y1/m5ceSyp8gQTzjrlrMi3n/nNVoc5VwVNqolrW0
F8gxkQoyDTUDTV6CnwJIQs+BZ0wUrtM2zlmFJXEBKAygqAuMa3KbV982l+2IKxPIbeOPc8iEjwaL
7YJoRM6ENBhFvzgvo2euHzPZLx2SZMLauGQkk+9J0wFzUvbj9PpeSr86iexmdhaIr5sHvuRv9TXA
HsdFwIlGlmP/yVfWRT4c4Nl3M7my+eyzI3IHhZjJwichqmXaCUhTksT6/r7Wa4okLPq+Lx4rD7jC
e7KMVkbS5eq/S43aUDe+2/Sjs5F+NqX2jUksuJ4Dx7BeD9oJiFF66fC+479Wph7HvrHyZ1sWxdKA
j6I7lp8rfD1xC7FiMbBX2rFbDLIqjJtJr7XJr20aTxlM+hkZpo0yiehNnl+LWWNtNXb1+c0fqiBu
X+woLG/GBEbptJ+FaLSrtYnNGgEXXY/nvOnFV68gFM8nUFedoMgrJyBJzC8s2HgbFd63yoBrSfGO
x7IYOls0gYzsbAqSwG41vwyN3norCNJZiS+wTxHApYGURD3J/wZ+iUlXOWBQ5LB/kBDky3kj6iar
NyIJlashmFYzkI9EnJuFlpf/P8CyYqEBEaxG4DOeNa0od8o8A6qeOXSHFg16bjaUVDOpYrfNQx2x
ol7UUmPAi+9N0eWuZFw6sPv7bruPpdDnrLmTSBMWAbqbLTw1x6kOSip0+59Epp0l00B4fwn2PSr2
ouWrr7Ql735HnbUZPRdvJ5zfSgEMVXKZUH3nYnKYmQCJZ1GsJrKPOEhKtt383WucElLf0iOLTRb8
CNzsy4lpj3zf4ZFNH1RpbFaNnEkTXjbhqB2SSJlnSjzMOgRYe5PBTt3OvHJVH0LbhKA6UZzhff6z
VzZ4HBsNJeNyhOvG5pe1yhRAW+W/CQU2jyyBR/ouORIB5FVkNFrb3NQbe2IymBtg1Y6DTPQCSf63
0eSMTeSvEx4Ief4PBO1bbNiC/pYFTzJNX4tLshNYgmrnaP/YNwxQTTTwXxZfF3TJpwkoJGHfxt5p
Y+idhQW1KtILmVygRu9rTOAISxsN28KImo4OCPYO8zN1VB1s/1HpcX/ON3lH/68sCAX6/pwAlY6f
Pb79yVxPhNpbk868j0TSw61NkREzHitfd9xAOEmnz+Ru3E9VHUeY9+H/+QKh+Y8XnKurjiy27tBK
9fIwPwGiGlmstn9aYqiBrTaC2volA52y5kZPScLD10FmDOY8jgDkZFzQaCEC8MNCCF6rNfxdHJ4C
gV0sXsANbMNTJrO8TOlQ+tHMcEZXFZyRKkpvSQklSGJ1rjKvxrBwyI8LKE25JacJXHdGh4h0sWQ1
WRsUPNRrbh0RdUhd2Amsp6IFhJ/a5OxN5D67EfjtixwJ2Z60OCjMh+wot+jhBH/uv2XY0G91r/Uj
MX4KsxKVCzDr0zTa6aa0CDkI9lmzY+ysUkqWPmJOp+d7ozT2l6XTkVy0qUD336+ANI4xtf1/fVXh
4sHOS6ioBiDurd2iQNgbe1v4S3fyKU5izgPkO2+DgU+CU6R5U+tGq9VrzbncPSIEP5GC06A1762P
MZYgn9LyO45CfJ4thYywA6z7XAlJfEXJHfrddZ5WpXjF5thNt3ufKlWdPGcflmEL4pc2EeOORvDK
z5Njh4nGW2GtOemWxbviKkF5b4k32G9BAhPe72fucMtISroNQDih8sw+aNLLX3QJQJIonom+xVji
tNroBfG7XQjfog+f5lGdKkheLWaJBxqlZWDjLrdahEwKN0TdozBp12/sks2xXbILsawV/J7xUvQV
bgrm95TwApw1WyqsJD9n4Cs7eQl0iqXuNOLcsvq/tEAW5n292EoHIDad7EIdAvRaI2LF+3lucfvy
EuA0j2aNhupp94qJUXwTAzkAwNE6uCnVnWdkvUk/Y9hl8pazAj8jc9wAjzGpqcyW+/HQ+7DKKaEa
8XpJCA5a3kDFNPHeDdWY33nzIltSCs0+QuwYDjvmzYj77yWCgcloRwUe6+6NmS59dUDp0JszxvDX
pXmwUWvOzSRC9jV49L3r4Bez5p4E4/Ft6ENJwXQO7FtOMRoBbKLsFONgwOIDGbf4ZJaZBbUNdJ2S
cfsU8pFhjGZ/kR3eqosCh971ft/GlbQBVc2zql+UFvIPyxunN97BZ077EyQEe0upOl5OyBlxc45s
Qr5kwNUaQ0XP2tQduj4z2kY9IV+gVdzamYPmKyibLD0rt/SN3KDssPS+w5n7lw5Nx5kYGqtHq/RD
U9fmd01rENqT1LbzJSN5KigdundkpxH9hISUJ+Vbu5Ztibf/V3yF485/oadhXtLt2GzBVj8cGLeq
bkbEEmYgK2JBxTiE17JO9rljFHHldZl1Eff/wPYT5wJGlZOaPx3jSkomE4u0+SsJnXdaVDi+8bpP
pRsZqKrkSqRPFLZIUqpoMqWXmSnr8lTya+xPifRb6uYuEWPvI8QlzPsXFHwI1yj7zoXdCaqGDJUN
k4zJNZut6L+evWM4/sjRmLwcgnx9iyQoO5Qb/F8A5xDrWns0MLe9geioedJJ2+ngdf1xZOE+oOE8
veKGtQ9of6uvgaFD/Xt0JZgbwd/GsIfNyiGbgB0RFWLvnghyR0sisFmQJAfiRd0wSPgvrUn9HawX
wvdkHVC9176xr1+CKki/Qse4GaOxTF0dvkLGjF9ejZZmCCKbcsu+gFT/Ich3iTcuTGgoRoFaBy6d
yDUEMa3h6M2n7DmiJaLMQstUsCVfYMBS0mfI/RUHWxPtv607gmXad77JRtfDLUv7Rx4ECOc+IFvK
dVFSTQk4kV6PtCoPcTLv/7nLl/9Oknu8xEr0AIQDyWvQ0hy4rnh6+YbMW7G2y01ukF4caPM9yKFZ
ni/8T0PLzWk3F1mkOyUC9A1TJ9qMkP/hbAjGExefas9ZU0DX4iYPyYGCpDLc1MrlzuMFt8CbhANZ
MKJuzXwBNWx2IQEDZrVCwfIqNrwn7/ySQ7o0kXYxSgdv7IM63li2AaFnfulXP/9yAEWL+LeO9/om
YlJYfoSa7pLYxIb3g/hnKBu8JjaSEaoESXke6VN3GzrA0ANQ3gk3l5Ay/WbjvMduZ02mKaBC81eK
KSgoBKwrYpMS5NofT+I8wJpmLO+W6Vg2MLepOIbbk1JoUP42fVDJHRaQ/+cHxa5NTph/XAEsuQx5
6DxNtY5KYHsqfxaPj8uVVxQjwMX8o+9HmkuJszaQsXb0TZK92Xt3hTWbcDk4SB9f6vHgDH5RbAHC
qwwftbnbenEs3rSqwQeafgM/jM/cWwNaIUMsYptAmUvzrdHWkKCnv/pw3tMh/oYDop++4TbquuXD
zCsxNKLobYzzGyEAmDnOTuwhIOYAWIfsBWfljSyRqVF1X3lW26uFDs+V143r7ke+Elv+0Dpy9laY
F9x15Stjfb+hWlRgcBt7b4E5LkcA2gOY0OGIYBIO1xxuB8umkPlbqNqz2sDtfe8V8ZQLqi9EE4gl
xfisNr7LcDIiqulzRFZAF7Ti+367oJVOuHKkJHxU/Klr5yjuielJJi0pRIEIk1013TrGyGmo1+q1
h2AiV9ZiE0LW+uygJsxsUYQksnzoURybi/ZrwwCF3+7/30dEu1kKgi3LNa8mPs3IVjmuucu06/qj
bOnaVaQsCgZliK/zxT9LVRGWVOWinRPKTrDApeQH9oZrZhSPKtdraJtP1GyWK2Aow84Btj6By9RN
Us28ngJuOkKo1pr38hAyNtD2drOo2diyw18MiOStFLGC+4UMCjEi4z3scXMetwpUUV5xGpEhhS8s
Qd4vhgAZgeBA/gw1Xn8suF9/PlfNf1ygS6Dky7fY72lGUnrBHSxgQg4t9sWDNCXVKthScuZ0NgxR
g/0UCrgw7miKSgY30W6+JBZygP2fkEqvhkS4Qy6T2m9ju2RGS8tvJGbWRfOOm+0GVIWiO78Wd3Rt
MtjETEHGH2JEqd9Oq+FJb7Sx2Qb046icAokpf0dZV+neZOpkzSNhRyY1FcU31RMU07zK7niekkEx
xQcvdZgfW8ok9HqC09GOjG1Ka4XZhOfYEItnyDdz5Vo1d+my54OJGkQoeV2oLO1n1WX9DtQOf7Yr
IKdh1XuUYfAiyd5onI8dpgakpt8LsjsDNCZY0i9aRkwwmcCnmZaZ1i1HWZ5lLKkWi9+I0Czl8Uu/
F/h2vcQcW34u862fYTonJBLfXWt3Md7pnXD4OIrrEmtqHJ+C15s4mX7SrTBzPSp0z8XyOPwEfr/r
+SrrAeYBB0M25Hcm+HQoTjL6L1G9A/ikp9yFR2KtLNROro7gn834bZ4kJFzbBtVpmvy9FzH7AbFQ
WY4AiI9QmnRpYPd+PT/FffVMHAS3ue+MCU6Fb7criksLFdn2arIqDA1qsLJBwkbCTzS6pErWv7y3
1SM1/9U8xDwRHxv75OzpUdf5yIxJYPI69Ebm9vc+FFdjnbhufMY6n6rJ4aJWo07PTwV2buyqxlvC
aOLyC/ckfCurhCF2pbcbH9ctacCA95x/IHtvx5TEZ9cbtDuFFi2RYeeIXxU0yyOx0LFNAOQ93id2
BWA+vSOgka04nCvDgtaIxpyOIywPEVOHj+ZArEEQdyCzyJ6fiOniL3DrFndQmCQvGEM6tMG7ggqY
VWqAOTRvj6nNDGAgPFzS0hyJEpjzPuTTOrZqD2cDsHShkZHJpifj5QVUvnoxd6AGrdnA2s2rCoqg
Sxyqpt4vUn/YCcoqMuHjcA45GAuKYUu+YJLx8zRnb7/Op/YqwLcVAMT/7CZy5GrEsHVQdu7R4vpf
Uhjg7R9rI8+hRYG8OBhe0k7HQeQrwdYTWB80GFyAs32GyJYjl4jTrV1SFKtw8k7sKQOuBEm+T7HX
tdSjkhhNsxKFlXtaMmbX0/N9OwLoMZz3h4AE1TxPmZHEbvA4JDZ1MKbbhhP7LI1LhgIMDVpDVWF4
y09kFuyMpmtzQOO360kqOJdMtez0EsX8a03orC1/Cvw4g5MMDRxeWdXG2Ou/bsiHxXm+QGP99N/5
17XeRg5h31894npGlj+vON/QO1RVguT2jqj0Ihsn66yf4kbzbkuAx0PVK2wWjSvQz+rt5JFIsM5F
qEsvJqaImwMl6/+XggJMQvz02kWjdoH8KHu21RbL+OrImyO+8ULbMDaL/IXKAUnymvUdLA0brNNj
sI/AgPAgzkAfcdLEAZSEVkmA/smzl+3dviMx1wO5r1k8hKfQXwhwVWeBbv21Hz15Y5F0abk+yFMz
huD9o19CeCpo3qbaU8F1bnxU2IPIGUjjL4w/1V6fk2H3yp3KNowrtkgtYUwTQEYmYL7mBTz+iXAL
m3gJ1Bvj6/Q9KJ6RLdQjTsWv1lNTKcb2HPLuBBbnDsPjCiHjxSoV41AHR5awDzrfpRGLtHGVLaMF
mAHPjuNfqMyidCTR4Cb8JCUWrrNSs6+y+Bym8pceHfD+Qi4IuqBI0RmZd/4eR9dAKk1oPhq3gvlP
d5tIutWA/gclmK5Ytjp0s2+74KCY1p90HCsDgFB+CDvGJbJy2BQlRpa1stJYcVx1b1IuyPdlsOO4
FRF1Q6daxQC6771tTIqgLyzKP8GWASpH6FnbXmAAOzHpV1mIWVckgEhkFhfDo+1iFtbnQf6JLJ9a
vKterrucW9pSSJ4dX7CkX7IhK+tYnMjqKg8Nu56otTJd0CiqoVFJDJLntWq9JhAy6Dn69FTlbu6S
IihIuIgyAolynM12wupjV527qTAywvsVzYDnQUNuVStp6i6jzNmjvSAbePQQ3N+CGgoFZUn8OatK
C2wV55Ga9LRt6TtE+AVcCoWd3Dtk3QL9H6qfnq61T07wsznSomC4NfrRSVjfh1KB+s3S+dBdOsUA
b77L9bRyxNT/y895ywmCleSZnmptcYArofMuPIk83BCBB8kqv1k9DF1eKHf+OHOKrPdY2YFsCfFl
NoMDPmejyiFvYnkByDneJqxXp34Uk7cxh3XV6s7jMWt6dfoVKNRd7ioJhxFvYM4bHxsD6YXVadJd
+tC7Ic+6uVqsbCPc5korcbo7zxPGxCYz51Wk7kV5+l3ky6kDAVCXdLy7VpowX/82jLbrqZn7wO82
dZi/tvG94I301jkK7Bh4S1+sW6JEeqdtrl/3O2yNOa1urV3tKfQ+/sI+FUIwBGfIyZOG6Cfj+jm3
XnXWAhDy7urMxGdd9BXwt5b4Yp3C2NhE6jrh35k1BBMd3f8PPmOJrEibspWoAu8PE/vgyOsm339C
y881Yq+8chpuJlzKGiTnEUki4wDbMY7y5n00ZSl5hgaBuGm99NJPSc1ZA7+urArudNPQqRgYY+Zy
kt3gY3AiXTjCKfhvbS4AYAyRKeF/u4ndTtRzslINhZqXz+DGUPD3aC4XZ5kUxIriHiAHpoVB2fTB
d9PDnT5EQaHZxrlaN4f77cRLzFZ1op7YAFqCvFQzoOJt4G2O2ZFRawFyOgCMs7RQ1yr2xs/QUTgT
CpfXlb1Tr8fIKsktlI9P1DfdCu6n10pCsTVJTd7/PTNDm+lSZzwbKCBWAYJJ2lz+evV1/Ud99xjs
GGq7GU8IZZ+hHp1xTp34RPeQPKKwc4qiHN3nr/isZj5KPZTH78A8XgKAKvGJ2gcyao+fvpXCQ0fD
QbbNtfKZXBZPb0CMipQWIEi5hknJ/mkWYZ5FE421M6Sp7gFj+LKYhUNJgzanG1JZK4IH4Sx7s/+9
aDF0hQosjYqtN+cCmNrHDZm7IiSDlNlbaL4jIhiyY23d0d67kz6iycKBi9yeLcKt1ru+VSMgoDFQ
/fn40T+r2OioHP52+2GMgRBy+JIvDTTCwddjE+2hIpUNvauHd4CT/3mQ6VLbx9SFOBuRgm96kji5
/fACzDZp2C3FIZdCjDo+8lzHEM8OhBGn72Qw2PN+Q8119Zeg9Ja4KGxf6f+dhD5Ijln33umKSIAg
EBoYgWasgxg+wf5p+0bALhARUpyuQ9ufpLFh1Hb55yW95Q4rauQNt2abpa0j0OtSeMxjey/OleyX
M5X63McSFwd3/WT4IkwdPy2Thw/72KQsKUgKSxs+yvTRdm9NI+XBHmQl2bnxWIdUKvCPhisE7U1d
oNJJaZKQIrzlSWPLKx5TeHd4dgwsCoiKgBD6UGtXgLOxVMc+dXHgBg47VhdhfR4zNnEDRVSPKQxZ
82gHeldzst9E7WsUF03RYogJkvzMgaaHwBV8qM/6WyvZw8eajJTLi64PawYHjIFWJmtXVFDsF2hi
PPk48DB/xbEn02EjdYwcxPmG81G/WhyYoYlOIJ8EqX5bmhQRCjCGUbULSHfSlU2UzmhF55I6AKNK
0lxSnGSbMA42HsowCkfSI+pXN/gshduohQvU0ICvtSCBh49sxwLjIkS7A2Dvi00Nj8GlaHlx0odJ
/EpUX0IoUhuOvGv5pKAmFMnBWsBE7OZBbxMsAHrb4b60Ctts6UYXqdI/MJxV/tLUEc3+9XGvs2oI
ypxxwLutoMJxLej+VwiVCzy/JA3xhzG3XscuKJ61bMvD9P9CCppvuGgPrpfDkCBPths1Nfe1sEP3
ubqCFGS3mbqoVPE0hHLe04/XMWdd9lbJzS1vEI+8HqHvLR0vYo5VV664/Jn2wloY0x82rPXk3b7B
0mfqZDx8mJkssE+rJfbLO0cP0BYLc2TlBJjPteEaSJxNSjlAyjYmZI2cKdu6DyopY+Hd/8rfJucA
CguijQpSVNnUIRRQR3BenoGT2GVRzS3fY/cqu8LkX+icFmf5pZ9JEy+/SqRVBJrg4LGQkAK74nzm
wvDLgvtzpmHySZyJ9saKr1CUkJ2HjvZHsH5ocVD9deqgirM+RJvsfyooZ8SEhhN/rpigYPSDWgiC
gBR3R+3eEtXhG+ol0NPzjMQDfNIxRchYFUoM9B3o79gQEYNGdo0DPm8mtDq3wYwH9k0k7jozPYIj
qE6c5V4jMiNSXuBOiKZg8mvV3mHNSAFrggjfXTUOWkKVnjVqghS/AZKHazLbNxGTK46PxVMgYwDt
L5KCjGeD130158rXVu7BCQaTiNcWZats1jsLTRbwPLQGIgU5OnHrA0RW0g5Uvuk3sZhOZH5B4w1h
E7dKxiFHiZ1wvtK7G/cfimzYM+pU+/B6Gemud7ZLb2d04DdfR5xJ3W1yl0iEpRlkp+EvUBL3/LFC
Gtu9luyHN8zhBXcKHoxK1xYLWWLBQQk73CqGhGxNdfBGYpYGdkxhCn6zaDR2KV8tN01oqlfblrsm
oItL+KPCkqIHTIkrwSXnt01pHJ5vHbOt3WbaOKmllpWS47PrucwPiCx3yGfSXYj88b4yEVe6js9u
qaFy/B9IADH10I9LaslyZQ3DGT0dSMFVbjnh+BcD2wJuEcQZT090+2Jk5aiLhWya2um/mZmeILTH
3Vj4h1R6LXNi3dZnMqxi7Q827CaBSf+vyWcKIRSCIZWZ8HkI9aVdtdyirc47uALOwbeVkXrYbtUw
/yF3/pEZrLQkYEw3iiL7FqzjkvyFfq4zQHMEJ+s79qqQRsBOw+pnZdClAumtF3XgwLoOyQaZemVM
hNnKtLjGWYhAeD2D/I+PLkEonZDnM7ksG23J5TU9+u+r//uIAEkRNo97IdtdzxI/d5xcIAWpBQ6I
JDSbKVxRTP5SVEfq8bdhe/AdQinGLim5OvLso6T/PBL9VNDfruk3lqEYcFO5u3ily6WkK1b9syN/
oQQzAxheNddfEcmm2Us0RSiMAHEOoDe9kwfGAiJgjFe8sn+SFJ1vvZhRjEV8i1ZQMNAM6rCqoyFw
8v0aZRUOX84lx4z3eeHhqtH9VA7US55pFEGzoSeSEprSbqk+z3o4ough1PczjaRauov8Jqpj0bqw
DUG3R+GT4KgsyekzopuTFS2/ofkoslP3itf3rKAQ7Z1LO1i2dzwj3BcDoXzQyY/VrfITBnb76T2J
FAZmaVS6FGEgmVaafN3vksRFtP92eDMDDDK/5Et15tpL5NN7HWxJvWmUgGOthptB1qNk6clxizte
naJXJJaxNXpRvm/jj5o+xvxj2/IDPr0KwldrmZM053bXHkCKko40JRVZFySMvQU3tOIPon8LFSnp
ggX7p+IVcdUQRqSV8nDlEU8R+SnpL6o/Sn006hj9schQ00VVqTcoPe+kJZ+RKqaeh5aHw9f1u9E2
hwv6r4JmJRZ1PlZ7acO1/ZwOkuMjNaCVEH77arLuFhcrcub2tvk0hCWNJl5dhZAIolgD3+kUoBhl
9ltI1zZRc778tGYYwfEX962wcgZoGkP95FAFngArxVzKAimHJ3ZpatBmdCf85wLXFDm8JHnf4jnh
Ci5VxQ8paf0UOo0ZugP4/Z1stiK87KdkqW2JGBhBjOp2ei8niLe3U3n+YTIo2+72SQRVd9Nsfppe
ooViCfSdXpigdzF3sQCN9vq9vgFMyoqji9TaDntwlu7mlMpBxkR38jauoXKpo67lQZG0QK3lhIlL
5Li3uYbu9cXugkx+rOLepgjDe7zfIAgUHLx2XYQDZ+48zWVRYNoZDMPWTk+JEHkGyXxSvl8eUy73
dKMUNynZJuEXpLhHqEeQfh5giy5ElCoM0Xm+CFE4lyOaUbFvfDpA0zgzaSOrqBuOyzWcUq6YZC9N
D+RCbZHQZAprxsFoA6XqbdhNY3GqyA+5wGnEdlLtToBcQAH5T/eu5tkf9lyNtaJaMIPBZL9CE5vR
LJnEyLl0WUEftppSLJlmsrZhqZIN9z9pC42+bMF8R/5YqC954rYWgPnJc1uS7E5ZVMKRo7MK4N40
4nnv7Qn64tYslpYIlV7t5NVTxyxFoqMlQkoBrhf1J2nuOb0onI3doE8Lk78aQ2czX80qIAojf6lr
btC9vBl37I4HFWhHeXT5JsYK+X2rmOPeks+oOUOxtYEprH/12oZQ1Gsbc2B8Pt5mT1yCblRfqZuW
jy4smj4JSutLC3V3jrZw5IAytEgsqC9MwJ2lS1GETU0AZmM+YwqoZi4Ce23mbR2oVNgGZTcDBseE
HJQyp2XA/+8EUFRyIe7iDriu/TT5yFeN71B2K0DSOAKzBUsbMLXVTeSSvYP6HYlOMC3AJfeBDvFZ
2oK4k+dG1TnFUNJ500lHs86NIS9Zt/FuYWYdra1FxFPxgayh820Q4fPPMfoHNrYPCBNI11UU3lJQ
HzLaYqKnDUv4fLAVQQy0EkkKdBQvXmgofvKboNRd2FzJ6NPiwP+V/PS1bZIS+TtDO4nllOCL0gEf
cWWVREVUL800gjMXXYCLLsme/GhvgK98+LjJzEK8xY8lxoE80yzIMZSSnrhYAdcTpTYkhp2aJJUt
XeCmqc4pDQkyZ9KZ9CS/MZjR21dR+SdZ6jqT31A5EErxOCd/IkUS7mBi3Hu+EY1OZjW8X9BaKSNP
KA1UAElLeYCZA6YsNv2fHDfhMgcTAodNmT3wcR733n4rIsvorrBVeq2JdHv+F59DVUvp7oPkb4Tp
IV4KcnCOTN0dULK8wINQ7W1Z95zRRM9TEBRKQAwoIDVocgsQWWocgSHmOu90hUJ860rFU6u1rHcp
zCJItl+sMK2OCm7chYvvjWgO36PU3MH0JcYRr3O0STWAaqj05dmG8oacF47EdvFSetaLnO54zgtZ
umYlyNxH6w6vv7PbTjAy7GIWSZ0rKsEdifC4DG2LvzlLh3sWThbcA9s53uCX1lGtULOuoKtPrgG0
/1OXqLLl3v5MObqe1QakRNB2knysA1FgqSRaDFjZeHf4uSKWGjXNJkOsDVzkwvp/EVC8LLm7bwIv
5QOzIbGr3mHoWARZVVFQpe030f+1CeBftZXsPsWFyNSLdalgYksCKcCDjhIKP9cHhAupqAhlEMqc
L5STdq4zmrHVsa3wr2x2QHDqY6htiBZUOqMZW4kyrPN3IdI36uadKxbzeQV0aY9IEW6B+hTxQmAL
f8+c/EVOGdEz/pQF+6Vr/rLoUTzhqxqIxKa0CUyZir6eJYTqLZZJhMsNFC1NZqoqjw8VgNsNNYFw
8R/CJLRqgSx9Td5+MYDh8wgkgW1L6+F2EZAGrjW+k3E/Ra9bRuXGeUA50CmdtjA2PWU027XQdo8w
Jtwno+llnJeeWQfyFv6LS7HrL6NkWzkYbh2EsjS+D0yssDzvKvKqMRa8pyISINw9Dh+H0thilfI6
7ZUYcVffjNPasMyBE8KvgTRa7WmW6GJrxzSbYg3pByv728gJ7zTi3c1GTSmSO9GH9fqB63A4ljWE
8iNoaN9dy7Xc8wfImlh/gOo4KaGz7HjrNhU/c68ZUo51i4VZNfBZ5w7H+HT9U2aDiRolvmnzSpa8
iLS3FfUgb0L7yMxEBpESyhuoNMmPVu8akXd/X587+fpk8hTyt8aglcKV+rrX79UFd4rYnt1ve53n
VGkABEbJHLBzAOai/hdMwt/QU4V82HbIlyOIUTk7NVSeMf5VQgvAKlmHZskNjtf6A5UndpGXriGa
+aQrXFRqmlwt6xrSnJDhY/DXhDLmlXZMli0hgvfiXWg3xQEmVI2akf1Bu98S53/M286zjqFswZHj
Cv6FfT+AlENPXlK33fFLx1UTn7GpJ77PBAY0Qrayf7vukVEOQpQHPZeJxOuiGoVpI+mFBNHoQTIO
y+Wli0VIr9XoSSFDmCYxh3FTgmlt7TNyg6IMj+fheBJPC62S4RJp3BVoxC55H8fkbZgd/dFHbrVc
kQnaFmg3x2EyHxM8IQrrNyUZU/Bissa68mrGTSTTz00XdG6S7uMmYOE7du2xZ71Wid94N/HbkEOX
U1j82vYAJdZI2+Lftvt2ySSi6TugPjyxFHTCK7KmVncH4iI7ngS3PIn8sz4YUJ9MyDhQY26+/inP
dWJ23YJpeMWVfyRoz7l8IJUu5xAmEyRYrW3JrcaVkkLZByV1lKrnidLLieWqJOICnu4U3RAkKGJW
kvcPxrMfQWkPjsmWN6Ri4RbZB61rEEETVnPnFMBsXV8P7XIEZIHJl6i8FlNOzz88voy5G+pQYb2P
DttBa9oGFeEDhNIApjV/DGzuUwzyDQ1YdVGWtUoTQjba5LOpHxYVU2llZB2HGxFR/nGgTLBkbsYO
etjmPlVSjjWbMZuDC2NARlKc9fGQk72RsqjL/PIif9WDKmIfMTOOVV8JnyMLzU4AJRbVDZFGn0hb
U5KwsNM5dHkK73n70AZp9hiPiEJinDUdEURF0m++5HcWucjdAjjJ/EnN44gQAH31aFBcUiuzEftF
T9rVZrajpo9+j9YVJZLeJtD1WivOEfKgP9WCuvVHQQY1jc5yuagV2FurhKL7wvTTf7quW55J4Iay
7AqNijChLkbBqCqzkhuqbeCDW0xq9j9F6iq6b6pd6QEHz+tihdOjGx8L7fv2rc0QFCUrq2f5QUt5
tRmELuI6WUcI0dLCMgY53zwlyE7cVr+ruImlFjwerAuy+s86AZH/0CAUQOQkGl7ZyixbbZG/gmO4
0XwFlGADB78ceXsZIERsYgq7+82/49uTg3SvNfx86GcjxKnXo3yUVWqZaZMTf7n76FIY25eJG5MA
abETJXyVmOjelTvzos8Px1i+tX9KMWJ7Cq51RHM9AxMvPg7MHkIY1PRA9G4+4dxcz73l8lQH+/9+
9NAOFC7RFCQDr3XyIY8CZhFM7RZhix6Au9VnbkK/ZVMPwmOQ7kjEUHPhxy7HfihOv3Ajy6Mhb9HY
niybR1OfCuYeVrTlMcqKOwrwjku8hIrxYje7iJkP3dk/ZQFmWJojyg/tJOsyAVKavSz/nRE6uIbm
M7Ope15l6L2g5viF3wWpjkk9Y6KHqP6Tkm/FWoRis8OWzAbUzBtw5glbomMnt75OUkEgb7sIryao
nbutaoyudMbjMbbWADmgqBpA5SWew4Z+JmhsFjlJ7d6dInl2wwGvVaRpl79p0VJI6PZrORPQSTnZ
FRbqsYBTLW7OemRVYwt3pn2QjIiZ/rBQwEAWxX+/KTap6gdn4WIASOIkOwxD/yYo/T2KvejpfhQi
1JBiK4jXR4iB0/Ms97J3acfmOz6MlgbWyOTRBEfLHOUojw+7+rdg+zZl6BnVFSy0qVwxB7qfEUzu
b1ciD33/u78bD7XXj2k21Bl7zxltFZMA+0oUZ3D1+taTtWbC63WjJbEbnnfona8herrwUerIi7jp
xYonwIxkkJVQ/v9wTnS86BsmjnhUCiUy/36T5NepWVxzzKEJJkz22upFyZ/ha2lZWzQYPlRmubzd
riNxp/w7sRXh5+SmGDjwldsZMd2doq+tg6lCBGrrfCGP2ORaIjHZRJXI7uDjvqU5moxIWhXIzIaU
9JSeRp7pk0T8hT2KFQIGtMGeRGHNrBitCdbOcT6i+A0Z9LwTZvfjXFgYbeyLQD/wZv4W0VRTfmfg
k6I0gWVw5en6nrhETQ1hSpybHVFZpj2l9RsFrZph0co6kPjVxRDFLIdwvwuLO9Hkc7IUOxGGTTMd
3ZHai8rVMqoiNxP/wp39xkmotqqNaNpKylxlOpt1Kx765Nza1neLGCr6yUxgf3XM0bLzWeDSZ/6S
9nLsPpkWUXGc3v3VAqNC4ya7t++i5wpfUfg1MXscSolmIJ9LzQ0w/GpgywJ8woDSCZX7N6seWONw
0XFOFJ0xpIMw+mG8PX+nrlug9jjvVReKjrdtlXUEK4G5+NX27wmqedVOsuwhcB2+WlBhVVR+NOwZ
BC/G88hv3qnQOnRgbyQIP4+LHjrfivRE6QzsPzIrDOBAnIwlXYmbHoKrH23b7+Erujy/SC/jdIlC
NIvX6zIcobrxJ6y1OGfe9jbuMgREIZzj6+EGU5rdWtTACEjuy2iUYl4OkMUydAk+sZA32Wu6kXRm
D7zE2w5NV8Jis+eO5RAeEETT6VQFd55kLK1qFrGc4gNIMuGvivFHd85rFzWxwpUoagCxfESlS/sP
EwDfQEjNPhe/zVp2nPuWtnYKnvb5eOZga9rLEA0r2xG7teFq0nOWyqD8i4HubDwSCspbUhcGBFyN
EMsaKAjzj6CU+teEYNrJdObrRkkMpZqXZc1904ralrireMsfhlAkWXOtGkWA8soqkDfof4qk9G1D
L7O494wHiHFFBHrB8LcLGImSyYh5LYSJrCS1hVKk8/Q9NHmwuEwwQemjHWRr3XIYpfVgjtF8UeOl
RflrZYSd/pgynqTuJyLJjzht9NiKxjAFdyufFEQbYraKwe6Aeqwhr5sl1BqK65lx6IWVQQizIKvR
GG+DQJRYqN85m/ug8MLCOABdiqL7t1DXSWWkf3ZZTNUcL53fIjjmGTPqK2iqH7U94wSzNI6t/yVI
vpuQtOzPdusq8QInv6n5Qyl+EzAabSjojWy1q7ExSbhBH/SsdPcU4CKbOjXxcoooNYYbIPrjNfC8
CZr//dnWx8+kvIMV8Olb2O49eog38Ns3OgGDcml2R1r3OWh2nLJ7CXsm7lZUMIOpXWMUzFho8s0d
Aa7ExyWJLsH4PZfc/sAKiTGpsSz3D5FQH32BJeKgRfticuTJ9p/QO8pvkFexb30ex6rRWyx1D1n/
zf1ufN4jwV5RrdiqiggHPB+TrZK9b3Xiv7IRBCUlyYaXWhOePh8TQsyv0NwpKjb+PokuskR8QF6u
UYgSIsO36V/Z/hrReYrAK2iZOXtHH2eb8g/hc+M57Yd+UT2B/3pzjgyzyLDzbWYXJanoyrG9/mQR
DwsN7yUlz2s0sjRgq0PDoPyyWQextNWbFdKpjmMUp1ixt/PxHuqxrdkdfN2zCblk8ysMYiwQZ+F7
BAvs8jDcA20H9gu8FpYL6vcBNxKgBXgntwBPXhWiL9+a8P/gjSbNZ4ZzR/RhOcrs8YijlopJIZXY
IBlyr/uKcte4/qFqeDoCuWUFs0OZCHMphDQyAVM58qsSWJVOkm9y+8rtXKGrdfv5pdYB7IVopHhd
D8oye1PV/uOZTw1jM502kMVeTDMl3yRLPGhVZJwCxOmi7be9TVEQ4haCTOLcGaa4LR6qoPZnM6ZT
RXyIr7TTjPISLBT7vresbZGLmP3t7EPr2QUt3pzudwnNzHf+CDAcTdBb++BrUt4bgQ5PmAWIreyn
nLwsH5NPy+C8qsdsZ573nh6SqfSz+PrN237VRw5A16vzlj4x1N7LPcBeFVgt61D65ooKPSpOD/o4
+Exnlx9YjOX5xE6t7q2OJ8iVm+TZ0/1vrwQJImdnLjk20NItMzGAU3xiwXsIuUr6yOZC2k4HBoRx
Sa+n7xk4MzypguIV9WqPI3eZb2Hx9szO9qeSgEUYRKuwBkzBrO1qutpaOltyI9sTP9Eku+pHaJF+
k7mVAmJe5j7R4aff2kS3pHzJXyvhTO6+5wi2p73jyjspisuSDtQdNfKssyNIsC+hGA+CvVb3c0uW
uPw48KgksLjLyOKaH3NaDcUz2cyn7B/Qzaf7fnaCs9HgXuXyDfQDLkj5x3I/S7mRqf6iZLIMHepu
KhNUF6k6Or2NRGk+q4o91KJMM0rY2/Rfu8uCsp8eyNy2ihaidtwAaGuApQBBOKdJVXqAien1Xz5O
Bb8NNhFTDUGNR533Rh5sHjFo/+choxDuG/rxIblQB+KDFcypv/imAXXhVgtEj9I1dIeLFurn4B5/
ao+gjphKMdNuZUVPAjDVGgm1MsRsEAM+8+RNcWcHA6vjdexo2EBhd4ZMJyw0GRluNA8wJSnH0ZGt
xGLGwd/XHMVezBVc6a7oasWUbBIbJqAwixxfGFiWgogo2C3PApMG7gfSNJAy2FnWVwjMY740+Q5s
aO/sGcuTU60NMRghNEkVkCoNLgI/SZLfsyXU35wwMee8k1bixbjHE+74WFQmGcF2M17aGCscXrZj
LnLdgClAqwrA8G1lmUQkKy8+XmV4IK2HznZRnFTX6nJDynOe2wRuMdjmT1JGqgtRMp7RuBRo1fW6
yy/fu/w3OI/5unf4T3i2kJgQhwtO8SjREI41bnrQFQ0Lqcys8VfVbmirdWXWEI0YRwAuiviE1KPK
rrEqNAvVQ+sEJdhG9isSkvuyDQ5c0lbWDazI4s5nqPr3LNom13LXizwr083ZtOSNa9eCZKFoDvy/
tKoYXT8sjJxXEU66bMYmrdwzoxw3paR2s6Fi6tdEIJJpYQe/VfdlLJn9cBN+HHgmctp3qQFiX7Rm
edj6zuM7d6gbtEB1eCzgbXz4hNpyCZuntbyqjQHWFSwhd8FldK4a2vABeCDr/Nz1YBKJ9Z5pAAoi
Wf+EDlkuDTEbh+mzlTqQWTzaR6g4TSpnaDMCtRd4HA1wn5dX4TxwicZ5Gj19LpF6WUDX1a1IsxHs
rwzHjphzqI85zeeZOWzpZ97ZW4FI4gcYexjZEbvGDbZ8t+nhAPrUUrVyqx2yxobukcuoSGq21cDN
329ojYlAKsiu1fZBmnyDelInzChuNAkGqicoe9hp/IPi1QgBw9LCRxbaoOl5dH7dLE9ny8WDAD7S
hH+XM2hnKj+WZTVLneEFGxmAh31OPWyyIN1Zh/qjQU8O4+8EYosGGge9zRxV3FvxB2teBhRcIxaL
baLOHpUU55qaqLTs78vbLmqQe13/PMHjcj0SnssoOo/SDBEXD8HtuQuKl7xsiG0YdOeNx5ZFh3fU
BHB4NmLkPCaXy0iwlwy+/IFFKwq95iG7wISS+WvqWX9ZQ+3SmtegDH9TXo27vZXsOXtCMqvxX1Qc
xXF/FCusv3qJeuj2OSfWfJij52VU+X4E1+/P8b3V0rFn4lFmrGo44koFkKT51qTzQlyQlMmZT1VQ
SAFg69Mvo2g76rKs7cCyL8YMju1JTzdlHKqDUKLPCnBEuuu8yDtPt51nwSkU0F1Rban5PSzgVyH9
8I9c7tHlMnDKM7VCGqc6JZQtQ4uuemuXxI377zWIghZNfthcWwtV8VxxfpIiSNPKtd3Je6F6Hvay
tkphhus4NfHTCoDctThjcCkWqwd0N7D23Vx2wYKUX/Ax8dlWKSJpBW4OPqtb+eaOkF+z2m0yS3jp
CRDJfJLc3fK+BUiHk9ReU0nI6dBKcDY8Z8E7mJwC9CmelwiLcN8IcN7pxrFdOYZsgJ4tFlyCEhRe
1czDbhaMT+N5jNW/h0mkorLVPnMrYcA4Z3bO4ZDjrU9QaquQYIGG/+FD5JOYAhRsgjVhEvthfVt9
nZFEeUMz7WXMjA/sc/5Lx4BCk7JqnV02opUqlQ5Ewr0238a1HACm1xpgMtIITPAQ9f8D5dm5IOrz
Jed+oR9Cm43Z2oVka5uobIp1e9aQX7Opn3QMP0VpR/gKglsgTErKALA4RVNygBPBAGkmyPiLbPYb
bLuA+F+afyBfymwWVgC3lMNzECKigYQPGJ1Q/0Wb176bi5PcLvgEql8ThyUCHiwqkRd8i1BGBKAE
Ebt1vzNd5FmIPd/JeYs1DvR5shdMC6QWkxZoSvizvtrnFKHimx9/onD9Qp0I02hnDBIBJeHRmGDI
bOhwbopIcik6x2eLJkdQkdRh+1z+71LJY+igAlXKx2wzFJYCU3nSioNPVXDzYrYKQn3PqzuBh/8U
ZfngUZbqUpSVH1/YdYnOgw/v8AKog7ewRzD3awTdMBYPHdLoVTDxu3szEcHVaAQlEtHFIjkFQNsU
N65fcu3epgQHj0AnwpHRvghwgJiXbqAN85TsfnKewApV3p86BfgfOTHrofHhCzCBfTleOeQBVhRf
GsTrQBckP6lEuhkiEh7GPYaQ32fxSos+z1PwHeRAJI7ppvPzSEJ/0Wx6cKu4SKj7m/JaNQlMqdOe
8sqjTB6rw24kAIzdGY8JkwM6JS8yf0pVASx2MveCl/2ZJSHXCzyym5d/oQz7mQkm752bdBiAafB7
DWOmrCn7Xevv1nffZgLz70AqXio/cy+gptYYWx5y9qymluXV9eP9QJZBNq/LSKzK1dyXTz8+OCpv
yB+6CLmnI6Xlx/eUlSgvzgr99jxNon+6pVWJZWbmeQgqUIa3pXxhQGTO6qZngPlX1t1JMdubfLZP
9e/0hGfLbgzp1MrJ1YHwovBFYjQRtPENqHLv0lGfocaSwfx60lsPGzIz66aprMoFthwGnCB1WjXE
iiTr732powehE+pWyUu1IlFyayaVmE3VqmAgChWa7ucoRA2nvoAm4hkPV8GhSasMWM2D7+NKoAnv
uZlLd1m+gEYiuiy8d1lpDYQKT6NHBkUFrftRKNk8nlXE/N0Q2kxLvGe8ttkvHkSlocbrfFK7l1cd
W1MFYT67eE9bSCzQ7Afalo9xcj/Go92K2qyqr8gwymZMakMpLvPNO8y961/GdWQ6bBkxOF0Xbya3
8Gb1NzZh174kqEWkCthZHGaTaf/TugT9DyYSQSvo/iZRNkVkW114rfmz6QpB8w7yIoOWWk+a0/kr
yO1KD2ZcMksIN4IK1lNIDXx/aP+oTrdoaO/P7vUgghvBIjq3Gos/eiFXgbQKU2YNQ2D8hn7y5DP0
IOpN+2oLTKmJMxkEPaLccie+2UQ+YsOYjWlCasNZjLMR+u92SgeZD2yV0aHC/4dHsWdg0S7Bys3Y
gKeVxT4fcneso2I7Qowqr3SJ/l/c0tIzKJLG/P12lQodHrDmrLQMkw+DRDAhe3R6ZYwo8F9Yo/cb
B1iR+YBzSHXNWDYUbITA18rgFQwa9TIvaJuWeM9zq/lMQx38jHkDPhnRxZ7sMghIYaYASOeToPis
FTbvrjyC7agzriSmZs7sowjTCdhvw3ZO+ACILLTdlckFctcdqvMilmtYQxdwMIkvt+MbKspwmKPO
OvAWuL/bh1xlKFFXqEqjcsiXiuWddCwSIZ6o5jFXYqIyxVSq68idetnVq/VIiCHt2XzC/LBk+HdO
rTA1MZxIiH89f4LAalB7zwFGEA2YpY3GN6jKCTi2rRhBGJd01NJTV66Kzwpm4MtZJaqUZU8tnNrX
QN5qSMbzCyuQ2n/InaOU6ef3wp3iR1JyKSK2+Qx4W9OKSI2fDepqQpLKUFs94Lizh0IqcSGw5vlG
ExgPognmnguwW6KAQl0Ge0g4jsQM3zzDCphbCI+HS4AveDk3cc0st/201amHFpQobnPFqZV80UOF
qxZ6yVVdzDQlcxFRJZpt0Lb/XlkvHbIJW9sSRN/UWBQVcPPbKtiWpJB/b9x57ky1r8y7zSLRNBzd
bQQINMv/t1XV9r0F8j0XxIRfVhvAPvZUEh735AZ+ag2li5fAZmuEeWkRlBIl2FaJ1Owl/EqME/ta
yBLbVdEnCdkyDd/9BruPSd5wQo+bSy7yr7z54jcTpCtjub810lh4UAb5SX22y34qNSCuLB+SYCTY
E3wJKtf4KG8hvxnekopRU2e7953L1I6fvExtes9Y7q44aIB+9topBFOAe5d8YhH0cyUmGk1PJ9FB
jHu7g65e/IZIyKPAue7rf56Rij7mjAkVoej6R5Skd+iY5aPc/YxB/EYhAlQ8IKZaBzYZhn32KcZX
GAUuzgGZFoEb9/sOIuX07q5NUEdBboXEN+frBnPeaCw3ul7rV6nmSeT/iaNptrUNeFn1Qix9vb1a
5qRuxmO7LHD8/VBZqWSXxVotvCqI/qumchn/29rMWo/za7LgwACc7XlHXbAHORuZ/4YjdnIA4P4Y
JrxSdMmnSzF/bmI1Ush0ilgGpFbJNIUiBaNZf+3Maf4VpqKV0LWxw5AeV9umyLF8by79h399KVEq
DpIJFz5gFgrec1/x9LJDlzOFzxSwnvtXeViB42rh6nN/8UfUAFwLIqhsJLXjEk9hin5qrNh7hun8
WlyNayIY3XxmwXfpZIkHv2LC8HG4aBgK7/CU7BtQbzuwC9BWNpnT9Euq5bg54TK1+p3JaVPrKA58
ddv3yu6+r6bwyJatiKcIH0PpJmb2D9i8cd6EoLgeU6s/DaW8TFPAZ4tWbXrljhndZYpbUxlJkJVn
K9eNmZROyTpVn+WFEV3qhySJKqHABhQhwL81mWOh9UM8fxQrfFdx6wdaYnjxI4tfm/n9vkI0PGUD
tEMRzTQZUoIajbIS+Izl5Ia9IFxUn4AKDn5LkIJCDdHucpqnwh+non1ZZ7WmQZe3JPuissdVzm3H
/Cxe/AdeSynr+9I3iHMG9QvkPKT9VGesNd09j7KeN7QPbtk21tHxSgKzWDlA+XGIjOHVTHqh3O4T
6NfKL6OJN/PpA+d3XOXYmQ/KHFOCS5wi2GdPlGRS9Ixg/Q1XH8LaixJMLfqOo0ztzNT96BU9/5db
Vg1OXi0bOlv0WA3r69P0I0ZhfO6MQrMpx1SKRul/wcnZaF0dtnNxe9iv8LrWH2DPZyFczIDjoow6
il8/KfTq/4shDXN0SG77h9h3/e6/XlJv4U83vAwujPIa2ZQCl1gUiJSK/G7cjyVu3vwdOIfxyFor
U7WWPZExRssJrviXKisuSENw9U1/htfGIig2qDNRTdj+RWqKZfx1DcKicAp3UfmCT/PYFNdpBxYm
El1qWwvuQyqhhJEtTE16NBglVSqZlRA48HWF9MoJsc8BZ4mASr7mIGR0QRa6f77EMwVB0E/5+b7S
oqs1KGSN/Gy8hDqpU9NzE+bsKw5CUXj3u6QOP6I2OhEntmLdeYWKVo84R6QOHhRBcyxhnOpK2KO2
N/rNjK7BvkGJUrQQoEzfPO26d2GvZl1vHHAUTjtUkm2m8OPJSnuL6wvbS8yjPc1n38m/JS5D8jNI
dL10XWov6+9q1FBhk2HLuIuquJt5JHxNoX4eT2TxUX4xEPgRcnEokbNv5IpeFXQWBi/IkimK29Eq
Ihql4cZ+JW4JWnSBgNyDcYu6zvLYont1tVLevKMPxG4uoEbabASO6nLsZXbMkU0b+ndYwikwb8wD
7sc8+9HJA7NoWSJPhjKLfyMTkCxz05O2+cl1FnUYG3TzbW3izMXUwGeF2BWvpwDIgapsdkw6DM72
ml/t/H7DMoSp7K2faYm7nusEXjbTMdsoZxG8Q78gQ1Mt5HRimeLqBZXf5qx+66AZ+oYf0JJDALLt
hMcgaefg/eayCPunHdTUDVc/FSPEvaE6blBF+s851Y60pvKkZrdDzfrrPX9Lrt/uih22hTKl8WQS
0TBz9iE1CyEA7dZgMNZEZ307vkoo/ffxrsts2RXGo+bV7OaIkMHz1nhnZNCktRYm4kNOlJr3l5un
l60Y5paFgKS2IqZJZU/V4Gc6N7gR9H3cw39qswnFqxmVCeW8BFHoNa7Pg+Mi6bUr5g97puoDDTUb
MWxSEE0/5uDWgZFGm6gEHYCHcOOj3XUy87W4ESEJnQ+54Kbm3k9BMIoj4JrkOpWpc3rhjTjeFl0m
b2AJ5tuzvP9h6lrOeKMOjqHb81w0CkUUD3uofSi/eQUrjJ9NeBlT4FwzyXm/DPjS+561aVfJLM82
kwv0plofPjMa9shBeXGXtFNOEg5zoHGEdYXPX17fc40tvfQnGRtA3FYDIjjm5DnUV7juF7fDCJ8w
ygc6YUSoZKv4uQXiKdCkj8LI4WW6Pd9ukffPtFSk08//lFNJkjfhODkGohWcqi1MV5ud2RiNkebr
AVPNqThx3m3rzNK4dFD9YTPiRa3u8rUoCuhCoRAA+HkoiNT48S30xqqKbAhfJ9z+8CNIFGwpMGvC
8WcDiRxvc1RDDzaLa8LIqgLw6+VjKctIoZpcO0zTvUG+Q7om/PyRBJE9Wji6ElkPTBK1N4ALfFPp
GDZV1Rqpf2hWkutNkis0Dx0TyowIZYXa9+5b0o9ikakJMqHhyRk0RuFNzdswpCF5tVQQSFNFkSXN
VRAMypAYiziBJh29zYvg7ZgWgT04hRLwhggm+3p8DpPzyrEKlDgglDrfAGXvnP2/quTETa7G11z1
MJjSUcJwXNr9TfSv3IAwHU2nCdQ99AOZwdvi6TQCPg4h5NciV8H6dS9sKo8Jp75itqHTw2/Sjjhm
hYxFMfSIfokUoXPmgzlMNAeXobAG5cUTJnD1av05ykHXj0V8KjpEaAjLimLJ0YmHKaU9JzsvmXfr
Mj0/A6K4J7zI5nXVSB7bZFFEskvpnLoGxm197eUrMwrfL3m/+aV5OBRozgmkJ5aCbG9QiZ/rP3kj
LLT0D6hhMIMHHgTJnno9FP9q6W2FHeYWx0jll4O6J+XN/7uVMqXJuWuTNEhXDrxOHzu11PpTMv9G
ew7HQCJp3BwhfIj+nBv1vzAEQ8Sl3t6hAhfgssJzWTSOQgKeAZzUHWzaN1iKIybNz46SBo2lrxBN
qig5tRYuDqbDazHB+p7O3uWtCSfJOcAOoS+OvJ2ksJoOJdK2OT0OgvMUhJk+Qj272XsaS4r63ua6
zxZgEHxHo37jYZ6uJ683unS0W8nl8n/vumBqQlvtf2uoKqZAM0YoKNt9DCTnugjJTAf5Yre1jLfq
2ojTb7/H9kZRjAA5RYxMX6tCwUdj3ha6cVGnbF5cX7hCTzGEteFox/CmAEWS4B9vF7S1AcFxtPTW
WGVKY5jvJDduJsEFYDQap5FB0LmscYg1nTyKE+NrbYwn0tIasn+sEMxz2cFqTarhRtWyOKsoznSI
bE2R6/BrwKzlCYIz5YNMiZyisFlErC7XJM/vLjR0Eh4KuKqah59qHEOl6QRdNlr5gU32T0cDO1BU
YiYZnCA/xMj3STUmpMh1L/4aowZb7fzkA5mfnsgg/lTLZpUM2dv81I67L8O0jNgo0nF/X1dkIYGK
XqiORo5Ko7kZQyxYe4rHr4yrMy7kIuktxASv/iASOH6+iZIr2puaCabbiBOxcTRrlBMQKPXVTibA
eQoeauIbgD4ZgKlBz5tqXoCU3FbzBb0fGS/ra89bANtXK4z5hSHEYWCRWoiym63E6tmbXHKXDRVZ
GS2JCKuhfGjp8TvRmbNk2+TbKoeS2uKjfu/8wTwagMu29okuej+17/0mSElRcrbfuw3tKXigPUB1
uFQPHOv8rN6SX2IqYSUbZ+eiCnKKnQ2IR0b2mhNM1JLn1xrwsh/Af6/3pz3y6ERa+kJ8xbVYcXK0
3m+q5wttAdquvY1Tp1TZiwt+Ep2TS88n+lXRKtm3leLFR6dzyvSZtmAWoeB3sDYplPhLDdfpGjr1
oBtEItmG0d8w+3Wl3dyqnn8pnnFCTLUVZ5gcg9QMkDYz2xAJfRiUmUrJBiLX9CAzCqAaHDkyi13j
PQXBfO/xMn25Ac1CmDrNPgQcqxdysh7tTkY+TLL3fI0HiRFNUFGNffhQ5hgSlAyYQR0y1OTANg6Z
IvqFv3RMaWVsCN4paodIq7vvkiNig/z/xh2TaF1S53oEFfXpJQ5a1MKKNGdA728zTpUVFEi3w1bC
/kYk8J7o9gMJSB4i6ys0pcohAB0OanGr7P3n3J8y7U7dP3KH+N1g9c9kN4Q0t8Xildv6cb6sX9Cp
Z3ziwhChRD4hWuOgW5bza4yB8zSryFKgn6v79uW3DRWu7BLOn2Y/9w2BDQenOtIsdUiplh9NRSr4
drBVSwkAMX7oRaRieJA8X2hNjDS3b5u3IyD/htcpLXd9lqhwBrbasNSAKGVAQgK4vBVzXbzqhpnT
Mbhs3jQKGu9ppXgFNm8LpLpNe3EHvOb2NFl+46tkXW5WsE3Qc+Lago6fqKXEV0srs9jv70wVmbiy
4xRrlTSmXq14vbXpAZMXXPmO020hWzUGBNTSYKz5gKE+zLP0ukJRWlINRMtF/z4I1CNuvH0ve9rS
dj2xnsgNQkxzVQ0xDtNEU8aawHUsmE1f8urGaRXpi/FCXjXlQMLGCMrUoofSDHD/mx7wsjevhgYk
Hvv+lU9nULCt9f2w09rIlMBSe5cCcQqed6RWU5Kg8p+5dM4Yl/GEvJ5dFCHufPstGkz5Mo3uIr96
v3zqnK9oMPK/08Qr5lHxvtnzgCGgzhL/uue8H+KxEd9Kcg4Vr7dBoiHZllmujI8CXSC/dfic2YSZ
cuaR8hfDfX6RhsLxHWNUgRxH/M4CxZAyzfLKT4pdIBmQE1/rfgM0kxgR6JVLS/ozcxcVfQD3nVia
7AqTQ65ybGqxM7sThSNSgoa4ygga8YSacx/MS1dVHrlFP4ivXUuX//LwDePjzJp7CZndGi3/nGIh
NCiIxKe48PMcd/ie566oE058PD3tG8IBoVcw5khgzb08zheV7EVrwNEWTXkbMO+JyhVhmepDaC0J
2/X3/UFctxRAmDrlpHkh0+87gcnm8uLyIi1OvQS8OzNF8DMIeqUJzioZXLT36VRyTSvVRBs1V5VP
EN434XDVsmCquQPrjRc2SoQhTqipHLRPn96FR09WJxJ1DZ6d0BrJCMBPPrtbCYuaDIuG94oJ1RbD
QPoqEQ93AGaIsU2cKU95TO2p0I/dv15xYZ5bmmOOfDJK6AfDlLIY6UmITLuIwUDuNYflw3DjfVqe
fe8atRubzDl3Uikoaur5SHlaLPop5G/LIkxSKZcAVSrJA8G2Fxhxp8i7N2B2ruxAsQ+CV0UkCaKp
nl+cvjSH/O1qj5H6PjlmOYWMBlvcXO8RSqSp5t7mTadZdDLrVTRhHNtmouwYaUII8AAofsBWMQ3k
i5GVds/Ie9A5S7XYB/Oc4a+UbliZMaORr5g2/sHpGVhWE1M3gW0iSobbMY7fTLjLO0BLKI23I/8g
pOeSda2zqRCibV2EbgtJEXGYhGHv1z/8eRHhWrtByypicplrE7arbhkPfPR/95CgMb1/MjqJKTir
H4nbLVtc71rmtP7RrvBzk+aHr4B66wFI19Bif+9y4Adcxbsq1tRYjdrsjkWL+SGE8oqSdkKku1KI
peP+de8Plj4uwxCc0d9LykqUZ4Jcme8/WRttQrO1LwLneiz6hMFMGGgtsUomtvvFQj5z5fB6WhGx
P1coOn8sXwLdZJJQRmw+dFs7O5YPIBbuKVjiEu7yNzqX0V5iknZbpe0Ibm+TB7ZEStUNMIdc94Zk
+tmA9B98SLt7vNl/vS2vmZ2Rt881pk4x48fm/hFNjX+vKCXILS0PV5L88i7UIVnOL7aE+EKQXBwY
IGe+XA9Bq5yobslYXg+I6c8bQeSGjPEi39aYQ/+h+ISjPJBl/CFtj7Tv/icI0ytn6c0YLPMptw8B
rcFQWVtvu0bIog4Sj710QQtVCkkzKdREYr8byIjzsU07Q9iWitU2MTYSrFIpm239wKSaDeWQ5XJG
Wxpg4VWf5vLwrIBZoigWZrTJaneaxYYcBNwxlddzpSbgFzEgqYcgGEmAf5qxKYRZk+Xz4fdjglhx
u8+Hga3K06leqTUQr9rkxdh+z+cXSCxV8s6cMrZ9trYF8FXDKnz1oEwJBIkag6emRj8YNIzwQAtx
NWLVS6fUob7uZwJOkLGgO0SEK9DjgIEeoy1bdGtV12UcOleFBFnEhw0hzo22V4LMx0DNRo0Wqgzz
rB8nMsc93MfMos/PAFCOky4OWG4WBDleStGtSoi/XBB5HZTnaMJhn5qCXbshkWshIox6DvuHI/3l
DDzukuG5GwqE+G2x+gaazrISOLzLNI/f5pB86Pgm0WxPOT6LKvDMKWU8fqtZkJtr521a3ejyeSsj
O3t4HXGex6+7BF9a+QVdj1vRnEOff7g4qcowjyASa5vt5aQovWXOSnubPgx93tdlpWJRlZARC6uv
1qwS/yRUq6fTGoSOsIEeDeh2e5I9s9sIPbC9r8Ycgq1r9hZ0SNb9utqk6HO03DdBSo3pji3p5dVR
nbJ206IwSQHwD1YdrDR4hhTOKKZebeXo62QLQPToIJYXxgmIwlkggdyPp6zbHZnOcmgNLac/+Kmo
XVXrRzV2rdC4g0mie4plGe+VmczlVgJYDLfgEMNNIsw748iTuDmhBNdhh2MuSVlTBxrftjS6X2B4
M7qI7Dl8VWPjRosPN2JUK96R1aET+BL1P2bwPW5IHVFOz8lr/BPPVMpVF4mVVywTwIinXsXuY8Ny
/TGlZ6dOqiLSrfW6Xdd8ONjUb5NzvjrlHvLOZE8OThy0ag8noIL0UU70bKN+06oIKkkE87YBCFe+
mGTy2ST50TBNEOVdECGXKVkybm1dpDMsTOnycTlOLOWnLCMFMKykpy1vFhSqBSN6Ub7wehhpx+ZQ
CqE+Sg4aL6WuFtLsyibL85zYGuH/ToH//28AWhU5l/YFa7sAG1II/v2QuEvItA/toLLJ9ZKwYkOO
KAO6YU7dvIYDW0yWsH2OE6FtZgIy4Jr8jFxLATZwMCgKNvdaMDoEpvJcKYo38x++YeyzG/SN/xdg
V8CXBR7sWAudMFnEyPsFbaYLvzFB5uDVUrHQxsMNpcD2Ad6oU6zmod5WRuOBQ94ZJvDqKqq0DpFG
MabINZ7bdFqutluHdqk4Pbmrw6Ua/dq25WkDvuQU0Xew5Fk1za52VRTNXb7rpg88jeANI9hAeg3K
a88eh9QnHdS4hz3Jo7tS16iXjkDphzrc0ApeaKOxo0+6D1VMFa646+eNFz3bXOBNIjb9aISTLF0k
cB9R5sVC0hNJSC21sxlZLhWrAwrWnbxs3wPlnr2Vbi/oSQyJ/q2xZki8Iyio+2JWSEeRp65zcnxU
sFJ1ZpA5AoM37c4o1eNjQQu2VpRQLFpeXQNSrD4D0sPuDRC+BT66bCBgNrml4T55BI/+5oJVYr8I
6LHC9NUr6Q3htUYyyM5hyhKQdO0U4CPZ2DzCJWFLelpJ+1NZEo8zk+9BHONFNcKb17iVh8VQiIeU
aa3u07VIyCH2QCscmRh99vOzVHO4cH4Id5qj2jUk+IzjDF0NdAVrOtLyLIPx+P09xRcdcE9bDCZk
IAurbVDN0f5Ztoq81fk7Z48vlD4j17mgjEe1zLODlOt/xNBmIfgycHwBvPm6u4KwWmWiE/zJc8bf
Zg1hSiHxiHfCf45EjVJN7+mxgl7IHoby9Yba7rYK08HvqFb1R702dbuDyZF1nDHSGS8b2xleyMQx
RiWww51cM+j87OFaTIgyqpFnLKfPHMZOo6icwCBry28WDQL4jFh1glWzpz1Gcq1Zahumsxu8VM0l
pwhiNSDdRDBTZrtMgyWzLp6lX+EJlCIzvvRrFEBE5yZSnlZZARBSGAQ5mmhZJFx7RKe0EsK9UjYy
VlTO7Vz00gm/XsSOwNCQ23PSHch6HdHIw6JdxOyZRZ2vzA9o3Dlw87i9/QiKwLnIHkzm4CRCe5pq
gYNZEnMIQ8hJ6QSEkct2Hbi8u3gQ43l0poidSkT+Lod2Hb8hklLwcw8bkSjZPSDPc+ak9N53n2Bp
nwV9pMgCNzy5VBXD+DNimFabW5I6Lp2+FdCGtaj5riMnBzm9XzK4hTNy05QnEuh1tuFqF88Ex36l
PW/D3iOEMQvZ9p/wDtlpOeXeY/3aXVVstJhRUqJ8TqYYrr81B643o7zSCHk4B6vXCotQgRfJrObz
5DhEs1Wb8ivqthE1LuHlg3FktE8J50Li8xcgU20qvk/byOfgeHnjnatVMcISkkGfrtbiR0WadO5t
KnKMgfUsgb0NsNqYSe42++fE/k8kIIlzS/QrlYwzC3OICeAlbV1O6XX9vI4TIv1RDK11RRoQNzmR
P3jf6D5IsKItXCXLLk9jENKDj/qqAf4VJU33HLJlsgTz3PjZKbmbBhgVwzW72xcre92JkjZSyWxa
QxEyR061+h2KnYR9kGswzsc4RVIHPzYFPnrUWxXaHHvF3yYkibDJ7qzngVbq13KGpcrgRzyEpZS2
Ji54Kcrk4wVlSHLkjwJMDI5mfWKfa9WDAioW//gD2sXEp29NDTk9ugJg47pKbct8Sm5ghQyBcfRF
xisc296HpHiSKUhb5tWVpkwf5jbp+qkkvM1Arz6zRMK7nVqdvv9ijbc3jprr26XVxqZyxp1FUufK
uh5/lYXmyiUPw7SWTuYZNI/FLWaJZooEVQwgXEjfJcwbQBdk97uU4/XwA5D6TRk9KLhAXKwHy3e/
bqKOaWPUMTOmfS0JNzZhoHWqC4KUc7pA5qDA54tWvm1WhbYfJ2booUEssfADRwKkA76L9p7BvRwD
E9gBNBCXvLUh6uDqpjzYb71LMI5nG55EWC/8LAjWOiqymOltw/4cpEaTeFD8wSmjxHunoMFKo8dV
/az6xllit+UyyhUBbcH3bBDTeMW30pZluPsYxBa3QOrh/g8QkMPbO26bwwPGmHcumG3JUf2kZEs/
XrBzSVeoBF2mJKYMkApBytn/0PW8e1Xg+kKo6rF5+qGxvf0mdhvTopA4fuDdIhdmMBC4lYvZw72G
OY7BK/dJ7RwTPlZ6+k/CqYKnSh6nEbir5prPXSiGOnWsNXtwIrONnZ1HkyC3k5Mdqqzt9a/ZKLNp
hYc8ePb/sqhLA7v6s629KxbSH/guF6qC60uSigHAcIXTMaOJtPFfrb6k2ADHxLadTg2VQAzJ+BR+
RrCYAdgGf1kzu4ItkmLd0XoAhcaJeEKrxcRTRJpY9ZE+v7bV9cklebiZUyaXw8QFYysEQCAwNwcZ
W1/Dec4HSYuYkB2lL0JFCmkK5nhiVA4XbE+RGajxoOsiV72wovj6ifpximYdsc2+E8y8c966jxTp
5UxqSUKDsM/V8oECD/I9iyqSlszRzH2tay/eBTzYAHz5jacp4mTkxqNZ0cEX/pC5bIOAgHBRndFq
4XuMrEGybYoXLo59rWehBSjLeCq+FEh6DUm6WEtSkl0t4dDC0ft9oLAx9boW5DnZ2pxDFkJI8+jY
5D/lmk2atMyqf5uRgTL7Uqt6ve+PXx6JX6BnFsn/gr3rcBFCAIdF3wTldqSP5h+ZUa/ARIEmWyPh
sPjBFwjPcXIKaVTmKycd+FKfHSULda9yDv/GULdptjV3fh9Xura5pWBXXUYLSaHDsHwCJS9oHmtj
ZcQQXEhedhR4w6zu4mViJFqWCEUgs2XC//F5b7MZ2v2UfWchGxNWAvc8VnFNak49On24wGFQK53d
8XsFuttYkFJlxADEjPVgAHHgWgGVtnyDSWqFXqXUlBnLzNeYnpm8UD9R4VgVAzme96HLFN+MaxRW
Fjmqbb50Y1uogH7L/GqJHJa0CIHZ3/YKqoCg9FQnf4vlrJElCrgpYd6yd59YH7Z0wPGQcbTuPnIx
1OZ/N1GzWF+qhUTwARvqLqKzlf9J7A4Snsvt3yoZjku/2RPqtxvq294b8B6Dx0C0AcT70vZ4w4NF
r9TG45ZnM+L+lAWYH12j9LQ8MIycqhA3o2Mwxgw5yEJk6WwAQpn8fZ8M4KMoKZCioJS9YdREz+fC
3RYwTP+USymhYOnSbSiqayJkNlHwwqFgSnyMPXLTPBk1RHftN08pW2QXHIHp+7S1sZaqVXekAoBz
QZAxHfDNYLxG/YC82yr1+WRRtqR612zMclDHGW2XOtwo9B9tnds7dmLt/0CupIrOzWZgi1bwQs9g
MUmFDEW81EnOWvQEfzCLwX7uusgmqRH2atWUEt+LMHbwphsMPm6aOH4jJcuGg+/1j2G9OG9iGFtG
zIj54VqIeFNSiB84NxeEY6ZMV/J4MiQuGSJeYjBYRr5bE788CzsZprZLNL+OOpUTsrGIutN9q3++
mEIGkZFSpPwGh3o7BDHOAWNqe/MFQITQK/uyuy7cEfSHYNdaTFXhzv8p/nRXOT/IsA3Eu1C6iFwv
9uTcbYf3Vh5E4soq4Qd6TCudKGeaKDyD0vT8mKWqGnfQjZfE9rQHmagGKwIkYXLT3bFPOJwH4QRj
z+eSZrcbVIrqWkIvP8DxKjAuAks5HwPirEEd+HJXJGWD5F7PpD+M6T6SC1c9WTpZc6A5CAl7NLnY
fXiQ3qlscSjZa2iFXZ1Mi7OAQIGziahFVfD4QlvJDg90nQK9pphK/6Z62MLNTDixs1TtTHBX5W3t
D7q831HJNZijMOwbhOUit8dGulgrDDj1d7aXlwGTYdTzh60VnStU+N7HATjaAYttlt3AI7EcV3p3
8ZEiHoiVrqrqeKIEJHDgVAM/6bCapdD3wU7iX7OehBOk/br4UCkxTL2rHxtO+hWKxtz/n3YPzhtt
ZYc+nsoW9gROdJU8g3EObn7B+X62RITpfB1CvWQ/DJPPwcngZT6uj5C0V/XxhEpjh4d+us2GoD++
Hj0AwaCjiIhqzO6dx2I8+BbrJwjPWZjDdNup9SO8pclge4kMpkS7R1q+pi1Jegi6pROcqJaFHfnn
W8orM3a+ssqkoDLFE3qE/BmmKEXD6qI/6XCqH8xM0AQF08LunT3rbg6FDpV4WQEoRlgDkrqk/HqF
BaCwpm5MKsAhqzRSJY74i83QCHtYgT9DwJIwpUDkwC6hNkqsELfUdJWIAPDHypKvbBLxZMbqbHXe
yhqzLVtXCG5bfLEBQZsL3oWJ6a7uFBYE70+fKmx15gcRRbuOpZzir8xV2hGKDDzzadcMYnyz1Sxs
Bta69LAWD2DEFwMP0s5vXlZkfgm7vsvyQZYXCKwsRncMUyr8yHHeBrUqWPJL7vbs+YtLzvfW36WV
BTkJHwkqX3Ci5QT080dSjoSY2AYNZwgsz2dUPUNo1CMeTfDq3usS56WK4GMMTQDKGSRzl22FzoeJ
Fx06oHXAXFkTNjKk5B4no4/lwLBqolzY6RKGBMmr/3XxPeHJyJt+aUDjYTVCoIdv8MKcdAKDaf/K
Z1F53JoInpOcFSEzXiVaEmNR634pA4ZiBZe2bhaNECOSZr9u81tu84mW81Ig4TPbJh/f/U+Kgl8a
Ongg5F9plajAldzltNN2aDozb08Ii8xWOJZP8GxzAOs9Qs+hX9uCbfH4eHhpeZYfK9h6jXn4NFPO
8VVgfVnegT613qwS4BJnEZhKpPL9xIHNme3DOc6cMk2BKbowvMurGn0J8L1VDZYgEdytjWHcKcPQ
I3dmSXACd2bSDbqk4J8lm8O5fQ0ZTWVAv0AR3xma1Oirtz/9rygyKHrxLF6Wwk0iVgRuse04fR8u
zZAu6IuzWdHBQb1/Xxkf2HOH7AVF6L1HsEBxRUr/fT+zI+1ybDMgxOSzD1Efm0VFzYN1G+9k0U3u
rw76Kmb62KYMcAjafqbtxqfkqj9a36KhgmIuqWNtBp8aNgKpsffpMJecRLasYQknJI4EHZaWhOXM
/6tgWWPhkSITmw4udhC1CuLIO3cuHm1C5TUaTykccccIlVVkZr5uzFDndNLmyrDCUOEHHR9ARBpS
uW9oSTtKXWft7ft7pN8BolFCIqyxo3Oa0dUivx5zgtMiVM2q3bwPpL70E2KAbdDojUCIABeh0Z/5
Cnh2h7tXjR/Gu61Me8u5Jo8Wx1N+y6GrQD662cSmj9zd3QKxWdrz7TmimfMQWdQE1uc31Xz72Hcl
K7bc/f9twzVCQYzQVesZ+OPTyjIhLwRpr2ilASgU3Dv6xlnpQhq1cniFHNH0CJL0F62g3ESSfEzo
I4th9TD7O2uloppNOe+j2JMzqHs6PM43rR+bZxE5SB03T66lGMf6tqoswZRJIMzBIa1vBQxC4ILP
pQ0PuTDulJ3Mxfxb/MHNMGXWL+hcn/auX9NJiqRJrUr0RlXto8TX1lordPPRp+1yd9jA47p0T9oF
XuGSk7BL0X/DI4MCrPos6SkqrF0nEgtANiTgsC7e5hO+rGp9TqhOPVoUDWer+Z8qHjhvvYkczObb
LmSM58UiGpn9fLZTnTTzQnAftfT+CAtt7wObg8696HBTcpCJJYzjBqGUgVezdiCzfw3/0m49swes
tngk+bU/36nGcEaVdwITlwprcIjrShO4KBauY+O9cBEcBJgTQ1SQogyNNdCCpKq0Y18y5jbnS86v
eO1eJIgVP/Wc8kbVg3hmHgH0yw4fBuRT3cVeTP3RlZDd7dEStEnA9kgjm4uQA1szwDDTTMdklY2p
HcJFrp9loYqrUwyRBUNNYFkW0LX8jnvmGPWrc+7PHq1a/Sd651EAVQk+/2sBSOqiJXDKjLDxYsAa
3X94jDsIHqOcE6Dq5nU8Nk+eC65v3EiR0u5TXxf2weQjpnJj4aqF/SG/89vVaJtrGadLTXuhtgUV
4YwTvXvlHFRvctY7HV60T0O7QK4e2bkTrJGZINBimcXeL2fgExvbn8iCtEjdl0hdPAhQ3/WKGm2Q
1rwGpmY9lLG1+EypLQxdJ4SHpEhWYRuw5SFu9TCrDZlQ3nO3B7S2dqbV554OJjJL7QluVWDJH4rc
7AVpPBsCkAB6DUoKxWdajIdDfj/+Oad0WTQbQl3uMUbe1Hu9q2vKBFkoH6oL9w5RBaDa9Y7sh4+m
gkbdmz1RcGUqlhVfUaXDrnbZU5UasL4HT8U0RPViQRgO4OEis7ctduW8h6Y0XtzX3l7uF68bBoVn
Bs6CnVGsYObkj/NCtjPHgBmPYCwvhP7GwWtX3Sc7e+Kd/9drfC28L9WGo3tjjw9O7ijBxotqTeOZ
wsooailD2o2Quk5hae9cylo7iePw/t+UsklHad3k/jv48/lBnv6ByWtszV6cCkxSiZAyrJJHVQBb
SLzinVAZ/PsSxEST4haNtzYINxOJnFlqt/CP3ZzNTaCUwltrCXhWnpj2jn1O6jHXLtSxB5D2GcRm
vlKFXxZuYp/QhZ0FfBMfzaW1wu+7mDRZVXnBmKvjFtYeS/z3xHfwO1WzgDgEblEkcRmsQLSNznye
1AC550Lkj9pTkqfoJKLS7cOgVfX3qzXMZjvGimr0mu4JdSaVkiFU90vQrn+lh7kNsrvjnU+iUSmU
X+iklc7qS4YHjjLFSPOQebwn1UwxQloYoysaE/vYTL2r3t5QFndeBGnPy6JJYbHV7OZaRV/N2W7f
ESVitWsh62JlXF8sYiV2TyjBFWnL49eHa/lMMRfdKvUDaRZ+i2aHxL9eSAC8YVUmU84kpIK8qtWb
t75xEP4LliP+jio3i8GHxS3C/YMVrUUyRcZNEF76RxQ5h6qOv1QU2eRDbyAthzB+yjceLKe5SIj0
cR77JxzgvF19uGPTHV3LSAWVro892aTCwW8jDmj+LhCZC6ORuQBpJv9f0YcadxR2xb4IUnFb8Qkm
vNYm+u3vtRMUoLqte3TysKHJQoS8IYqhdCMaFmgBufmOVTDRHDIBtA4N54wncRz5wRNROp3P+uU3
0TTzJDo9KoUA+NTz33vavPpIp0Br0Ntxem1nwBKBdtQqH6TQFvUxfYgvUyQCKKMn0F5v4y+e7yH6
nZEB19+w+jBrMGeXsuOPXMLUQ/CWBiwe5of3JK7ZjprGDewHscMWpnqFu/WWQ7Uv/hyzj99zr3Jf
/H5F19unZjrb6ZD9g9bAkI9QF3c8XLKSwedkLMhUVK9D5iSH/vI9RsRx8In0BgN9eMcZ1KyubIst
8PmKLlrGIWRIrvxnlrRRX5iRDg4xpvc92bGdicYe2aFH0en4uNn7qH9ItB7Ui1/bwVfq9V2uqM65
fiCwc8T9pJAwKweU7cR1+eqtRD65Pb0csMkwG4iHnX7guaOdiDrS7W8Lhplcmo3uwfKkI88CMfSz
nOEmyg64s79fiRfR1fbdP6oKnalsG0D5d86CgDz7tvXdVgJIh4aaiySpCpozVaZ0+0rQE91Wxn3B
0ypg0ynSyymjGqevgOWv6ss2ih2KWLOfojryiFmQ8A7L/9ICbLBnEwMu6fCvT0MWEysnV3aj3Gq8
ZzMmJR6A7RS/uhVQWlkLIVtpkxMj8e1AgvXJxx5k9V/pasytVHqylUrRsKHp7pjAVtaayCSY1MK3
eaoUpkExvilRamksa/pAG8tEvjK7FOoWOGrA9qrlXb2Kh1oEorredrmuYcub+gQhUnEmkQ8h3tn6
2WwytY+3ena38w+lg2oo5JTZGrfgQtKmvAinCNM76SXhrcS/cTqQSJ+WPTeR/PaPpKgHaBdOEuRD
5EMcHxlWL/2ID+oI/A40pU8tt9geZ89rlYIUBSGbsyU3MASFGObiBu+ifu/1TwE6/euOa0797vOh
85Sf2ouiGuaRjQDBBn/fI3qPth9NFLCx9o1G1riBFaqBzoQFHZYmWvknqGU+ZBLagIvsd6bTCamX
jQ1erNe+ZrMtq/y9qIqz+qCfBU2vlptKI+AItvOmKtOhA6kvZrVJqxlcQrmDvSyCUD6phB8XX8CR
1fwlVQf6F6S+4r4D530J2B5rHiB4MF9bAL35TWNVfBM6SZJRNOGCwz/7apXrM63KOLrTVTZrN6Xg
MYAIRbiJnd0vSvv+Q2P16wqsvt3KnR8dhITUhZFcXm+Y5aHSELlk8sJ3qCyiCe7cDsCawCdGYt+R
lqosAF4HsygxrbYh60mzVBKGkN0am1aA655u+ElzIeO+BK4N2E1L6lVmuVRRm5KALUghSvOwszv1
Ylmixw1EJxShy/yDqe3s+dtPrzxwKRO4Z4HWxNfdoSGOY6H3o+Ah6otwbK8U9y/hKe9ARn7PmOj6
UzzGwJ7wYo97DBlgisLSx9qXZs93RcxSujiyBwumu93pfPLOkjTkPcfY5JQr7jPXgXcfDphGysjR
h5U7rCHN5RKO42N42zstvJflgC46768pVxhpUJ3gJPcLICXYV4qRVZ/Oobjvb5O/aT2PwYosWAJ2
ETK/edqpn3fAubLKun5H7/BWGFIwZp7vEpPJmMQGkRDNQD4Bk8G/JaRNQVhn2f9xLRYnuv2P1Y6R
hbnmQMuY6z3ojQ+cHGwepfqitnpVgCUi51LPhf4neuOa9kiQE3UDb0DOBY6csU61osngu+7S4Xvf
pzY2xihNVmeqt+SgcprjZrnS3dlg9a7id3y/axDppKT8IZzTAbI0rDsGN4ZoL/KnKQx2qC1tZUs9
BpeQDh5UDC0xIajvNyWZqta57inRWUxnntFNHyvAZYWrp6y4FFLprvl2VYDgkJ1sIhDidxZJhPtI
shY4lXBHt6Mr5Gxj34leBNtua1anXh+rLiuVXQ6NRBdUJ0IAZTEIqefIL0YEDbwjRBYcp+kTI8u4
YSFzwNx+Oc9Vecv3X+mSAHDudgMGzd1oFCbxKygZdJ4IzPo4a4EnvQrc6g3YmFQsfJsu6uhggc89
uSVtZ8PGLR+D3ZumR88uhpP7uZMIRe5yoih1UTyK/dMnPJbWr9wOI8O5g/sFWoJZQQrsW02iVLwU
+EOLMCOU8vrUmdqK5oIcldU3O3uk9M3fnNkvj4ZhGPwp7K2h38xOXYyXj1ikofscoxaoXBWkKxjY
CJbNaPdBfUgxOIkV5viF7oQNAeo/vRZlDXElnz/nr/W/8Edtgq/efxVUhf5IZfuYr1dzx3+E2vHE
LGF75npAtfUXDoJdDQeyW75TCjP9opRzhWGYmCfti0MIdVb/qCX8iYEmbFjTvo1uuXtkYPbsWsZs
9VfszEad81kWZ6aOmzQcBUU8nhYzs/JxYoRZ215FMhJ1XmAQGG9U0zvkTbwKsvK8MRKNm3+iWbXb
KgsYZnFGuY0AcUnvsdLySZ3bVZJe9orozULqFOw6YFMMCaBgRkrG3Nz0cSM0pIRI6Ym35RWltk8k
o85oahU2dmBXwlQAf77zjHjbeYQaR8ZE4QL+eGVWoeKI7SQmrQd8ACy0tNweaxt1IQ/RwYS67aFA
xkeR3jpomdBMXzdF/Z3y/8M9OV32RId6qSBgchfFW96p+XCdEGHXwtkTgsk88d0R79hBz9ZK2T+4
rJhtBeYPKHQDcNAj38B5yYYqSAPIzLyL9RPlITm3/41EJBTNUqhYHgQXs5GpfcvEZo7GfLNC7MBT
6D/ZomyCWzlEWUU8ZDrHhABCjkCMpeqyG26EbSeVELO0UGvJLeVJW2wNshexGLDdonv9lPS/neTI
xPHYVK+2CgB+423syTEXk8jcNqsvtRDs+E2gpR4H+6UkQSiBDBSXtMhKBVcjLg2eL9fljVUIfdt3
1Aet+m6KOYIVv7DLpYT7xqkWcIBJ9tiuc8a45ELU7kdht2g+Eunt6ZFXeueZdXpBu/HmwLZgQpSA
gNESDtnd0BlNMlu2hEesk8y0s5aDSeAd5XNgu4F+5KG9538lac3ORvf0Xjz/ooyP6C2mrrcmSbE2
SX+FYCOC9HRlUY3zskrS6957HkUwdeIOLkC5fgYhuKTjHk7TKJ9TcA+5Hwy4fjyajW1aGMg7XTfs
2FtLHuOHKrzV6ycDPdsPP/r643e6ijyBPT1Em1UsagNm4w8D8fWIEe9yyYDnabP2aoPL9Shh5Rc7
EoktAYeGX2TG8/Uvwk6ezeqfpB30PhLggrbaFKIv6pzvr5mBCif6NExKdtE9BdqPmS6lPldbQI4s
ZMmhJcFfej8ISxO8mwELxznn9Niqr2Xd4oKlTHaU0zJdZ5aGNJFv1TUpAs3+lRCyxsWIRq6UmRy1
IIebCtmErqn+/0Z1FSBvkLqwLtlFU1h6FO2n9Aka9zrYsA7m/BeChjpndp12GSjDdlsXi2OoChHA
nnLrMs08TcTwtI9Re0Tz8nq3grM0EvTzRKdbGiMgONnyHFeEMcXz5WoolNzrW0tEeH8xjtrNKsUD
QIVQ4cqNWIIx+2oYP7APzRELIxdNslgIn78Rc6ftM/jDYpnjZY8DUec1WA6DtT1Tv05EEn/plO5u
8/Gx49PlM1HBYORMpeDpkQHjoI5cYYSAyR9s0cuxQ43LmveJiCWpq8kqzlLGkOtGUY9ZpAv6BExW
cVKEgFpew7YSXa4XmUMyxg6UdSJBfxPcKsimK40pgeWRhcwnsnVUWbMSxYK6uMgpelge2aQ8FZAS
JNg5DS2OuhGHkbqDoQq49/nCkaDyOwKI9pE6ZGx0ul4Isn0rd6QA825afIhe/rqskIZf2FOFQm7I
Ap/c4I8BQi3A8i/ysXjXm/5Of+O1o9u0mkVT1WzTYyyw328QiipPyoLs+iecov7Jjm1HhPK3oeWy
nMjbXZeeF72eF79qFsA/crDpg2L2Q0LRk6vBHCSExmuxV45BSXT3lC4K4APZCNGF72Bs6+kX9GUI
K7gn0s5EnNHadkxsKEWtT7as4ODQy1PhVDDsDGIzxNIOUPYnSuXvtq4IJGUNa3NnlaGX5c3KZf9y
eXHg+h0X8P1BQ0tx+N5+b8OG1ZWGpTjZ3gLkEYvgySUsfUjuDC+XjE4ZOqVtKY52tLBANNxN8prd
Jo6lP4/pga9+IPbWCJ9UIDcH8ZUIS1aTkWc9Y7cgZ/fSI1OTbA2Vh72vwtSYjGI6VT0gbusCqrh8
u9oTSarAKMzZsppRYPBJ1bDUvLpz2Qps7jrz+JPmQonoyPpJ77eHJ760rKhH8cIKk7azaZeCwRKo
12cwTLohL8Fzv+rkvVXwu86iV15qTBEUsJRYP/i4hRwmXcTEMqfH34fBVoFrOI061YyhaGXa4sDi
VPHk45RGEp1cToVbqHW9fFPGI/uWVSqt+b9Vu56KxubflxIw706bupqXkpARlsEYEtqoeJDY0MQI
TTRnX0C3bvXv8yz9e9NrSAuh74aRkK4/RFRqrtZy2tpYqqtyl1tvog6JJzx9gnxF+MNOkq9zPeuq
CCldUwiFAWvftULohzvNH6oH2dK9bBg1Tn6Tm/cILqWTllWTvalGXldvMsa8CygKaTItHmgBjV1i
gcPCA2hP9Weo5UwzC2IHHjiSbdpMI17OOrSeOsd5O7QVKZa1lHYSvV0LgDgFtElJVsNfDWhtAzUQ
pe+tUrLCUb3xXNxaf5vDWZybl3J4WcuYDV7mMYjWND2tlZPPTOtoVz7FH8xoeJNl02nJ/ezA9QA7
jHw9zhpxzvtJ/l+NvkEAcZ0m/cW59MBU14dsH1FZR4xk6mMBvboZ3EUvNkK5h9qnbLZsmzAaWh1p
ZZcSzoyyISo3MwBI8gQ/FYQCQwO63Nmz2WSrde2K8r5N0a2aPPizMY+/6ph9/OOdp49mOcTWZkED
Ow9dHZqNPo4jLodD9X+Zz79lx1IIuX1TvKTzzn9x4S3CNtKLtAChNKD7E4N4N3ewr1xI66TbehqK
g7nlXP25uqs9ISa9KCo3MD36iDOSzc8RaAGNBaUJIuJF/gqeOKkmR4lpFJIkLLBLLxIh0KXkXXo+
JR3117Dt2uf084cwWhwa7AiUXpLnhLN/Fw7l18jnJ/9VskDPfYh1WbgZkjo5hMzi6Op88SbcZm38
blUqPAB15kTV/HKWGYhhDNl4VEIr+CA0XcMjGQKFYs5NciefbuK6q+qPvsrrq7Ssk8lUFyG2zEiV
vcCMnsH/xJT22RptQlmdnoQ2gs+359Mt30Ku1WVs7Fmx2LvETQtrHuT2vshXwiZB6Q5wu3Nq91cV
cpKYIPY7hxF3qWPvTCnWHcgimoiFcOk8itwFwN9g0b7eEkUazFn7T21py6PE9lAdT0npzntzyyFx
1mEwYTV9Pdh0BQTQtHSZJNQct0R48nWhzSVmE6+enIdaef+Z7pJ/sC8ZumwVlI4vHCROkITnKZdX
sED3df0+9XpopPgtJjQyGurbcpDwCcC9CU1KwuYSp+XeCNbYD9jKt244cAaEF5YUXqVY2DBTTid0
reuDc24xaoxTEfnFSuOAEtYQo3mCdW0wiImU/BtO9Ne3KnD4VyL7LQ+qoXwL2A1RLYaB2Vyg1He4
/kFmXYFXis6mfHIngWtTm7tgQ0H+ZH4PhY6lM2SDGGmZIWawr2QbZFDsEeuc4YhDmXERboNc5Gil
es9lYQcml+6DMaUrIc/fBnnBtSp4pzSlcQvN5EWC8el6GmZyzY4DRdhq8DZSnyAHYgqc/w1TBi8S
JGLGa8hZaX1Hwo1cw9NA0oBEDmzrieujTGTN9hIXyTCHmXArliA2zTyjiFofnx6wal9z+0AQZT6N
GycKERCea7vtFS6HUAwTYa4ZkJ+DBmWlbOmrb/ihpwLcBYX7dP1ullyuKdncQkdalkzTTdmMEc58
G0XPUP+scQTRUJSmTxHcy+Q2L9UIpKvEBOSgo61aifLT3UCkjkkuXZUx7+oYXaPHG9IyA/DgbKTX
5jQ69ybdFplenm7zCT6ZmYNT2H+LNOVvFVjZv/zYHodYDfIAZIrV2dd7i76Tv78PrYBDvYSjvtVZ
J+ncaK+uzNz3XNERqp4U40UlvmXDFIa/+oaAGTz5QgPBRGmm7DRQwhlpOQqA9jddqnTt+X/KVx5w
ZOSVd4euIzfsOEZB+T1CYPADwbO2m6vYMxazXrStrjJ1V7CpqOlWDQ2wF9LX1bXn7xVDJdTyW+tS
99bgvf+fKTMIjSexMUXDtlobwcA/T+cUxZ4/tuNPXdz90CyRUgxCpJsbrEibvJ8vEQIyVPvDB0AK
ptHBIoxWmHKj+mOu0VR7SFvnXm+W/kHbQGnfOvnDWsnq3BucAgo0X3chYFh2EbTd8dez3IGhrSIC
q5v/iZddiePnjMP7e+I/nfY5D2vu66o35EZ3PSQzkcxOpD95Qq7aS3lq7w8z+MKoPsKdedHJS2Ae
ObuEUX8wt6o/cTAExXbVIDbFkGaQpbeS7/SC9RKUlqFKhWJBPusLTNT+vELgjURF4MP0ssBf6ybH
qN2Fwb4TOY9EL4dnt0wK8bGljO5Y6QIU8qUiMEiuUL4Io6wKdkoxngGdz4KvW1ecvL/3++l2Wg+1
I6mh2pCKFYX7d4UZG6BIxvMEXf9x3ETLRK6VgpRG1WX4P7HP1Ag7lOi6ckB/NAdF4erUPqzSk+S5
FGVm2nF1YndA/TACVJtrxwTJeAx4rrWyJNEkDgSdVAO0J9Ns5/bwL011GM4j0S8S6T/4uxwXq1pB
mHxvU9VCwVo7xHXfZX+ZsbHYi6xTfHW+K6ZclhpbzpD9zauTxOtUvticd5D1nv4ctWX9FrAzrw2a
NR09891c41sP8P4xEQiRJzc//3E0EeumdJq16T3E0n67P8uLqdRquOuB36+LG8bwbedc9nrFSEH0
HUO2s5FYQZZaZW+S9iHsx2jORxHQbTL9C8cEBG0k6CHsKmHR9E6IiI/mpFQRfzJDFITIYyyLpur5
wdHzknRHRF88DYyYPxAxY/npNycihALr8neOf1bPlHfhqh/QFwdQ7qtMlf3wNwj4DvdgMCuHzcsi
VLsBd+O8JdI3YsI4D/auLbxyf07YavxROIKTg8J0tj8JcXTV5PZr1Z+O1iBY2DBkHoZZao7qrok8
NTxS/FJEnhXiwYp4heeQqEyVtKtAtlIWeCXRfKENZWypHH6Xbiqd3Kq3saXl3C3ouUQg5Zyi1iQ8
whktMFtLLpl9dIb5fPqZw3onIizqYRFH3n6NfppPl62Gg6HsNALPky3qHq/l3hk6Msr/aWi7JrxS
ppS3sfYNQmF6H6LYlWefH/mauDa0/S6URGfTYGwbcaAKdDv377RyanSX0YRmzb8Q5alv9rG+NmEn
7XId/226kacr1ME79+835Rmz/GWWJUANQ+82gNBHwve54kY+zMS0AkRbY77jyIhDM457YiyYxlPf
Ek5qAM5fDJzvOjjlUXlnGnaAkmmpCl4iMIgyAntyRJOS8EmPCCXyIVOcp1ZrqnzDZiKU06BwEtBM
Y9cRH2ZgmBvCoVdv8LWIbaiUhs9l5qI3oANBca+gWZX2tfBWUIcFHBqbpMQuys+sgwZQotZolOap
0h4SNDtAbGVGaZOhn4y+HIF0NQ9jxfjsUwVHRlrW3CsR0fs5waAus74OQQRw2D5iKphaxnA/2qYb
ZEz0umQm9V3ksupMTmhx9Ts0YV1P+DXW4xSFhB6FaNVuOsvnwbw0N9hiYTRS7BIh18xgD3QZ+TBv
LuDThqZ9A57TMzfVWxsIkYRypk4XyntAHbfl3Qp4e7BuWGwniMSg4Wsjxhs5lYjoSSndIMOiXszK
h1MmqazbidqueokYjq4AaASbVJoz5Rf311Ykhmdj6WsBSqgKql28MC2UIvSMbHqx/MoHmiUDMtJS
xzfa4LTu86yI63rN+8SKxMH1NOiOYxmbFK9mpDgMbZK0xcn3cR8x3STY2NNeGf9bwQW78e8o7/nJ
sn6NMozeWCTKTSJLXptEbHjS3j+qlX9U1j1s+kv6wIznYi58Y9sYo+U7bctN9FsAV2FEiVPah+va
Qd+M16RJal7U2nPXHWTv89UmShHDRwzI1k2nDD+pg/QT6/Tl+yoqzrIC1DDY0vKsLt6LG9h1IEfs
k5er8n0gmvbGWZqxo1zgaOYajHrsgXibz5bJfnDr6Dd+98fze9XwRGIeapNBDFob0eoFMq1ZMFiJ
BGvJEBTBCfXVzUULLk5ijc3P6AYYhnLwTxplHCU+97nUX5mRb4F8gL3b5HMXW6KKtaflBFKyWyRj
rnMMAawkMF/1jg5dNrL+RdvtSeXyrLSOHXI5kWGJP2lYI0BhGjRSm7s6QokZQpbMXScud7cztTBB
vK80o/gX8VzXxysOuatkOmdZRCakYCyk/s4+mCfb2TgoYnbsyif1bmArILBYLgE+UrwCeCkyeKI2
ShskhJCHGkq/hBbwMyhZ3IT3XgP2XvCwq4PcRq7+KSHur1kcpL+R1mhbXXjM1QKh15Zo/1D/RooQ
MRQXP6VyemPFbbofnCO64zCQvCNjK0zI939K/nI8+0+EFbpD92MIE1cpfe9ZT20q/Xm+Jzk4sL+H
R2Tnw8MnSnvG0jUmZTztmhTA81mk1do0egNdkVDrJMInw+lnIfQUIK8Q8OK0tCptfwcVJ9EyrQiG
nmbTJ6CT0RxvA85SlbOYDKxADQIp+cuhEI2aD2MVgpCPIMaKp/O42DfCQj/4gNGLIRwPBSowNTp5
r/UA4q6Xy8+jDMoglvd8eSf/iVilc5emfKePQoCbsj+w1N+lt2OcsL5cbI5VikUtTaq14QWwZh5y
zXrNc5HBBG5Xw4EUEvabAhkHGqg5TquPzeTavyfEIt138KIquglF+Za17uURShEIEY4ItwDxx0+u
xc379IRYjpEOlHadGXy5croojLej2SjOB8Uk6J6bvQUm/5DDFPP67Jf7AVR66WtXqp2hn1f9sdQh
hbypQ2yI/MIh0zYUvoAu5jGxqkw2Vy0Y0ip2hBvA43pC4Y6IpSLwSUGpgP5nbbuL8uYqKSWae34N
Yf3Kv94Zqlhk0Z7XRehlM6TpFkBgwjS4eHr+l/dQu/oB90XSdKLorIBfOykJMhZyoiJFIdgyyKGV
35+U0O5LPN9qfkfG+hn4UzrBIAlnkKVtpolJZzGS6l7hgIvKGkqfV1rUHA16+DzrH3IVPkSHdEHM
yNBo6+E61ZfxYTxs51yDcxkf6FJxOMfdUC8nYYpnpFT6uAPgUjm5bqz5CXZ/FnHPwB5SOSZHPhBq
kRoA3EhLH+jdt9XptAAYgEpe/Gb2NBEmFnvaRJOf78yYU8UJUBFkCwdXfitI9h5hK82aTPxpOoux
8jixEopMLEvlgVLZXZThjkPbXfgQNX7w8KyXZUGBhLYgMqeaTOpvtKf0rWF5+VMM8nAI9pJHPRMp
/gLCpF6yijRO7slKsKErDf3OtluTPGv2RdiGneLDvpVujXE033qJrLIkbg+M3f1xE3+ZEmM1v0+8
c7T+KK29ks7KUefQCQzMELl/8tP53wYy/gpKDyK+SUWqjxTAEWP8iUwBPihbqKkj+LHo/QLhkR1j
NbBDdfiX9QEQU98HKKJSmWTDvEpSx1QbmlSX76uKVm0WaPxQeVvdaqBBsGOIJ7SZixP0ezMK5C7f
eZfZ2KWN0oAyBQjzdXnJ6Wxt3Krb8SI66dGDVvRjOFsKkydkShX57BNawVRFeXthaV4FZ6exw/GZ
75IsxFSx0FUMyAGSTQIAdGkDXgWIGQHUadWE0JS593AFoMCUmqJGKsaWIytibxEIj3keUDyGm57H
cTSJv+z96zncZNj4brgTxcooCrefUA/sMEpN2UjEbd2pK1C/5Y+ua+bLU+Knrb8STcWNNoLcQD3P
jLxqo/0On2HF/pud5EngwN7sdtH0+nBct5SAnAd9frOhfLPYv0k2OTZJwv9/+SzWiPgVmVdqzRJ9
Op3lSAqtnQbDCjBSG5GT0QvT1X2ty0vQa2MKr0KP6O4/dQuI3f87nbGisljfRz+/2b6p002mrZcl
3XEEfvtCua468Zamgi9SSM/gVGVgsctAcxNT5LaozUzJ8iD/fJVNuR95nyARCvnDMVSj+oYYiNSM
loYuzKw4HNnYr0GVPD7e37jb2SoAyxwGO/dkqnYmaHkeWt5F4mhiwgSQWnE/67OPITN/4YdJVfU3
PVPhFC2qZiWH1PlS1Hz11z/tZxznPlFqHVOGZGVCXn66ciXi45N/tHATyMymxOsX7y7scEyh3huU
2ro4N3aOnwDtAa17JU4EpNxlk3YNJ6XLH6ROF2q2q+IOkHyQx2/52jG4tH6PrEQ7rPeaCJwv9rrA
nZwQrSy7obuHDCoA/iWdyYwghTPOvoNyXhDdqjFi76Epbzf+CIvIPOXJZIayVX5gKREI4Nxv0AaJ
dVIK0+A2/aexWh9h06YM2xN6fcUacMtGn3oNz/76c+r5BK+2ByXBMhMlv/3u7QY2nDeasN5Ucwep
RoNqLiZBEgVpP3Cz2me8hjtF1LYiKh0in8HBE4r8k6My0vZbF+g2KG//OI4idlnIb+4GbtWUSX2F
W/VpggzfZfP1gnbbjfpAImQ8dP2GbYUv2pj9lDhz/wDQVR8ZfdjwZYe/AtfoJhBir5wqErKf4ern
Ld8Gjo/08eQ1YIWYx5g3gJ2kYnmUgL3MBhm1/KBv609v2JPShBBxTFHB2g3SN8VzkYRTcs+eYur0
T0n4iBNe+bOue3BI9Q+O7cXVSrgyLof+LVIejIjVPDXt9cYEqMYi+MzyX+6UWX9kD2e7Yl5HUhN/
222renQE/8tmTHJrjd2UqI8RvhXvE3fybYH0ibrCydcpb4Wc2K+zzCm+P3QbxAtmVQQB9LSNbXMs
fbZxgAELhHW4qcHbJaTtDpn33FNbZU2ojmmBBYL5+v/RdgYLkuB0o6ChPtrVCXQV+FDv1aP2WCSU
8saXcOLTAdkCTMXeMPzcwyAajg5ywKVBMR6BbB+MfNK7QAscfopt2+j7PTHKDv9ZNHbOXS3mLxDn
3BUkfBN433aMYfUvRTJLACVmFShoiLqTkA8zvAEoIa59yVhwzp7yb+6APC5nBxrmLrobajAeSGZQ
lrTJp8xCiclRKbMLtcMDrAxvVpx0Dlo13ZqVSwVs18o+44iUP56bE9BfKQjAy2t3ZjjN65/EB1fi
YOpXqiKduyxs2UYeobMLSfN4uGrhR2I5cnVubJS5ekACZq6+gv8uMidd7b6OSWXlTaJmAihUY/Ix
yi8TndsVH02lJvgMNDZaTU66/nJD9tOiet5vofSOjxuBeRrexLSoSgfn9znnCdRLp3r5Ac210btM
/ZdQneRbiUyzW8R9INxzvaRIueu3AEhrL3xiqrEuZwlQjJ3v92RNl2EfrXQ3gNHOT3TGto3Exjqv
tm3FoRTKcoGhoVsQQAgpzUtR44e4zlDrjFr0YcoEAEm/hV0UaLGtj+mzUwnECH42EP2kemIRXVAs
HtJKL9EJyB0oT00i1bfLCNw1cQOACvHQkNqBEtPp1TOo5tQarF/EdKTEQO0e0WYjiF+zU9AnC9yx
dkbfd7S8QUv6slHxd2hK069zTIDUYXoE5P9SbY/RyoxY/z4IcDGpmSzMR6BwZoSBbyXR8lhM4cqR
YRKkOT9iHLgSu810SGgfFpPhzdgR0SbcmW2k5X37K3q1xx4/TyvQshz4z+74ar+nXEAZe3J7tFw0
Wh1+rIyLBXG3WP9XqDmehuVris0QqQd9KJvOtzuTIZIrLynuZGEwAD/c9pZ1bN5Q/7mBLB/eD0L8
N1UZe1pOyoDzAnsDB8iDpCc7VPX1pAjcwWy1eylkLnnWPa0pZoAFDcfO0lTyYxC2YOsUMuiEwtUe
7NHa6xOq7bX6sbI+n3fNSh+vyUUd6NC86mTbRUpnRbrnX3WHR1XrRozCWNneHGLDpj8NO8r1X7t1
zMgxEuNM5sJlxUHJewycyVaHm2/SMKCC+wqEdIQGXIsb+m9XNFTg7dpOinICti6zACQzgDVfHb9V
7NVyaYQy2oDXSMTrt3AD5CpnZgthdx3Qswp8BQRfM+roMOI5nktaY9HetWPQNCzsquha/Ftcn8oC
vYgoGxRFo3finoiqYjmlVAOHysz/JYUk9MPMQ+SxajMYwxC6b1D5WabZZcskyQc8UbUsQHMGuzkC
mkL/jzm/Im+ZJbd1IKiQseFTLAeNM44ft9wD/k1QNjUYTV/quPrmpyzz0LlHyGxwezoCEyLfomyU
+9d+BFhpXvfqk9RkMZbWsF8gioXBIv23KJ0te3OVTV9AusohyTnlzIsg+sqFntGBL2WZANJ4P+/f
+87XScL288EjfV515etY8QKHANX7h97UdmAWsHm6exGxaHUg6PUSAUDCqQJLVX9U9tOUi3p0T9Zr
tghIHvcCrHlM1XoY+eVglfoc7+zDepWa1iAH2mfkoR9891uAwi1nMcVd+mMui1n5qdyHYQYrpIOK
aIwMNtNKqbT/9wmeLR8HDdjdK7QyKgkfpQQdl4K+jSTf4UXFQa2CV1F55wxSeyt70RjPQDEqA2BH
uU50EKEEH7y/hw36qkdy+CHjMuBacEBPKR3c4L7aGJ4W5IgMB31hOsTx3w5GjHObm+iYPLH6bxTi
zy2Hq7jKhcU/UYoBD7KZtNOH5VNYDOQNY5lwPIx4wZuWuz4XR3IcaS4SqiBewT5qS/QtTivwufDx
6YNk8AULcD2zQWYrtePxyYt+SimrZgAsU/topHCxI01GjzGdkmO2yWrFnzDi4wYEPlH+3cEBYXCw
vbrsGjb6PxIUJMu+dxIHTb5oT4qAcEETK9eLuUIFVkU9moZVNy2/tyc1DtQIBhkPq8byiwYLVKo0
1oJU6eyBPtM3Xg3FnzXPwWQqI9XEQmem2KLmzXXTtjsJTdBo/mFwKVCroFf3u9WinRsGGKF4R9CC
Xd0NV4+1A3S0F2iQRD/8yWoV0yVEbU6aX5VmOnolZelrn3WL7qdUCGedtbzotEwwrvMltLGzkq/J
DQGjPxfZZzRjhzs5MDbhXdvmVEp0rYZIHy1Lrn6bS2GoOhrhUw6pjVSqj5jkQwAVdVwU45sDDK0x
P7veUsNDQC5Pkihm55+P5NSScUhTplg6guJKZvhTPGZWpRKPLRKe+iXco2Onj4MySbCmNb2bll13
nDuuGOHzbzaRhME+tzi6erMjGEe2prlSYrmmML9sw1AVckqtJ+cFxpq5sRax3j++S/SZDXGRy1t7
JasIG21E4A2c7RpyjupFxFh9jCf0evSWzApQY+QG9zP2KnwlbRKbfX/eYQABeX/GowFbwrKj7gwb
McG+ZbB1O1i+MdHmS/2GHTuB4B6CovBu98Ll90U+d/MUHRqQ5yHHY5a0AXcPgLxltykm+JT6LLmT
U8JHUiTrW8MXOs9PyB5ihd0OLldMkDmx9Gp1zQfWFJOnF0sJMkzN+mHXwf+8/t6Yeq+GEplhcPQF
996/Hj5c2l5/4WbLepdJkY6BjR1/rt3/SN/2Sj1o4Ik5R+GRL4UDIHezYFGU3wmoY/QQo4mTVlXl
lasedLX+MvqxkfXZwOiV8nx4nSVgvxRrJ9bfwQE74yozfikXSJwLa9w3OKxIdUJdd3j/njSBP05+
FD37aOSYAKkp8OP2j1aMskGpECQ9Wy+RJKXVlORvDdVccrCR4vV24BSRziD0yYIH3ZY32uKjcBud
06ZhNcz3Wvn26C8k7AhW/2nrn1qtdRHmDh67McQ11SZkOOOZ6XzLAHLDASCc0LA+V/8kFP90BqlV
0EJKX/+R0/lr6r8lzrVhl/bMV0sZpFyv4O9unGJNTo30lkKBRAW0KIKTFiy4Jm7dYL25q1qbHsLm
j81eY5HGf3ppBwSEA2sqWF3o59XXXWl+r+3Y86eP1hybcLmTkZ3xFWxHzEhU60pozE8m+EapReR5
NCCr2c1fkU0rmRFIPLGYL2zxPaNvJ3P6F5GaHBZqyabAUN11SsNPEc5n9v8/sTKufURFqOpr73Jy
z6piieyepWbDLXX3vdIpPje4sDVp064qD37yGJAgCf6g7fnhaFSmey+fVTc4/CrC2jtHicy6v1+G
r1ddHHyc2hVgnVho417XYTQ3lKrgVr55+DQ4obPyNBFB1g1HEU4zHO+n3HHOS7cNOYhRuPbdCmNs
VWbVAaV7SDK7/y9xUh/CT5z+576IPXJobN0hfzH1CEw9g7Sq4/GTNT7tKRTT2sw0HtH2GDIx0oyp
DMW5PeIYj5txp+y+cy3T6t67PLBKP31ZIvd7HIHAd8BwV0LPD+JO9DEPJcIvtCRsLOq9n2UVlo7R
iwkbjetdCCbkuelghZSBycyICPamIiPowbnNm3UMAc5g2/5r8CqXhm+L5bkvV9XZ2Om//W2ewtEs
NzujBTtCfZQJrdz2cGCx58scj2yaN5t15kTmzsVWkfZZF7+9wlb1Anyjs+Ge4uw+6XbMMYCfA2b8
LsbvSQYKWmXj0leHh/+rDq1PdxA6bDwF7e+lziR/k6qOGLYrC7x+B/huVIzekfQOYG7bp6NZ/9g/
2/5zoYQZ39yhdwqV6sWAVnfG5L3zjuO/WlILIs1hJtChcC6YA3c2WEyUJNF+V/qHUZDrdIImp8BB
Qt3h5sWM8dCNb/rBBbhRCirXL6HjZIi1IjobiU13AEdYzRB0/+zhsjsZOyB8dncrXd5EWb15ugdL
qFuoVpgdl3utRlSG5LChv5lGDpAV+Zt8bGHS736tPc3lFwsLp9V4rzujxYU+Mvxc9kRU9Uwm/eyP
IiL1E7UycQvfFrKGN8rVzloZ+GOpNSPu84cpX/aUOoLcINo7v0rViYGnEJQD5LmPZ8S3XhLKYed5
G8FDuKbSPliXS0aSqpWbPJPr6LdgY3bC+o597SYo7Dlll0CW6TLy3mKtaGto/d6D4ehZIJVHRjcb
EB/x9r9eWWEiqJhlhlvb+L8ssvD+OFv+0tfIZCrjUQrauVTmeYy8w2pGhNMo29m5pF0SqeVIfN/3
xijaDDKS6+l4bjAEHnWcGyHVONAdijpcZv6Wy0twVtKqv3KQgHzTBfRP3a6XYu2b6VIelYgqiV8n
CRpZGgJH2ReC75qP8D6v+oiX2A03C8XsXt+xDJfhs0II7tg9rZVU36eT/9nPgG/gZnO856FcHbSS
RFotqOMvj1p8SpFBKyyMQ3zMKi8m9sZWW92pDbrivDpPyUAwaezii9n+W3Dhwc9SuDcSJq+mhOzQ
X5DpnC+XEsfesBkkACJKC1kLAfqWTihlHJYNDQNz7XzDGCt/VHVeoDmD2UZLYhahNc5q/fqOFKWt
t1mraaf5nRCENY4+abFOxWj3l5X0l6fT8wpzM0OGf2hlS9Ko9qr1U6v+IX9gz8Z9ALDw44ak0NGM
5icHOdscJKfBmpAXX1j4PVxyDFY9XbrLXXRGcDM9Ud18p2dcIaLaEXcl5wy9uvKEZ31Aafe1uLxr
175ZpuXqv5V8GEdykR74BWX1um7w+AYR6QBwMzUAsVvKxv+Ztjy7jqfYN/1mwgqoWuaBIWNPPbyc
ndKX4P/vn30yNBCTrEr7BQnsNST8k6m0hiD6UjA2g6gLG13kbieeNQTK5F9xhcQizHgYbVj6lovH
rpadfe2m26sfeiZwhBzR8hrvh6d4TxDRDbjdJDDH/FmNZcjOuPByTHxNiwu7MN0hF9B3VIQVm8zv
saKT2ilYzvafy5zwwMBH+qxYB8SHg77YO4mksjEoDc9pT5UzBv35Q21NzRoZ9yH++UufpZPbwfvN
E4sin1wq9SgRkYc7LmDBYWodH4+OallC8WrUYjf6upWmKaEWC3Yn+67Kh1hYr9eP10VHQC8OnGfh
kjlksOGFkBBxXKFr4WdtYkJsFYPHFewHTS9hNO+R35Dc+GpswMdnfH+PIL5CjkgjMdssTFYcaLI/
tLvtRHmWXj04CgIScOBh0UdWgsDPJ8yDLl5LilQ2qd8eXZqD4AYV9r9Iiscy4iZg7+Q86V2XeIep
sNUA0dNdgVLN/d6qfqplqLCSgWIyEJuvERWod42VuY7FfTSadTxtFhbewb29+gVgzyyRaSbQ4nbN
kjlgZdOM0oV/KfVJAPnBbcxMnS3fnKmPr3arG4DU9POFycLaKr4gxd9/F7N4a2369dso5m9EGG3c
RqZvpk0w21lBtm5jNhE5lswCaOL6RIA4P4M8hAEIEN4mDU5BuvUsp/6lwOvmysNkICpR/Ui1gf2E
m96iVty22S7gxt6WtCPVe1XyiLAXxaBw0I9Bco6A6KFB4tgUED9MhzondQnVUiycuvkIkHux715V
W/pjeTN3VeOkISj71OTdbOTXhWl75Urhecf7eFZLs/yN1L1KWLM/v37uPEXEVrNtjDOOLQcmUybq
081Jpls/QU9V38H5FhCKnzevsZmFqseijRX6yNen4eF/y96Wn3+CjTiReIttUSS+nxQx71X1nJAY
jT+cr2S1DADR1LCBkD0faU49xrhqqX7BCJVJ5oj238qJBumgjMp6YZRAOCWOJW6B36HKDE4pj+Ey
Po/0LxIV/BWsiFIlB4hO2p2dAop3FhpRP1tzGYHJ7j4sU7KY/oyPHCYO352IN1YEDH+wZP6Yz1zu
9yl1IkSo4QXsPjgquAcw1VjN4O5DbwqC9TyV/EwWr6y6iJWx4CW93f6HdGgjLejIZMXMQDUnvffa
tF1pJsqzDsaDsELUgpLnUjqbLmFAlMVHfWPUfcn02cqqO7Xv1j2oqij3MUpdNmtliBu9Dlhgp6U1
MROK36oVRH/41yGYiSCvSEuAVwTlDsiGy/1wKqPwXlJJ6iD+0y+Pplwfnk0Aypen1ReIHSKKs48Y
4j1ugJpGvBZE+hgDnkpcqyERRc7esJ6W9lz7hIAYWeWVR/jK3OgV+eVeXNHj+F9Rsu6VHE6aTQR+
Y8qnylBO7nokyNN8Hl8yKTyMqzLfaTJxxoty6IiJGsH75bGz8/J/YXhauk01JWcrlQsLpPQSKHi/
S8AOJmfPePFS4KWOlLsx5/vCF3nu+E/xLHYIVGgf2Vdjk60/FRiAIrpfFxxLvqT4Bzra2vGK5BkN
jWFGE5SJhKsiRF2Ef+oLVMpQ+zN/Npv1P4LeKLKI1QRjaf0dDdYF+nzDcSnRUnSexZb1/bAwZ69f
fJ4RIuf8mRA9fSFlvlENexSqaBM4An2E5z9bn9iA/zE5Q/ifEJHVDvW0n2XZKk7y9a/RhIf3Ai9h
knltQgDaEj/FyWpR+3FJtvfRMN9sfxTKmNgUJyDCsXeb0R+MZStTbtg5+VUfVZ1NsRtR1ETj/A1n
echrjAc1Fqv/R0e4MxsYubH8qFLe1v+EHRNggPY0Wd0gNZa3OfCJERhkMcU7eveL/VKH+jmQoZIt
Ri7ss9zpDmu431V0N5hpVFmHc0u/KXNd+htuLRxZWHAeYWJRmjw0WZTsLd5nilr9G1tuMA2jlwGx
AtW3Xk7kgc5ZcqRUkglnusyi84FGlfsFD85WX6sh07x5wQqxO3MvT3hijgrBda4n8gRJ5Cd9V6TL
2C9QAwuowkAzYU50dIjjPQs1BD+Kctk6KIBp8wx1R4x3jqWFWIuMO5y+oA/4x1he3z2b/390kR5Y
D64ErssrfqRcG6QklEo64O8u27Qp4GNiyhtd6aExRs6iop0HOzTsQqe+mtA08didKQePzK00dACx
zRtRvJrGwd8L/no9H6XfxK8yizNu7ZCaCJBvrwvTu7JzEvrza+h4wHqGnyERgOlRfrgDkjg8TVWu
rmpQelJ7OYpGtnJUAIKbIM2kPyczuZ/uXuJIUma7E6RosRhg30pOfJ/wBQjrx6wVIRQ8nS4/cOTH
t1VDYWQNLfHzrwkdjFB7Q1s4WG/F4WAt0P/j3CW7v6OPrh1wB6mp78N40MSskLKT4p3jTOVTo7xR
yzbZDUEfnOWIhzrjG4m2yg0VED+nUlTqa2ExVDsFkms1pvOkNuJpoFyjbTPOvg4gAYkh+kD+IXcO
gAaxuUkcx+AAevoGld3nPRIBKR5HWKckqBQdjvuWa95jbeZFXCO4hJA5krYO4AOPTiVH9qruhf7P
PBEm2Grdtzgge/VoUF+4R292s5Za+20FrPSSSkaXupFuk24e1+RMkdn3dHhuOAPnIw64hJouIMY3
iZwYvj9NBIr73YFWLXJ91JGlsyNSBp3qzATSZTWV7NvE880fC4xDDaMvhfnPvIh6UVAfRUR3QtmA
rZX8VL18kaXrJ+V32VkpVk0ZA6DmCWOC5UXdq0/rBSFH5m5RXTM3t2g+SuPYonLfmAIB5I9HVaCQ
3YN7rEv3huUW/pEMB4J0WQTV27Z14kczRc2fc1U2LeU3VywaPsjPZvIkH/enutL4ohy6CUoTOQT/
qC86gWFQBKehbTWi+CskWh5+oUSoP6YgLA6bcTOLCztcenbIeNP1igiJIRioHflybmtTI+67dEYv
sWf06DsRgbSAZTKS/hiRDCT37t6Cxatz/VD1ceTbnnKaL+qJQG2F5zON7Wi72xNzMLJh8MbcTYS0
pcl8We2WMUc0O+QeEzL92AHkgp25vcOQ08N2fpDSVTUpfM2h/KYaYaumeHZsnI5v+JAsicwuWQ6I
LH+8pk3aqBx4fFdY2oWuTRFMQe0/FLsopLdaiX0+VW7WxIrdOD9cCkD7IHe9I45J1mBQBYWc9x3m
SvOKm0Ua0YsElJu3ySry1VrTXxgmDPpfY0w/9tppgBtah37TbSM6uEpKRX1b4NIQpLJJ88R16+X/
JDN4CkOybR058UIi1d6tVkKH0bldNed78ZKhN/hMTe88hYqf+2X3vFH4II3JhtF0foyTYK49YyhR
DIbYwvJ971CRsEwsdX6A/80HdgjmdQBA1F8aafRstqzS091wdGqSxAkQ6wbNM087fRjWAyDEJ6Cn
f8q7HDDPtxCZ3hTfiIfiTKYkd0AMK3FJ7gmCErpoKqRIwr5zVp2OMnQWziqYcodxqgjJ0/wKplYY
BBf74ARbAo2UVqmrXAks0ZtFL23nTSu2EC3fb+iE2OLDFYeZl+1zciOOP1EOGnpUJdAmZ0rfS7X1
GpktCMS/DcTvIchjbwGAMxpqmCAdWAg/ZpfOEOGgaSnpQniwrWsjMwpydTOVktrkDZa1YApwegZ4
VLRQBnJIs1WDte6+qM8xDAflNEaYgtEyfqRpm0IFo/z4Bbx98aLQbY+CChhes0AbOjwAUOI7anfo
/F23oEqYwEBsgUGBBXQyacM6iam0/GG8Ifhn1q6eoTKSq2oQTfNpakryxA11gplnnuK0DbMK2vdG
6H10xSXwuJM5bh5fxlD++NJmaouKG3c2taVKdemMtVxt2TEUeNM8Xo3eaaGNGwm5TRfeNhAgcV5Y
0cNl0lp75tnmmo3Iie58Ve+snAIbqIDOITq+H5JHc5JRMm6FVjS42ZckojPkZwOV8oU94RY09V+j
pNlzfnDosi5Ai1kRGEcfMVMpC4hcvUqhw5wEgosDpZNUl3u3JafC2WvczRjVwo61TjjMbOVLylZs
iiusOgqNZq6tEhqytUQ0pBZPg70kZoReAOSglNGYmAqrPsjdblw2c96g6pXbNmjE3ole6Q6XtN9W
TGLFxVGU8mPcgjUcmQI7ev2kK2zh6K1NGFfWfIJ2yKtri9U3Po4VCNx0diDVqdG4oenTmJbZlAf7
V6lrfArlKDDcvUYYjl+ZJwfM4NX3N98Vb+XLktEftEvKMkqodDakf78XVJFYD4xRSSGaerXci3dy
5r3UvL+qPRLpHEndSaNnpZJBogMg7PnmKvCnqJ/o3PA9AbfX4pBN92ly6AeYU4J/46BxD/PO1fmY
hYPXozO5RnxGwSTWiO/iHqu1w0dAcl3d7Lk5iIVpHHog8kHDlslDuakxzDtYlAaqxz9FSrzMJUaK
EYz5TvMjaPjFmeqKClH07qoEz9uauVob6ADw8UDiojuTZxGfAwgFKdm5lBRuDlFQDR4WT9AiowLl
9Ml0VXioFINyMgri3qP6IcUQN+JOTo8eIQtZ9t6e5i66UyCXFIdGtiefGb4KaOHwi6nMgwQI24oX
WZxA+jl4Jn88cXgMCjUm8uWc+3i9l84UaEiugUFFEvcgIbl73y1in4tBJMBZ0z02DlMsFcVYeGaO
IcVDFs1lZySGaavlWcgA5DaW6I+xk5aSTEjqzpUs7nUHgY34hb/s7pFOdnoCrQHVooNMF80JLCq1
/Q/UvfOLZw6B9AESwaXkCYwkiwRmb6juLvt7KZ1UmdFAgdAhZORYgQbtL0TqXa9grBhEbovklr6N
IXM5pAqic4BrMR0wvvz2EB/lIy7m9UFn7yoUEQUhJGL/lcss4K3wEu2gpEYVBMNDfJ62f+kau9Wv
vOkFofJNpW65mCVftSnjY4xu3cUWBdOQvUkYgIUHapBJqn12gOg6cZq7OWfoO1Py0PmYrWLe2OTP
cVpibbtAhkNOd9y9PQPncaheaY6KtmX2RHX7FNCbgUdTmCkGXGtVStbRxW2Y0tjB6K4fG5+NVI7D
+vLel75fmlEAJ/gRMeVSwiKOX4pZ/+kC347WdM2P5uQAbDh3bv6iK5Whn+rA85LoLJQ4BLNr9YEY
5iZNFKACiFwbmdheancChpiK32e9SP+sk9mnQRUy7EsjQ9pAl/AFLN+od6F9dm2N8GVm+vhOOxK0
M+w3MZ4hzKFIKh0GxZs9WlPpvtE8NWDCl/ymn+QVi/zLmU8pwPGDdAqt4itnxELyOlX6oaxdg03+
g1ZVNSezmyp7t41eD2eX0ZgnzJ2VVv6yb73aSz0zEg9okPOuOASvoEYMVLV8X/BKxI6NzTriKfZv
//IVLfM4iNbBAC9isRUNf7a60ft/NHmR72ovqTFRjErlpOe2U4OTOrgDIPUc4j36E+FF1AEO0crB
qycPFp0y3Nujz2c+/Qo0O1xRNPNM5QyYaDDuyij/ZOFPbKYo/7uJFOBSqXObX5JyiEiIF8hwRn2Q
cytS+/lB5hWYLDgsaiW/vHkIeUqZxCQniaw23A7rw3vFKHdt8DY+/3HS29uwH99z0oB0wACKVKwe
NAsEYeOeR7QZHDbN3kB3ti2KNRiS+oZ56sdTO/2b+bW/twfZs9tZjykEpO8TTJC5oKKOhOf29nx+
WE0nHHEOoCgfzytal2104ZeL9AAXf59ExibEU82LKZBUATRkfLs5iNvCYigUVyK9RsqsX2X8nn7+
CCJ8sPnz87ZjCXIgmWII0wEgA5YQfBhfp7uo3jfCEcsoOhIIjzG3EXcv0uedzhyppHtBGQ3ZNNiK
5yYIDYxQ06iRVy0Zh4vEXIZ0aBs6EgkBXFaz3KBl5P5Gfq2vblnC6yQs6JqMGlwZ62+OoI2jj84z
cyHZWxE5tjUOlmishHq/kzbTqGZsobrhGD9P4tw5EBmlY/VPCdh0Hkbi82ZKv17u6dCEZuMSnGmQ
PGml2gCbrTf8JSLnze5ZF4CO0VrnDctbBGraTdgrBXZHtvmKoBIvK/Wn4FGGLrYp0qw+AL8bUsoI
RxjJbapJN7jKur5vFGr9e4ZZzlUIdPn6b/j3iMxE6r5qe+QHLCeVa4RgdffoLJNg5cnro6tnhLwx
K4//x2MI2am4/BNDpI2sGqooDG9l+8w8sha7JnGhVXVgfjjS/vM6fZTHPBq4E0LpeVyqib2QjD/p
AabqVeoqrFGkvCkTuBWqSv9WNyXG/I3uMYfPzbictvL+a+VgY285dtStV3dg/OixDWzmJUqcm7QK
bWe3UOKb4FmMWFNKKdOCGg1zpGkaLYkFO6JjFLB2yHQIVXaNMvhY11y88vfPS5e0A6cWt7BjyQQ3
17sWfhH7mDt3ZNAoqVeBkBfk059B7wSQ+Y9BDZTYkGgpSA3wPj2ZBXAZ83jIgmfVpK+UYSjMPNBq
tFlBwYxRhmY6MDe4BYIZDE+rCaIiXi8bZqBwE661mfadKLKiemhTAIGIWpWNsOLbITFvtqbxsgQO
wTx6JNax+Vm2wHhEvTiavridypFnUGqRFLCaxlzyDkn6v4AjxEap1VPrhNtgYwD8L+6CY3PwpPNA
7mRBpEMDFbGmBQQLTrjB3OL/wA/zw0JLF9iDch2SDnqBHInbTtaEinjbItaoECqUCtuP0iQ/nVo5
vKmeWYupukt9/hLBAKkdicNqJhf6Azx+jzqneKqpiKtUurldRg0LBPnPuVr/YD/yvyZi2bkf/h6N
KLDbeReqSHDK/x/VQqIxiEOdwRK+6+elMP7PLDyUpIszJ5ZSADM+6kti5WvxR0bQN6ZIge5ZWdhJ
mT/L9Up0W4reKcKG2ziLeIoDXLaVQ4NQ7Qg4X/rdQjqRKJZgUL9LlAG0eMm3pgJgSF5JSEYH0XyM
CoxlNlmMO7GhL30zHtbKt0VziM8oYQoiYz1j3v32doPTU/z0dQPst9GRQ25hsfwhDXf1klTUDTXv
OFvemLvGm04QEkS+63EkA5lBNZebQB2i9jpfmflqkjvU0jEd681C1K5ZERIktOBrYwD0XFR+29Xk
vzPb7qjlxmd3ZwciX5acvOmaYqAansfHTnorl2tSBXAgWceUu00fH2Csiii5RYIHRRRHg5F1Gl4t
6X9Q7gh9GvbzXkNQR0e3yJmHGu+VIgfgWKVOx/WWdquMyUPfT+jR3JyemCrIBP96mOIadCHqNaBU
Vg2cnntwgntqykklb1LSCLGdvTRLxmECMcxf+OTUFMyXtaLENN+IXGyG0l1pNCGFfFpSnzjT+Bwm
WOKVKvuYgfV0xWH5YO6a2ppe9HIxljJnCYU4FmJvGE7H1RYT09BgGP/JbO678gg8LT/cOvIcJeqf
55wHUx9DOc1PjHKaUnQfEUjpakPVNOYdI5q3dcWp7tFijzowbh7c+OwIxPhBvzXGfgSGIARvYwkU
N6/AdolDyzJwrY0EigMaErrabLEnSXqilmWmXoBiN6tMPUKA6cWvgoYyY3mQTm4urhM2uA7Ls+A2
IwH/8nYYpwJ2gdhJFeU7GculPdMEayvTZ3Wg6ezYyIG9V1eKjm6wme0bdfgw4dFja4lDfp+o2Cbx
p39sjWHDxzZoOKi8CD4pW+IcNEMqqVi4fdn7cuAT3MvsIGFmMtR+F2VVRCcBDMkTCPKrHumMR9hE
RO+0M2MrewEuhdyVfCCZBRuENsiN7c61VjqjcuOChxaSz9Mi2WuJe8ZJFkxyuJKhZersv3+HvTXh
RbWcssJLfj2vRgTx1aXWbwVRPR0UykzsYICV0HZ4vZe7amy4ElCb4RZrX0BGZEb/546y3K7Yg2v8
z7VKnuMdyFr3uk60m3tykp0ReBB8VZzFeHZo9uE3THAHNVIrUCiofJzjZFk2wgascLy9Yz9z7aRh
Z87vJ+OB+LmPe3LHimmOjmg+hjiUvVFRsHRrnQJZKn6bYsIcaqHvXam8pWl+J14OE772vp+Ll+Gu
61qr5TAz0H9CUuil1mLuW6wJd55EiRpUvR8DYo5RfuzbkSee0TGGZrledh5M+dFJwiO9I3yeBcSm
BEyinrA81rjh6fJc7qWwtvYYfjuPkaPI9kOweNFB7VY206rJbwA+cg2AohSCCrfD5iCtK9ZzUy6/
ZWub15imj2d64oe49e4CV1G9dd8gFgfvqNlkejvSFeKUkG39YEU7s6d7yzSaN6iyHf9yPSu3pnnQ
n1eVHxt4OK4Dd6ZabFF8LBNI60+Bmoug5hRY8WcrMfiAym8TgHnXa+GSFhzQv2X3CFYjXodiaal5
oFqNk9FUwETdku7Fg/7jW9zZoZN5XZBz4tGH5jtSOZ5pg7ymAjQHP7gAu2FfJEg+HS3OQ4SAMqPO
ZKLSFedaZhYqkkSPqOqFobwJCeEVZ/cGvjeW5X4ycr7G9HC0DvJZM/5GaUPBGB8hqDHszxZUfGWl
MqNRaal0SOReUEGYNrSo6oh70QMaQQcjBDWX1c7JzSfunokqjLYJDa1HP1vFeUhtqfa8g99KX+F3
UiBXg/zT1Yk67RCN8RLdLeU4dovzz0G59tnmxxZqUfxqPgAmqhioSQFAV2xWsQQx2rqS6Ah0YCiY
NOrnfd4cPbxMdzH9xMTcV65Y2vfb3dT/cNIbnkITTGXqLbfBCuKw2/KPLRetS0rDcTX1sBa+TIki
0YDPYWb43f4muvk83hUrYoaNmcMIw0paDRSoURnQ/9WLl2ymdmhUrXyT2Y0OEYd/Vvsc3iYbOX+2
7uiq1nqVvoYHY1XG+1sDO9lUHX0O0f8PIIcKWmEk5blSwDPI9DDJ5bhKeheJ/1dam8ThM8RwoHio
5yC2D0PWUNDJ3eKSdbUz50cBFAQ+/J+KdbN/Pc99TKInloab3D+ieGFI6BF/f718xxKelEiVLYJ5
vyiELFO60Tgj+wr9jfILZz+0WKa1SUzP/xIHJ7RAR+T53MEqJFMKz2NcjUjCUCbdv3THoHBMZ7Ro
vjQeaoDsVRts3rv5gk+JWDtomUKH8ljFsQpHfEx1LA7xUMn02dUY+WfUisupBPK54aDbqE6fQRBv
Lg/4AuP9VO9lhy3NeqPOC154mrLTOg69y/9v1wDQPQeABkBQTUxwTLWREeKR2ai6E0bI1O+KKSpY
ZBybb8exE/KzoKI8jBm8cKNkfLoIZXg1XSLSD6IP7FJr1Pha6VOnOGxIPDJitjwq8LUEUvkGp15s
QsJO+MVZ4nRpQw4FqMVmOgAftuKd7cyviH9SQ744Y3cTKAwHsU/lE6I2+WsVWoHheGn8zA8ltfS6
wYQKGl1pawuNfEZsInwro7qfTQbr+cqVEaqn+ykKJVHZjjzdefjg1A1MTJX+8rdVgLa1m+DLw++T
lARSbhkidA5Xb7VpYhEW5nwmV7IAT41vGpVh84BegpUTiSsypiusggkOJ0iAGye8oYrAhwHihwCm
2396/0fKHgWIfHNMY7PMzJkmqlmzLOqP0iq+F1IGxRyVFZ4H3cDmIUhDuATlas2CW005CmHhvvtJ
qaqrFGrEr66TQ1RIbQq84J9bKZt6ubjOcpZeey3VRR3Fg3zod7+MuoHoumq/IF61dwPvOHXo0Jyt
7XZlsksGeyOoXUpVSa5lfxcKpOJnnISES9mi5E+DwslyQvqIOdg2Dvows4R6AbLzBc4Q+wOFRG56
XOQVQqY2LrSAXdJAcdJe6LFvxNKaEqPdWYAxyAnU50HQST1SZVpdWnUjThDnKyXjFDJnLua0SoIc
fIuKU1jqETQiTWLTRdiNOpxHrFAHHNFyz0F58ehpgg9YPuBsClN0sv1+lQ2hdg7nWNL+b2L2BPAE
LVhi76MpliZvAtuGoCkQmj64wWPRRtW0bWQsR2afS/YYvU6X2FHHY8qW2kSsQ9Mh5tYJ6aylNBpi
GZKRJdt1e/puN4/gAGr2sPfY+GxgTeyyyGEs+LToVXVnSLD6irXb/5Tt/xauQcb93OAvAbZJcG6B
CXIUxK+p0l6acGlDlcv5I3UGw45AQT9++J+mzv/k9JqTlIAhoNZFnFr+0HJZxRMcyavN1GaDZdsd
HYdLymi/8duvTuJAVE2f7XdWDoB4HFTEBRwXBN4IfS/bf+G+neypDG4WB9WOlOORhsLrfk4JVXSz
3J0WFUv2gl7DnPfb6QxV+zu18RnLVmCIo/Y+0x7JMLAXRtSgnZen6slkZRMRX33c+/qMf/FJF1M0
tYF5Xsvc2XRYst29eiOi+94NRV05QD7fFEWTqfN8BfsLgr4cj7+f4yaUWaWSR/IIyaoNhpxbI+w4
fNR0KvdhwPOoVaQ5x6qcxbyNEzN+8hIDiskxpPRQqCa1RiNOoTKYuUoXjKjS60MG4Tgx7zi0ErJ2
wP3InnRVx9u8u/plA7sgHx2GNQK4o3f5vOeHTsSGoAQnslEyTZDByPluei+8V59z75l6ukfio79A
qMV6cnmt2nAYmIquQbOjXATgQkycIcg3zxivdX2GJFZnni6pKTnXNrtCTVEN5BxEPtnsI4ni8ztS
NSnLltHpbbrZbdhkjVKUDp8zSMvOsWmDD6XvCZJ3XEXVb2sst3Nv3iBHpInTNie3uMIQwVBDPRcB
iBNnel7pKW4l0z4sM/S85zOJeKvnzF9sJgGYcN1eqOUwYyFjeN8LRdXVVZqpfjyoyv9iY5If8jkp
vtj9fRVOy9Qp6IMFmRA6DjWuDCDgfb2upNxu9pgqHj56E3xyqhVA/k/OhJG95pb9rjr4NYE2xsl4
ttIfjuSMF2bUSIx7732eWLkTTFCIRfcMnNyVNqLxhAraY+S0N4yRQLGzH+h3S4q35C92ULVzdTAc
Vf1OirVvQXui0l1sypqqHN/MGBboOPKPBbwk2UFt1uxhD3E9Jg4Y4xR3aOHpIm8wzW0puNbG0VmR
z7Cq6QuX+41Y4r56SrcT4goKsclsaWta/JpDZ3oKVz8Pol55aI8pWFODy7x+et+QaAC0I5B/EQcf
EJ1N2sw/Xy+SboANPWPxLTQQly+kn6kzM95jl3aZxxmSyOLZPk4NJ7iZrYKPSIgCvnwU5bD/kCZt
ns3svSVxH7gOzWeRUVke8cbw7e1Gl1pr9wy0r2ZR7zHrxh7GBs1a196A84KNDhir4vLZYlj2vkWJ
evNwedasv39IStF7XnibEjgeqyzINo4aKRhzRjLdhHdhcWNuXb6WUpUlOhmPT89bks0zDUPHmG8o
FitpC2vb5kygTEK+ijlAe7Mvw4cPXK7UhtAqKuc0aFYO3illoeb35ndvaqrRgt8Pgti1w+PtHzeh
JtzS0XUog0yOrygnXnBRvRGWjolDhGW05KbPs0tpef1iVYtahWTCtRU4ImUAbveaL7W/mBRJKljx
q4cCEKFmdH03C6o4/BV/eMhH2Kw2h0mnbYa0S2Ub5Ktw70qBCVUzhR1gk5OQVANpW6OZkMs+Tjd1
59bCHAto+M36T/S2u4I5vY4rWiSIlX4qGE1rQbNkyrJhHEe4aatUS6HruKMqZ6SyBfZsmFrIDxgf
+z7pLltnEPmUyxXu8v/eIhKNl0s8la20pBmg1HdSxYkYlKxx56h0TeFO7plT4XFXaS40/O+jI3Rh
xv98lpLVreZ1N8jL2fMsNkoTKA/jLtZXimlJj0s96EEYvmhAsmFySKHSNmMBhCSI0VwIfzoLc1vO
cX8QFVQts7u+79xZXO7QDoNN1puv7/naIkUWESmtGvQ90aavTZghrYDLGn+WXpqBIzfj8Hy8NgRe
v+Q+hfX8e4d9aSwyMQ5sUYKpjRg9wI1T9BmL9fflugr64PPGKc9DQsn3d6wp6Az9aQW1/oKzA8vC
HMVkgbQngzxKh8zyrqWRWO/tKuIoi/iPq/Kxj/rqb6cB2G2a6bdA91XHAJNp9SIcPNH7NLEICmmi
IIP/Id1zPc6SV0rTctbFF1h5h5D+GVMz8k6SRTdiLWv+RHVBc6KNC/m/fsp97i9OXENaokZq7IxR
sCxFl3QSsbDSXDTdDaradDRqPvF5MV0P1OrzBPVm/mELocjpUT3nK1IJNkBsvoyTbr5NJRwxSwZo
bTQMzTs8psXlGwoEZckhebleskRjVSWTDy3JqJs5v+jJIfh9fjZ98zZebYaaFzt7gds1e2EXckG3
6LRP0wqE4CNNAzrIR+Xv4AhRISIhNHsPPWdQBKKHwsOXnu0BxfbNFH5R4/pjjqyiefEyjc/uKSSL
rtvoJadrEa4m7aNQHRDEK9E9i6Dgw60XqgewNj4nupHuox4uV/2NfVCjK7Edwug7SOTtOUZZtSHK
WK61rRgTkQLcjAVHxXeVmudqE5XY83jNO99xMo8CsOkDRIMMRnRoGJCnryPKmKpxO6KKWlQLFmjP
32xJy6aw/zbSOV03gQZw0t7n+AAUgLjn7pC44Jr3S/6c0SV1g15Y0Yd1m6+0eLZB7tsa2tf7q65q
O6E2pWta2TDWudQfqHH9+XXpNZrS7qolOvHPw2z9+v5LH53x7ayrBhcQDxo+4xcxt2iKpWvNrNOk
tOg0T91EDIjkgWl7Kp/I02Haj3XwaTlvj9awRgm0xrECCBXkLxzFtBsH2RUnx4Mr9Gp0CQIg8Kh/
Xe9k1btUwj3zzT5hnHQIzWT3HUqQylP5wyzdwdrVqQRlRmp/BYpWiSLQc9/dcRIWm7KL1+c2nvpe
PH3ra5nqgDEWiEKfXM1cdd4CLrn4RjNEa+orl8nHuYxB04jeYTjfYXPwhtRpSGDQTNj78cV6VSoQ
LPGcyPkZe6EgAQjMBK/4891VYp9800Jmg+7qfUXd2dCMdB/NVIpCIdRv+7noAHkJWLajqjPgD+7J
hSEK1omU26LVjKQnf4xHNX4+iXiqH6ir8qlhPYKxYajyIlSKorbClQE9BuWvq2HyqIL7SA+RQy4U
+2gduHaWZmGZFHv5F6TlBLRtJc5ige2zxhEZvWd59Qmq8g2OPTcu/Rn9wVZCULQE5bCW7tIpmk6I
a8I9cx4Vm7ixWsCjTg6TeweVD3QvDkaNAVCX+wL0Fp8esDFwIcm1OqeNEdRI7iNdCuVr9yjcbmWK
G6cQOuv1lDkcOaRcLe1jtI8wra3uJ/SbIDjzQV0Kxx64N6cryv37a/pwWW8+IDaAgPV/w/BrfkAy
pOMHZbErpmc6bbSvv/LzUeILtA6/60lj4aPFWmK+0JCAD+yhzFdwjTlBohn1Z8vFv1FKDsilVxjd
s/13uaHESku5bJSlfqoGBUMsOn+OCaZ3/QIeQRj21qLvLejJEaRcgSsR4pcOU819FxzaGZUVUmaT
EAjn4+jiAYXVeS898hXy6aWDwPCWqLT4Bjl2tcHXLtOkuSSA0Th2Nmyxir96yhRqBc5z4bZ1M5c/
fkEDOKhkAlvf7uyxR4HU1k7LrtUUSM1bsP622RP2aVAZ/UcN1vybS9x1nC2Kx8vG99XDNb3BRq80
fqTng/132hSQITBIyq/G9qG7KTGt1n3M2TU80IrZQTCaPz5NKJLAi6pED3YA1zGMg7fzn2lSc7yq
exL0jQhdwkPUdr/PPfqtiVqofNOgoOmoPgxAwfdSzumKPp7zthPuuyTnShMIcwKs/Q2VUc83oVCD
bCHF+fQDOBbmlLusn79rplk5i1rZWAVcyv5o45AL1KDsnpM9xHhPsgzR4CDW+jipvjLKqO66Rtc+
tbBW4hfG55KZgTWv2311Nx+RhlLRm0VvHcGUapcaFDxC3M+/gBGqRmJA4cQjzpQOqH/L5DrTeAxI
0TFPLBlJeavdQc+JBKYmCJIXFX+mcTNp3bMAvneJJcDcZF1GvUpzPRXa2RuioKqm/9Kopkk7kim9
YgCkFggJ0xbxyAHRtgyIUzfjHcbrCT9reKl5VLmzIV6kTtLAmS5zr8ixLciKQWrzP4JH9D+u42RV
y2qXQPVha8Ejatw+lEGrUlp/H1NOMc/2kRomXsvTwhjCQ7DBxckie5xVU/ElSHhUno1wa+PERdrg
yYdQgKx+Pblnq7E1DiRyx6Bh4YC7CrU4OnwOTlJQcu2YrtMfWHjEWyq7FRz3ms45f1+xg/q8RQBE
yMw97PhABCzgmIpJs5uEDduiEavwQ+CtfE1tlWk6fKbJfqC7OlKLPj31kA3NM+tWL+8VNdUX5Y/I
Lvh/s/JZhp+CkkP31IeugTDAamBGU3dmofv99dKOgBfk+SmPMamEPSSxil7/fMH7cCn27fmAuviA
a0Pzp3tx7RwW7bCc+U6pteXNPZvd+Ce6gSImSxwJ9yRKOXjkPVSNna9+M5Md7GftfqZIjCrugryW
Pjjsoxb8CtKB54zWgxDjSL4HJWcaHAgSHL8wTwA8FJI/WUa5fb5+myF/DO9TW5U+AXg/EvCeHqqv
JtqFoniiwLeD2fJqUAO6BvsXZcu8vNBP5gFBGSQTTVLTyJMNV++A3btwSdj0ZLF27gTUfGU9v5zg
RonLiM+QMiNsb705Woko5wBDjPxwzID9yjdbWAdtFPVcxbvjSSvpT8Ciq7F0cAqwomut5JEK0Z5J
Kmy5ZoNlT8A+flsBq5pWkFrnXpPha56OOFoNWY1m5Dke1DrGtlQaPBTiRlaVqd6BqGAMd15VSCc8
Km86/BbzIOWhIlCtkk/rZaFIEl92pCU81/5654QAnS+vVw5g5YHZmDnbK77ucCFiFJ3+a7Y6HuOZ
f0jwxj+Vd2e4flm9hPUiEj6wZMWJXptBi+pWc2d+OKbHnWJm+0/D17eImlxEUeDoOWgxNOOGqOEn
wtISRfi2hBkPRe3CeM5MPnH3xKUfVRWFOh97+P2CxgF+qmVgiPTshvDRFpauajGkCPoTojm7Yp/H
zaY/74iMXc4A63iXv584OkdZ8BO3hAQA4IvTEgNnLjNVBWor1dBuWNs3mAFgtcEAOWa6L4jp3Dg/
8+Zjz8M+MF4N4483r4WGjFhNzxmDqOMIir8a/CE0VIkpinnSGYwmjYTS97BsVp64aYIwu1W3ohTO
9YvFfVfOv8eYPJJsAV+S3w1UVvVhSfz4u51ARNAF5Toe31mohdPKkmYp4oaufn1T0GfwwN0y3hkg
pvcApdi9TpWr5NQ27jUcVMzvp4hivlQ7j0oxRUMXqPO8qbMIAydu/WCisedFt8RT1Mb/rhEgBbii
EWpNnEx4v/TN820g5u7p+8Na+3uB4lG88gb0iKHu1iM4oip5BhyFSWBVVQGDKsqlFPOZ9lPukpqV
njsnHKfqVsW4XbZA8pXF3tukCa6F36V7eE+WQEuxvQSLJIgTq3REnhNNtLIycSZ7mnodjMdYK2cC
sATjLqAz/JvBKVQWJl3HEoer8+35Z2JuNG4ws7h4qhWwqyg8kcGu/NAPsjxKIYs1XaUDSORBpPpd
F4naOhhtcPUhhHy62xbvhURLFo4UWj54nZBMKjRqLwClg8eD/UbL3TKql3Y7DW+djZfakFEp5of0
hgTGpTKAglDWMl99KNPDFzRWjrQyKLADCLayUzvMqe+/rYi5Rfc24mmQfZvI+K4YZ63eI+OCpfLW
WAqMt2XRUSEfnR3jAI3ylr6yShWWKw4jsB940d47kar/MbLmobnvF7YjKMEUWVqNh1/ddqNeYATI
eUhCs1Nvn24TOU1O85xP+V+Iofww3jp3Oal7tLLV7XMHv/Ma0em0Twra0tlLwEC0rwgvBsvOgt6z
JF4jPzNG0JufSnTwuxb4kZpRaC1+f7RFxApJ/86lMn2TaiaBZt3HBqYMTvBOe5bwX0eNqKgGRILx
e+P+52E8Kv9y/kR106mn2XEkihXgm6eLWe8f3saMxwzMSuc5/vjOMPaN/2AYV3PNqqBzyIFMJCA8
06vTaXfcTU70CbB55CIU+rb5Cvj+SeanBcHMf01mlRboMr19ui37PPthqPfQV2AXgiNvIN0nr7ii
1FKQLE8772it5Htjgu822uNxKXCW+9K+vuOGq2GerUfUl2lOWi/o/dO8duNTbSlCSNexp/+d4qcw
zSr6AJnlAfs5FA0umCNCuAAL/SfGq9T3wgHRl2B+o5O726vzxKOQ4+APi2/toWVmFAPhGnzGyJZ0
zdi840MPFUyGRDDmXwIsIOYt31jX1zuvrUF1uJDS4zHubwpxW7yk7adBP+EY1v/n4NkvFlhxKO8f
rZHpuEbkpv6gKGF1HznPF2cCSaK5zY52EldY+Y151eRjj2IscUwKH4Gm/PlFGI3W0fb+AS7sZBJZ
O2vxRsqKCaRg1ievXFUUM0r/OtNH6MVE4WcKW5S8EdKocaGtn91g6k+U82jO0RrZ7tjGx9NzqTJL
3LmpArc8qWLYz7lQ1D49V3PzV6BigjgweDuTCN4wCS6K/ZgxqcvW/GaHxIOSmt6ZwN460WE9zRfU
WVfwI+temBetNIKMC+McJjSLUFecwkPxiAuhW4hUNC5bKKaf3lmtY2zGj+TePEYJVQ9onRocJHWU
Xfxo55gjbJ1zAcPFhw1IVn9eUo9dfCCOi9iPeVcE9/kmgBg/+TNIt4fZ9ZpXdF0Hs4BNrCHHjV8P
ZoACqnV8kzhFgwRZaeFHPjwYeTcTZCDBwy0Rk7GQluPq2JtkDvn+ARGI295ZEVB2b/3Lg3gRKVcx
t6Tmsz8OE1dpTO6g7XlJCK94D182sZ/EU1NKeIJR1xfDvH9S/Is5G3qpaYM2xwqPEAMIFmM59aFN
DumdTA5jYTkmdGTW+XRILwsUfruB66ofSBqN2qmb6DCKC8mdZAhnmvOm0Q82SO/lg2WxdKRwud5N
81VZ917CSCRdp/6kFt+gTZdfEl1NBp0RrBA70oVSY3xochgrF5AzxrvzQmOiEd5UJuyqvPqpXugW
33vsanmg69/h4Pc5V6N4brjKx0vEs4r/aScxpshVunD4xIK0usA1vpwileY/5DQWJTvXyDPJOCRA
3AbJisfs5GO0qO5qHdEKyZ34cAQ1BTw3VWe36sk5YTY7tzoj8kiDNOkH4SxQmE2/PTJujvMuiW/h
uVYzTNlKsZNZ3gGkvT3dUne95ER7FDdT0jwY/s98dwgHXiWmOSBoyX0tTCs3lkYOW2mdoIkvcNPb
JhZzmbNzj0xemZK4gtttVZQmFOUt1fGhysI5TyBFewi49ydpzKM6Q5ceSp76LmbmZPtdCjqS0Fg/
3p80eEoLIGBvsYw+yn+4hzav/L7Y7Pd0vtN9pAtQcsr2mB8Yw64V2XMkFlAIDV1WiwjCZZ8Iws5g
lUm3DEv0o8uiQAaQolU9NtkMfnB/3mdCsVFUpESthm/puVNy5N2ikUBWIUasIiGpaGLFHYg5DtWi
UO9bwckZK8qPeU+QDduQsuWD0gobmkbXkafB3wYG20P3lUhj7Zrdy1FXt/sj+TPWn8TemqiRrr15
+6KxgnZ490wNqQcrHsejOB8ZClGXGGwkQPJm+j2aNj+YnYZZ7/2O2d6Im0svzYtvVJelpqjqm7G3
/cvd47udF1raVcuydbT9NmhqG/dh/R19m5QinJmtAflz1I5ut7bReCNWn3CamC7zAAyaQM6uxI/i
5XlaHuHBbdTypTAVkzUje42gC8ehz7Flo1wDgoisp5X0wIDsqOKAz9W7C0XNhdkrmw1YOuQt6ljH
JlBf1hQWrEe4zUZ+nksPKIGWSGApHPih6/ETEKGU9lK6Jna05S3IUx5FvUzrzmobSfY1EL/8DPRD
Hh0qCRqZVCa7q1hr7+CTJA+YdPBSAONbUdQqqZJFU3yUtr+depiH/jTiOJ1WsG4HIL41asI7KX3L
YGz19TGMDms/lh2eWh+mP80om+s+RR6AxaBAFYMCz2uRsv6oYIcCj9//EOCSIJNn1tnSn7MWHWVi
iyUTYurKLYjVr3wRr3xA0AfvMMypWSsjtIBe8ljb+jgoSr4PJCxmcL6YFgvigXkQ2IxZPhv4C8/G
bsSez7TXX3p7Jbvac8Z9RgMXEqNnPluZG75HnzKOz4MD5lWEcEzjVoVr4w94YNB+LWhrDontbMpf
XJIXcCTVr7XO8AmZ0ZWzXCVX0jw5gA0dGAx3xOBCLl5W/2FA/d/1FK6fwSrljWCG6vuG9fjgnD2Z
ZQ7m7FooRAVSTWsXAHd454nuN7QuwXAXfkqBOzbI8FLOz2yjmpfnOOQwD0gusULu5m2ivnl3OPgZ
BzaiWbvRhvMYGaihqKZN2Snm3XNkSNau+T2rlBfB0aRxYpjGYbocBUA6ZnLUArUY/GHdW3/uKdft
oTiHnbx23iqb00+mkAgOkb2TMO5A22TJhAw8iAwGL8+jNeZvRUAAf8GD9RwMFMTpnVGdga48S31R
/bK6USH0EcPF4AqcFcVwFraqeDBpsqis/xTrqTZJWy7LKRiqD0yhDpmY4qjXIM58jz8q16Eqq6Sg
2EFfdzRlW/9Q6y8ZPhUm6CzQb6rvkUE5uSJN4mgrt1Ir/grx8HFdTiBlMErFI7MjD0sXqVM5OJaF
+hMlgehK+kJWEFTQTD3FZRzHWQxijrtq/IkW0bT1SD2JUOu8/p+NOg8ZY+paEbVX1A9d7bkMzAYf
C84Js4/ffwgRm5lGQVjDHaw73/7k9sFrCh8LiWoXmY2ukoG29KDE2bJvjiqWeKVzA8ygvbGwC/YC
JDP3I7JHDPJIMunXoQc16FJIum21ns4koYN9KI94JS0U3sH/zkEC73tjNTia8qmY+fOeOOQP3p1/
cVtln0UjHmtm4K8L4Cgj9dMXfCwFTk5eZlTbdqkjNID3zeLQ7OFgFmCzZUExVrzF7zYfVCPsFDgY
cbpA94c62vLb81pDKYwfZcbVasTOW4qgJ4EzQTah9bz9w473FOOBTV/qbvZsY+o7HgbkxpgJsVhs
t3TodDGUYcpiEdhVBKiSm39rqYk7yV75xDKVbjYnGtVCLyeD/gcFK+9X3olOTN3zILJshnszk6OK
cEcdu73pEtreQiZ6h2REAS50hpPDhS3GvL2JOn9AvNB6CMp1jzlP7FBRDhMFdgJzVQY1mU3NJjeh
YDE744AjkGLoU8TArOKHNeYVWDXOYPLrMynK+c7XIysoM3SOum03RGbtlxYOsWIxguR/uGr/NfuJ
Mt1xM3WsMNAp4JjFBXAzAVQvFLpijcrMkwn9CaxZWeRZGVzP3SpiTkbR4Zt34znhNJz+w31LriO+
+UylM9tPJtHDkYJmVwc3ifLapz2d0Rc0SsdvfFAr78fLi521CizO1lyxP3F7oj1JhYuEBtUxz7a3
5gQIOfQgQDqx985JX4R9/xuiOJolggHICkg/1rkV4aoMAO0hpKX+b7XEoT0z1BlBCekRcKrqk2p/
d+4AuwVwkSzsCKQrf+WZCn1rRt8YfiCqpkKlo0tdjCCmblUM3pSUEfnYB1x+08xyGP9XUahqK9Mc
8oMh9zn0xLm47Sv5PJt9nSLucRlEYmMripBAA1IYKo13eK2OXO5KQk4kfD48oXLiExdvUrEF6/AB
6A4brLvs1AuFe8xrsHW8as0iLtyb3wjRbXy95L3TR92WQGa4LWVdWabJ6gDMTl5m7+2RUhIJFsFR
mTCSEHuyk2biicjkncxE8vppPoXvg+2DFHjvYbGxiPAbvFtyijL/BfbyY44/SCSnUZQIPd+xK03R
wC4D1K1OPENccvoeZHdPcQ1s0tZK0TUGKJg7RAXaoS/vf2uBOgd4mzPWi1dRi4srG5lIbFhauzJw
2jYa6p8s07dqT8Qebj8VDmahTLU3hfeth+Nh3GbkhlRyW5HP9+vux6eUdatpBo77BW8SusgXfdZ7
zlkClFLfZllXUGGmXPx58akTqyhzYpqqLkmCjP+4zoRiU/f52oCtv4PdWtpqD4v4wQX9sJ6jzTPN
+JpEqvt4YC6uR/lpSbRTS921FF5ppzmp3XWN4c4HLVo0CbzmATl+bgnzzxHCXyuWmg4BFoi0mzFE
Yi5Csd/U9HqBlPtwfLIPwCFOqF+0h6Q6q3U+NwKJzR58eMLTnDTzrSg4Th1jFneHqBOhCQGnl47X
pUx3nLrrlt52Vho359sVZsvLPzb4k/XjPRf6ChdXthROC1kPC5eH8w5x5t0tTzrNRj9CcinvV1gG
LG/6iuQjLn1cGs0PaskRXOsV/Ti7PGopyg1KvwFPomEbuSP5I2K6TThjtUDfH9ctw0oPZRE6Zd8i
iEbAOtBzMytbb5gl54qPqUvdpoZy1x04lnxVgRlEqB3UyXADTA9oM8gWGn7igRzNhRec1kIQTSZp
gJblIX30+Bx/8y1SecG/idZVnZ6+Xo2KJIvBxnkkFHW4O2oz28p2qEjL6qo068YCRRmTcPHZ1Rp6
rf0WPOz27KpRoPmP48Ta4xVU5FYeCJxanjNOd/mxKYsxmmXAbmGpSrXoBZwgIL11dSK3rcy8DsCd
+uOjL68VzQB3NOVhYigh6a1DMcM4G576N9y2D+4dJLKvh5EQz309dH0qP/WWEI+33zCT+yglYcyg
hd4rX9PA60P0CMNIFgDjuB3XNCrWBrRTfe1+nK0yCJ0Ma+R612MOmGKYsdHB5sBSSIdLUK3kl+Uo
ig9yN5fbIOoJX2b30unAUQICNMiNAzCl7zr8TPnwGSfOrLWmn5/ZaQaIhVWKLSW7Gct7Vq8ZY6zD
KDcOsnwLxCZ7g1QSRvBrfRRmJSM2D4+KkYNML3HDNnOIkguF5L34bN1w8xnlxu1GgjIpJjMnxLfM
1Fn/myrWp7JIcqxbHWhZXy2xs1lWUjPpVQHLB6i7duK3oVD1EJFoGKlcwEGmGwTBIPqYIQXI60iI
Y462NvXnBwAmgNIy7O2e5CfQuPd3sDbi8aYdFPXCL/JNjldEfxLy0m3iOA+Gj0w+ahUxIr5kECQy
oX9n/kzD0ERrCSp05ed/VtYqSKXx5nzfkaUc9fo7Qvo72V50mKJJdvQdCOBfEnHa1gpz34Bk6IhG
ykmjEZC7yQgtAXYp/mCBsl8kNauwpNvmQ7IwtGa0GsuEYFt9qA4ew2XXabZ2r0ECuL3zjuqlD/8l
5sDMntP7Q4bipeBKirNz5YVZxzVTX9IeAh6l9MnI8yzHjfeO+mfzzN0yeLh8g+NfR8ezPNmkuiGz
k5Sl2zjm7VfjNka1rSDeS1HAHBupbCNOCSgW14UJXgkIbTILnbpq8cBkV8w6jVt3RAg29Za63ZwS
4c6dWnxbDI1cDHc3aSkr70slG5OPPaIpoEP8SLDIWou6ka74nQE8Az6ZiY/RcrzCHUjwaCyj2PaC
ROFU0CqLrIgOpenBcryllR3FhVo02g7nTlWEdZ44yLSgW77yqCmfAQ2uc1ANmUV3NWYR0I7dqQYg
PVnqUymVVAiIbmd1MfDalI/AmimY/darxet1kTFgNXoeJqcwSxCJWwB5PI22BniU65C414/fHkBR
8hNbMEjtheQEitYvt2fFM+vtGRLcYSsosnyo2fpLTSsqFUrBj1IeW11yilEHav5g+RInRDvLXQow
1jqHSukXVWgYYoKtL0LAlRSyu/LY9rfj4bzgjpKapyW9tgEDKQnvdmLsU4DvXc+GxwRC7pfz+4J/
z7B+x2laZgz/Y2AhLyyq3lp/OEyDx53WNoB2vdbtY9cv6LNGxqzbL7E6ZUR4siFJh3UFH1Mn3vRA
nrpPFviZ2Y+BEuOOeUjBokHCozBLgHMgepablpRDsMUCuSaZIEC9rB4+FxvJXWRoA0Q9G9c7FxQh
vDiqPWryWEFJp4nZ29JNtxRUaI4aY2tNndbvWDf7qGx7re8LM6++HPhSBCcq+7g86z5mjQsJJqbZ
Iz+ZRU1p1wfnJMsLL0rvVPsykU6if2YeHwdHkLnD73A0DdvGUw1377bpVPHoxjQkdSKkSMJMK1Mc
TwQhotlMc9lnts8FzhhomLpfQD+ffqYgejxeL7tFjQTVYdMgrUsmKeb5N0LHEe8AMntuBeLgh0I3
TcjWpS+uZ0ZIPeeZ7ifTA+56rgYVI6Y3u5wWKdaHLzwnkb3ERYy9nfXNSV+Imn7PObxvFGz5CKUp
ZGmxVNZ3d9TYvW7pch3d5XgT8dLh98Xz7btFLlPGJQ/joVDcpmw0fXvFP+25u6SGQI7MvIrKQnXs
9C5gSohJOtaotlQ1HgKeuWR/fGSJmzrui82DSDbLbxtLcmp9T5orkzfQoqgYLb52jaquoqgJLQ4+
eu6lCSnZCG527AdqLJPKqkLMn2JE2aPhkMSXSCHyaeXSP2EOZstC3ZuFpjmxgKeDnF1jtWtd6ss1
telbZNzxY7tz9qu2GOZvLL8DCsh5WHvpBcnwa/zbGvQ/DedK3Ucp3yBC5cXxecz5RbkL9+AhP7fO
+uqQcPwmFexUz/Pe6E/qBl3zgSpo1EA+p2nbLzLQQnCy4KancxCkHrgQq0ZksxEek4gv/q/ssL8w
bXDRxrJYwMz+G4wMP/rjkuoryKvPwn9XxQ/ztxtjnZ96owPA05saQQK7r9PzZ62u4JplHXV4pP67
nQzXsIM96raObpUBErUQLhBOxZr5LMkCekbX/jfYuESmMLlgaHonEG6PexNtIulDPiIwvAGXFuci
A0s3KnCNqLrycIFDb4xOZkT4tFqA5UPqOt5OxE+lPIX2TyWpDpPZJ9VZr2+fInqAoDeNV8xiYc57
eavA7uwNjMzsm5Iip6I67jvuv6T8dcudJTVPqliJbBi+8ZgC4hPmjcoz2bnPZUeyucBecugTJxBI
1Nj65oECdprlli3rdBpX3D+97gqkagiD4yK9/cCXgxaLgQdYSCZwXODl78hMPAZRP2XPT4rzZ6/G
WAxzt4KcZWS87VO7aTOlUCui/oqFv+4hxPqjiU0R7zE+byQXAs2YS/AxC326Plzf+UaLV6HvT7Sd
ox8bcJptiD+3VzmgKvM7GIPOeN+55JsIe2RnN2rsQpbUaQXOEwtTtvSP00El6Iqx08+7e/bM6xNm
ipTpUePSL9AVTFxaBe9KCiJ/ikFkpAdbLQtsTGxmLyZ6HXWljgcT/20lQ0rAf/ZwlOgN1s7x4MLA
Ut+hnQHiN1qo4mCsUC8CmkGYyifrJ8UAR1r3uOAyzy47uDqqSAId2jh8xzova0lgGpMnanAEKtUU
pVmg5xLS+PYx7xK5HeSRpKuDYTnBEPdKJzxSZC0jvwrrceep7WTul5EVQmixzWSP8Ik5oij96ezX
V0belNwvXVxHT/fr6TIzuR/OQBY1sx7g2Pwbz1+eej/v2tmPlirZyCTPKZjJLlbKH+YGDDR9X/2A
XdRwhvVrq+ZOImdbuBj+4Tl43I4XVP7eJpbAgsEJ83pM9NzXopV2sR/ka+8nzTg7XfP6RtD23R79
alHlv0grpoMe2uHFJR5lS3AaQcB4jhNcjIAlA8QraRAgQrK6IFI+44QdqpEMQ8/B5zD/HsRKqNbQ
UeIev9kSywdEtouxpcFzv7ZRkaYlmhKZVbmVX3/dCR08uwCzMZ6V78f2sqVo4DuKuse4ViGkBshZ
qDQxXpPWVoFaflBSepqlmO8bAPgtRhiOax7Djd0EzgpNIz0yad5bBXBO9o4qNFERPLZvl4RC4D3I
p0OAvSUlGyqiAonF/Ut61vGOCLr0qRTawTJjbeTbOGR40jjpBkkmshiM3JAc/0KhFENit3FlGyh9
W9vbHxJP9IYZXzyU5PuphCQhx3dTbQFLV9FzjPzK0tigHuanPlpYxUKEIiJiv8JmydJR7AcAfExd
ZKMperuHF1RK2RohoL7ovDY0mgL+VsinJDmGpnbJSztsguK+4joeeIWQvj36aVaN2jxMlCGIeU/f
BY7DOlZDrQbA2Do72laJQKio1mIQZBzxsHud4bT5kuaWSDYm0o12UWwLwCpEoHVtUeb+UzV2/fBm
9bXT/K5pFYy6Wqsx7m+3kIUXNJr20Vbzx2mS5Eo0dRXaLSRvC2/q/Uyu9vxtstzYY5LDxjULi+Vk
lOHtGi/5Fiy5RVtXdbq+dGcgD9qGbj80mOR1DvRLfVkDXmt7o+KKUCltS1VQzAhIG/O6OrAqg/nz
s6e0t0LVU/ip44Bk01gOgyx3/BruSXyPGkWS8oTa1cE6FOt8OVlcQcoB1o7oPGp6BeuE92QyRizd
uoZMRKONh5y8ex5GY2DGPSBH9T0CodBlcPUqSNj80q4tgKrw7JHldyYGa7Tm0w5taBrz1qCbL1df
XvI2nEK+cEOLosUh4NGxtnwgb9lJLz+ns7KCxvCNEj5FlGSWinwveXBiwEodjWIWqgLKNdlOUz8D
MgEuCwY0xVzg0z2P5geHqMsUB6Ns2Ba6DjwG3OfFH3TFEkQ0hn/rDLB2WaWfgMf5dhAkUNlAzaqf
wUxIMoElvNCT1Q8QazJFsc6xSauDTkNNT1EPK96WUzjB3uFrbeSIRGPdYDFH+uNXdN0SP4joephA
VsuKCB/auKbzIgm9VYZaWgnJlanj0PQ0VR8KyZaaKDKFh5+FYZpnQjDtvBRFzgj+H0Xx3FdQF8cf
T4LYvmrWfVWYC8SYdetjCS9LZmqwLn3LRuuLJTg/RFHOxk1I7umz0nn5aQ47S7f6wek1To+FbV6z
2NhqpHeiTMNBP25drLBjnqp78Hm+HTm/y8Gvog+tRvaqnl+7B6mYT18M3c6B0VKMWI+zl9VObnEa
Z6o4fDBvSsyBHcYuYx8j6aLGz7/bIae3mCvgtSECBQ3C6Ie+3oN97Fcsv5n6xEN1RQqnQAkjfJ+U
zJfDYKIfauYFIb2R33bx/n5NchjgADKNQGk1qdUAJ6YbPBVkhO2+JBz87yVvAVvuTfJc800filqb
okB3d/LIuleLlZu5qWBcBH9ERO6H3+Nu242CnNyoTUCh+zsDrvZ1Pb2LehbgxKxtIn027GOFHD28
iqYqMLAPdwnzDFu3IenV+2w2O+xG1VTvkcuFC8hImTcqZgv5/nfamtwkUd0wdzBx3IM27dVQ49eJ
cZiVoKSEpvrbd+9HUT/Q67xp6H4bYBpRRS+s7sPGVnTkTm0dNVcXR4xfpGF7IFsqar8d+Y49/FwT
Un/hnc36sjKXV7856iciwAgesRM6123ZYW9ckdUE2+riMz97lD9+jI332zVJ64wS0tmupnFBuZAt
pEOZP6Xolq/728TaZQlIm2rfErOrPKpZc6K4fLPPuJZkJhycOPkXb8wSN2OG5PxtHtcxS9Okg0jG
9Z224rgw4yoOxO4db92N1ZzWj7K0lvKLhLbB7Ittdt5LqGeYzgHCfm2AZi7wZ+wzYkzNU5d1jdEn
mVAgNpvPDXgA+yzf2LNqFsZhCUR0IN5kgaKtrh79pq7NMcYSl+eN6VlSCIM/qg4nS0zYRcrK04Gq
aYDchVN4IjllEPhlvtS8Mro2smf9PmE6CXITH4NLqmbjhRlwp24V2lqbOJjK4Wa2Rkmy45Ih8p8Y
KwXQSmXjyVzIK2oZhCKIJAfFIRiXQ/S+7mlAI5Dp47AK5b9BY+vlpRc4dQFkGv/WN02xtbHPCvxF
cyfaF+MMFPHUHoVugKlfTOo9djkDu++XN/GL1b/iPco527I8eBiqLYv60TN9Bn8nZhnpgKHjZgjU
bUAsFHNXdDfCtukF5upEcppoKe+VbjbTsPnuYcXqi8AKnIaMf34RTuezZN3OmJNv3Bc2tYqWaVDl
aQyDZYgCOrlausOChUyinHtx40ZgeH0NxhNFb38aw/2in2lvcpiIkYjEnM4YB1aBiiQw30rDccu+
fPZtTEw+AvPen5nQ5CSJJ5BSBnxN2ViWS6tLEZGc71aIfZ6iV3NytqooKuao0b/CwL+FWG5LX0kl
gz2jgPjDgWqYfOxc91oH/VFs9M0oYmU3D4yaM7kSxM6s7BGs0wq3Mt1qbi7PT3UYoBLEXpJeQPUS
RJHiPu8id+W3ewtmVfsHg7zHIPLo6XQjKNIYj9i9prNix/0DDmpfIuKtcIT+MhSZhl6BkIJ/BOMA
VfJNIm30GnLCoikGjU3KeEfSyfQyItT8S9XT8fDpK5a7e1aTRyPJM1kpUd+7xS8wnuCeLH1ryNXj
4X09vjQLmItB1ipas2jYM55Fc+OtzgX07Tjzo4AfaHW2FgsblLtoVHzEub5xcV6vK5+0clWPTVy4
EjHYdKhtil5/qdSrx/i61Yhv1a8SrAqspE6pyjVRP7nQD5n7w/pg2x3LSn721xw73Ctb38qmzj28
x8u9DxCgdrdCYj8hVwwPGG/uqt59ylwfT2ZC4sAKf1j4T/R6/LeMjr1baafQReC0jaOy3MDoPV+/
dkVMjjEeKBzh6mgsHdHvPmUFqoqdv1hoJVtht44xOCpguLJ2+LYBWlT48tssxWavxqgOSZzIsFvZ
loVw2moIF/A0XMTUQdQT4hje7FmmrR8yjjzy6lRe8/0CoRmOARW/RaBk2mX4SlYzAWGjAtwPa12z
LZccKuDqwmB6EIjom/H9XSiAAdOsweb03oH2xbmqx9fs+Dd5dWZIPn7SHYGh9z4UyPW22frgB9KX
/i2QQo5yT79Wzm0iyT+bCDEMsaIpvvuHY1W8TNfON/bQQ4DJbD88PH3QrWRFy3Vo3hyEm74024Gp
Q26QjIRf71ZE7nsQWoO8gXkQVV45ggGtNd9FGt9CkHoi9BuF9vnsBQJDe/Yf38xd2I0LtYOPh26Q
pDyq4KyGzbqnZl9LaCusEdqpkvPPTLm3HKOW9gteEbAekOdugzXHFuQh+XDO1CHYGIg8bPbANfNR
xyJ5P5iXZ2HqxA5+Ne1zgta4FuDNBinWyQYryy1ZrmXl0fb0IdK1eB57nG83sOF4gVHmk9grOxnJ
ulJidzgi5GFQqrKEstbUhw57YOPCc07XBxS7y6m5tk24XfAq0WIYX3uAG3ejS8GYKGtTZB3jpONa
9Adg0fboGocrjlGe7VuxnijXE4n+bEorXIBQfGjBmLwCPILTI6zu3Kw81tHVfcCcKw4EVbxjI4zC
NYkReQHo+078Hik64sbc+YpzzygY9FdlgRVBfm+gIHP2cmE39t4geM/qiFyKUQrr2jrcKGmHmyVF
GDB32onWQEsu8qLXNBeZTTEZ6vCN97Itm1eykCvjZNwaZsH7BtnZDYDLk7uI4DlXVxVvdGDcVQPr
YylvhCp4I1m40gSVPbsLaAPNeFmXFQ6GLFedGvptiw9e3RSfRfxjRFzt57IQwZLY+b4X3xNIrxd6
OQOaYTH+YemQJw6luMNWbecQifn9hTKk982P5XGGMQTf05VtP3A/cvYJO7V7rmHqIw+MXXJKHQR4
Rq70SxCZ5CiXWcV9YwXe5ZKxTM18HCH7iqYdRN8/3PVeh/msCrXQ0wkDDbNAUyVxeTftuHnl+nmy
HjEgrof6hdYCrbnXXOJdCAxtoGwp7EPhJnpqpaVVr8QwWVbf9P6AzM5pKdewZqndpwD4wcWWxtsE
CFbuu7NJttI85QmS7/+LCB9t/k1uUbqQWWqK0q9kOL6qCawrbRY2j0R1xVqfZc9Wm/mSzyj+kwpX
JamUA8QYWYcCFXaS+clwHF0ukOyx4XCzHhzK//14AEglo/FlrDgsTHZCRFIfJK19MIjVmWCsCeSL
laymkmWMv4GgKHwwCnS2Iv6XKqBHzgH4ZuUzLieOrDqPIYHTfTp//W9uoErAeA+T3T/kRcwbBh+W
r2NothGrsYgPSJBwDIT69HxfRyPfKvhgODkMB2F8ZLzqFE431zynlp5DtOpMQawtge8qGER08mdR
zY55J84T4OWu08UOxkS/qOhRJmci73SfabHUZA+OvHLJS1wAcDa/dnpc9bq1CQVOSinOXdAn6AlN
jWrUtgUn0oBtVQBKDtZf/Zmm59K5MHLhAWnFVgvOVpebTHClA8Qye+q/fsR6P/eUlLIKrpv0ylYi
mbW4PtqDV9WXd7hefW+NT20dLa9YhKWd2quCwR2YEBmZpEc6apf6UkhRDCAvRH7tLESox/3Yorxf
Fs9y03wqDaFvUQltODXpxrtjY0gBvWSb/iinU3ESo8JT2o0aLuPdBgSgwWEyNjQAcHKVmHmJ+R9d
76e44XW/1vLlIpOedqH91N9kdTmqnpxrh/I1VjD0vMGY5jNh9qbPLSmK0dQqZP46PeZdkiQdg5ub
8iihwDETl/mP4/fjlvmxAhqE4I0+ieosHJcXabCmId3ENLc/KI8t6rCd4KMtc+vZ0MHv1DmrDhi5
3CfbKoLmFL/+6NUxhqPYM3tiLYWPdvqabtfiy7qk59MeH8mOe2KIFzrYXqw044Amb6TU5s6zqeOF
WRcAD4GwaUiomk7yviLRLkS64yIekAH65S/kx1UBg4H2OQAXCsq6qXE/3bK8Dw//dLporduh80RS
+XMVem3DxlYvrIRJkXhk0XnobRGAMu3niO28Jl3ZjjaNiD033Dim8VFju65dX+F8IsjxwH4utyyS
+oEhSMTP4dBrBwNMIhQrUkG6nVW1pKh3NGhr3VJeI4Wh674RsOTq9o8K5AQ75XWRdJ5xlIvc80tC
rRggco28P3dBHfSc/hVUwNsmPM0WvxoFLjRKcxyYJRrNUA7mpo7wQ875yI0cYhDKFQqtaXd7doJj
h7JeJ+tRO7Zxp3GykAVJsxqfjO6FlbBHinlsUnoI3IXIbcMkn1QzpdSU/pfQJQTC15z3LoJZCcuH
xJOBiH6nj4VvfyD9Tuj5sZYxri503Agi+HR4RBgXfqEz5ZJtajou5TMeajdGlqHmkpvK0ush0ixq
6L3rJLsGzWN93D8DazKpjwy/hDWV9CJwEfsZIKVSIpy4CkwkpxnMDsf8ssIEIL4w927A0cLJ7xBA
sx/9YqB0uXV+h/MnEYvei+B3dU66gN/1pOa2bIsxDBKeLGvzI8AmWFUu4HqCGKy3xCeZgzzO4r5q
eeCX6FUYFN69ucZrqRW1N0h043VmqeEBis3QfWFokqYttqzmNcO0JzG0/xvM9NhajU1lmaQBsxI/
KvWU0ucqtPZpL7GqR4judzi3MldKGhXebvCT6twLM1TqgH+qmc4zGQmahwfn6AxJKTmTsxExRjrN
8xYJMvXE2kxwuiQKCaWm10Rn6MhKNtHDkF7i2Q+RBPwky0tFzyYB83J8/wTBVd1KXQ5TTfPDr/ss
MgHOeQ6EvcngddCNJ3R2M2Hae+GdpHGaOytMDVEgEH6ZimBYuu6xm0kWIAobgaUliQYU8ClI/O/b
DUkLtAIhwg/IIOtArer51zYu1Cj79kqQ98m2dn+5HVVeMCSwzCejAFpg2rapb7uu03Oyp8zircpA
aNFV6OcdcRrUO5inmkMr5Xd8UlDbmu7c7LWqyg1F9Y6SO6BefJ8+mQleMdH+tlsOt+a/BqOX1Tjr
62N6a/KHZMJjCop9cQyZINVhmjXiXFLUE5uq045w84iP7PKWbIR7nO0/fADR2l235egIK1t7Mmes
Zdbqn2o1nvXVelYVsU6SCS5gBGqMLjJhDAN0zkTXzFtHHGslfeEZk4J5qoJxCsIsXZ8gLLA0e2aM
KxbAfCJi7OFex9ERPdrnzuZExchbPLVwdgbpbfyXwDzVdjc5CxPluwUWNhjJvllVcCYUrkjdTHn2
b9srRgkJdzrxxyMJZtb1nJb+OL/XEfNSv5zJeZTHsHXpv4yU6/XKfwwSfql93QlZkNHPjHqeq/4M
u6b1qvsIkWa2VZaIgeEzJHMFCij/a7GnULBrxcX/HVtv1CbmT/DN28u+wknJ8vbdLeDHAKqsYHJ6
9H4T6//G+gNPpacPpDUSZNmOtsahAEeaG49bwYh7Chp3dbf+O+NKC68ZvlGhl16L8vKXtsyvy9s2
QEQp64jAw4PSBG+pmODDoF+eutuKMyLH4dn1LmlVnqSZrnq1V0JdWaUYDy5C6KiZN/oZbwXNKC8g
lXiRCOH7VAgbmgIDbow2nmBfmW9louZlzrdxSMwVHRWzoJ5JxPcIPy/Y4h+vz4hUTxIwjrz7/OUM
trKxA8pbS3rhB2M9sCk6OHNYxYaNWN/5SXn8/SIJnuc7mHLdD6UXO4OlWiZAlYOTIq2P/+t/9bU0
UVAUiG4wSOsz2y8EvFYhqUArJdkd+m5n1gNeT/03ABaNQG3BqpESj1WRwW4BJO4mktirfvlREpiy
TzEKQ93PrcUmeWd+b29/iYiYw8hRj1WF5no1bFpxuSMPpfzAPiXpPD3FP0vZCVFunQbhuDjeIJsq
b6nIWzALxjxzRddGuRlIl/q4ubXvUGPZ2LrfAliDqrEEK8gOCugXiq+sdPOpgCZtLM+w4My0l7iF
Ur57q/N8NV/W6IXOuhOFHMOkZ8ps/uHQ9m3mRUyzJwH+Zq5qNkZm/0aT6VhRuVR9SX1+eBtJiCwY
Zg7Ta9qnmyepmZWs+WNSXTuNlrl1MussBsdrXw01OZQDpMeUKb7EXCbQ+egBeCrRN3NAQp6AbjTV
Tr6vBB+ebwLbIIp5FLTfxiyVprEXxmzGJmJHsLeBiJLhDDLRs2XyCGUxh1HwjLE9Yvr78tYY6mwF
x7bJfttcTD71b1L+BL8Iff+A/WrgUgaXyU+DlHmapgFrk6T9zSLMhAt0ruj8NAxY/tlFBJ8N8KmE
h4XevZ8nlDJtTWCEnPY0WmzSvEx2oqVAHx0oP9Ar0F4BhujF/ErTdAhKCta/dPUtgiTBnwZcspi2
XAt8BWWM6yRo3QNka4LmhmY0NSl4wOvUHWqVwEa302q5YCd8OMCzwpqIj7VOrX5WwE0aouADYZfG
r+QYjDdUhXTsNW2fYoIMku5739tRFi7pjF2at1oRAWc/ce+BclPCXGt3Zsd5ddHjsMzWSiElbiRG
8IbfQW6mUN0xqwnGovhArB2nDct/A6ZWWPR2MpkFKtjFHjjzIG8P50ZK3dvTsWuCw85L6VOPH2Kj
gq5uHpGH+qcPmYh9na9ybh0/8OfCJFBJUFBnlXFs5zETe68PE9qkiqe/qNmif71TZ1nAZDrqFY1w
Yk6BPr7dKt1naHgJyrMM8LD/t4nU4fCYfkBghYulEwlNfNeb4drAnvCH1A7CBPhmvdgShL0nohUP
raJFXv32W7aCPLlsT/OWrjZfQrl7/fWQIcd31iiqUFSJ7PAVnQu4n3HL3cQ2iZtBMysqGsrBjD6s
+9Y8IXam8XR8DQYhT+Dw/nRM4h+/RFHNR5CTcPTOxC/osfc9HrDwIHY4wkk3FHFGnRDhJOZl/rDj
o4UwHFM1VQEgDzbY4XpeHkf2PgwKr5rgx9Fdg8DLr0loHxvfvbCWvCRlACqkvZi6Uk0bTooWRFwC
xbxKcVIhteD5RoA0jG/IDICIaKEVDlSGzgu8ORYaZ/a3oUKUQui+CH/xZmCZ5cCnRzmshYv4gC8f
MWmvAd+3PAKxvNnfkIZAsFdYm5d+/o9ZqBPp4feDloNI53RE3ZTUYMEQWAkbo1GYyCmI2AMH/05L
/ZTA36cdlpgHawbLe+4K1SRFRWKl5nSQmTWQZdFoPFZ9qzp5YtWQDYbEGT+ISZPL2kNy6ad5Zbn8
DNZcU2u4hv3ixbPVyV26NTKh5tS+/UMHT1ynU2ISi9TUagqSMKwcUGs7fnfQpWGa8LS2g8UpylXQ
VM+UiIwaQQt+qbQ2bL89sCu2O+81IIpFlOLtRsxdV5G8mHdici5kYNydG3YMrkyOlYsSrzH2C3Uq
pyvPFlBAecfC50Rvj/1m4akUNfeN7vL1kNpOLm2F2mJQxlRIBLqiLOiIeuTb8qjxc69Y+V2rK+Ux
dDYrp9WlNIrubYbzdxytvj8i6/EUx9c6LPbgY8r3uR/6+aifY8W99MEPlznz4D1TjGzya6OjqwT9
dufjNoWylthnJvLLDV7hJtdkfibQcoXuSQZsemXAf+n2QZU8nG16lNwxezYzrUSEY7hiOD2YmA1i
kHQR/6J8jMZbH0bdoSpVJnA9ql4naTC3Mk7utF56T5/9H14VdnTg0FPOGgK2CJfpXYyvDTSPqlGU
Ju/oruK/7D4roqovQBTKomwBcUxWZ2roC+C1BC+RMi95Yvv8fd1Aw+9unH3FYLooONsGhNIGGulV
aGotiLDIZZ8PiPBmmWf9G3+uqrtp6EIyr0tGKQuhi49+RR+31+rPxjfArU4bmmizH8U470Dpvbv9
H39Cx7saNiTb1IPcElBG9VaJoo3Vzqf9AkZ6Nm5CE0uKDxL15ngxhSbRUvzMZfF3QQsEItNnMh2l
N7QEwPmzAYhbrGvlcGsjSuOw3LxFNN0YGN6/VWvVwQXLsTl351MT2X+5flwwCoxzX3KmZshnESXK
sE0ARXo07HBrfanpskR3nXoIG5kiDV2v40RMEfWNnqGc3jXUlA1YKCc9VSy0P7WV1+/bwu+0P7rO
9k8mYLrGT1ltKIoPBYA/QUgCyT/V1Ea0Q+ziZTV6OftDZJbiU9W5xKn+UV1UkecYx48G1ndbcBWS
997h/4GhvLP0bJ7QODfAOPz7XL+hqVB7K4gcuh/9qwSWU3U0tfWOKcN3EDz7gd2ZUiLRWggI5j/4
vw4nRAWcKAGiWyNG29+P8CUM6BwyYFntcbxXisaIlNXZmSCvSxr7WEBbHlZIXV4Jo2Mh3UXtHC/+
J44U/58Pz9shTEaV4oEIAp0huVfddIPoNXBxahyEPLHJxUZLwbvuMXIZgoXF8nL/bR57rvnQ3z0l
ceUoIw4zOlR0lUq+lj6oAOyIuQUItJtKnvhhHi5j4byXFO/RouVzMUhESUPop/AeYsZfd9T0hk9w
aWVAU3wke82lYUvS/wY/JR9+/8l0CShIOk1SgWGg9jFVTtcgBemN1ZhlbgoLWWmo2P48JA1O2MNf
zz9QySwKL0UM4w53oxw4xlzezo80YzS+aImShCqSYG1jususvGjSjNIZtAw1QzI2X6mvgOM+9L6y
KEj40W9+pqwa/i2kitMKGgoz7+nmniqc1+XwVnXzws6ErMwQDoIAWzugD30UuUfJqN3B30c6y9FB
rls77XYv6btr+Lqo+XyiRNUSVEfSeIh9wwPluimxslMosSjwqpO3MWsEJrSzsb0VfeRDvt2BOrEl
E0nCUZjtniyLMl7hj5LwPA0PpOJbY1RzOrydIF7ZeBW+Yuq2oNi6lNQD65lWCXJFWnFlCvBD/76M
P+OKxZjrEZ8OgTnrkvL8c8mf3bE2FMa+KjZrt+3mNSs6F+DwvAnTJ6Bo+qtVbdExDhTV852lySRH
tbPCG+HamO0R49VG8c+1Ah9YUfYx+ZPfZJUx0OqbJUxjQtSsg3YYPzrM0vGa0tSq9o+an82YX/jC
XqbRMKx5GHCuQqvPE4Ha/wp4H2saWf6EMK8mqJ7QoZPP4fZCv1NB7Ij/mfSTf8JTf6KVCgZaTlsK
kknmQiL2df/lSY2BKtMVrXHWQMvNefdxIzbfur2j9lZKkr+8wG1Z+2c5MlPNDm794xrPwgsha8Vh
PibXtdj0o0kAv7DDJ2gPYQSnVmraC0HHP5ffvV4dIshHEEQ+MzPXx481AjuEgAoMK0y6adaT6lPr
hNouN2MreAhvzty7GGpS/IlFLnMhCTjsu/qxJeBsKS6xCRDxYE1TT37P83UJ39VLHYnZf+DitWGI
IPwskpfa1ld60HJM/JAEfHxVg7vLwocDZaLMuq3c73+n8FI6tzdXHeIyo8pELse1mtqD52JrN/6E
LvIN8c4ff+dEGhdzZZ7DrKXV1g433rPJ3nZErSA6o00hB1TSqj3Wl1/DktyuVpX3WvV7oagwTfow
ehRIPrWzC+OOw61PJEgSR7PLFzvXqp/fTvGv01IrE/wD2qX4iiGUXMD8SKHJ+QC4XR91zJ5u6Wsy
8GDg2/iJEXF0FStiq4R6Iyzz1vWhLKZdXO+pIUrNP/OuwuX4H9xjfe6QYHxDkBYoVPK+bSFjnWMB
cTqUcjLRhOYNfoGjekgJEDPbv7DY7G82FWnkDuusFi7CBvRXVExxOH2CWZpqko0iVPeyvUcnrkQa
wScijVngqLhDDfZpIkpjwPP0SHS64YbaqQQbYRcqXgAXfVco08mf2tMpKhs2KqKWhOibr91ta6CF
7YPlWIPSuoAan19hxrpytGofcJkLUx+93KoF+4cAUzl6D65GmFCYnrKLLs7dVVd8AkGDq62bhXcs
TxkwE50IWl2ZKrYS7zlW7pz84cuO+IIwPhkiyJDgj8TEhBX3A4YMT/QCZKdLT4ht+M84tZoSLwTw
TksU5E5cH/0dn7MDEHtR2YEV2LckwQV6ZFqQOo4TueEVlKYIdUFmC2xeUdupbiIK+3B3eiKhugDS
jgoeECqJuMZQF0z1IqIOk1D7/EpV9RbJX8RTetSkOPvFyfdnZoon72XWHgGRaDopSV1Wy5AKsjpN
9zxF/V2zZQ/6XTmmghCclI2zBOxURMyMuAXc5fugYkatT3yVXOMSHS1P0eWvkY3vYI50LcPA3ke6
DA89Bl708pm2yzB2mz2R86dLLMCBxLaO6bR+2JcL3VfdjAxJWGbpx3DXcFHbAwvBByOH3Nb6Lucn
Tsu9KLoZP/x58E7L6lGQq0f1kyUFiHHIc5diRcIpIhyHdENhpuepNW21Khq5whV84++jyp71WzoV
xBhpaReSWTb2Lr5/X9uaP1a6/TvASbIguz/sU3pgF0PLZR4TZ0PA3pWAbqANtJrrELJpQiVn3Qm6
jsolBprCVs8beigJbr4VIdVy9cKeru/XC2AjCGMBSTwXyLZpbaq1jsnja6lAG1WHxyAmCvIrNZMo
XsvPLH9sJGnwJMtrL2oQy59NWQC4TDflq0ndn/InDv+CE/SO7S8Ts3+RLreRhzRKdjNQXObn/lqR
N99U4jgOjsWgPZEXn63GWYsvEeaSmOZ9nbY2t6nFa4y2pxNrWX1TKa98h6JW5No/wi9/q6c2LFYF
irPtkwjhkWTRAHvW+eqeTKH+1n1xRubbYqhaLFsfNjSgYRGQnNaPFc32rR+RWU2O4gB+eHqHsxvb
kXPwGi6ya4C9Lt/IhO7F8yDFGRwH2BxUON5waiswxyFR1EoGuCNBm3ykaSM8mejOa9M1Fgznr0J6
4jTGeRPszaqDt0jXymmL50/6je3HNPoaTg1JiwFzvVwGAU9c8XiXfV1Mc+xEzrGJJnxJZuPGCVFu
mkRMpMgHyADFNMa9cJ9PmZzhqshF8B7bIPZLBQWJk8xp7ujjDDWSNvRVwBh5oQKXHXtg8lLjQ87b
DHrefLh5ONhfuBgQ9nKQdRZ/AjvapP/2qAz7OWo3sjffUzSiMHv6SRgU4KHMrMbpAZnkRqn7rHx4
hIF6Pc1vWOZnAvTi13+8sw6+h5+SKcbsAcMoO/EaY9IMOlJ0+6lhHj+88tMJRS0ArA1x0C46/vli
pQaGwd1Y0MSu0RMJl0Cz5JV0cD039gVw5DmzTUbjVzEQM3CAlk9JxGxNaROv9XMsQ+Wj5ZGaFIax
Q2SM3q7abjuAJLn1q1+pdX+osndSmtSEbSoBSuosHf9hFRFcn5LKm+bvmUB8N38vhI0EB5vbxBvA
ZYUtMNk3ffI3WCfKGNIt9t1EK7rAaAWqwhizzhRhc7iEn97LAChcKfUGC2UTdyPDfrw7QgEpYiwq
11exWZwG207RvjTGAHAKAKMerg2q316dv7ZB4cUuhjqpYGzY706MxweU5mCuYqRypneYKpG0qMni
n5KYxd0f6/xJtF9J1yXSU7nMDAAGaR3O16mjrsuEuCyEGbf3qCgShS+0CICVhBWsluQYHubJcW6X
hETvhQ73CLuKhE1HKr/uO8I65oa0YI54MjN1WMOQ4Uh8Wiw8UuK++GHaw6yN1bKC7y7Ex6VTmWqR
JvaAEw9TbrAEPiBz+bYoCEV2HP45tVK6gPg4VErY0SHmOszdrdur+RxgMfelYeXzHTF38eJiAFJi
Q1xbYRpT8Zm7Fi/1PaKp646VwM3b1YD9dplZlzfjkeDNwUAuef1TyY2JGA4ky3uQVxHYftTNLa7B
6PBcuKnCsoLF0mBxLGBER4vthy1dfa58pn38WzPo7ZqTko9qwqKvCCel7/IW2b9b8cWsIsfhAUHG
IlppJpgNB7fDwx4RKkdnV13gDarodbfAYQJOmYxjelhRioDguyGw1OSmkvaMwqtVqj+d3ce7Sb69
2HfAbBdJ+jmA0hkNUoVHrWr6pRGfVg25rUTt6aP4gAlyIO43dMalLCgxBJHr76ojr62Oa3YGcKbx
FAhdYOMwkR9Q3FQNMTvdIqf8AyOvnnDAWrVTnSaWzCQO87zxnXhvW98pqNtxe3mtK6I1TiM1teUI
6NPRkdIdu4qZEMRPL5mt13UihSUkuJm2Jj9gkmmZq1HTz4f0ovG/lYgIXG+h+lyZb7VWLDUebGnB
ocuJbHDA1oWbqdxbQRDwPmrKActfr8r4dwJZTRVeshmC6nwgTdy9ieDKGP/GWI6gHcz3nfhmoG39
n5EH5RgM9QGpbVVRR/DU/KpdaJTTtBZKesihjjjmLLZBocnICr1IlckocX1IDCdkAqhEaugu+PBs
8pvdDQZlz69YAXNjyBkjmDvy9J3zAlw+ZGmVQhMPtJLyFaS3w1UYPY60jYgdVsxQgnc7Mq8iKjgf
iffU+dg1cEQfdGHNnS4nlGWkKpRIwZKs20htFjruJ+HFuw2+MiUYxCYq3SHGPNMmkK5sKQDMaFmJ
AN+7pooqMjHZabbFiQSGp4WXufXKu1IU6tcN+KutX4s/gHV9vA1DWtugSjb9yLBCz+G+Yo7yHXop
SiG5Hdpe0BgNt3TltaFvSpE/getfKm8y+OZVj79kmMkYErzqDZYDm2PhiG2mnDmoXUMV2iWvflWE
A59ZSRESAnGtrcWtYAPAyMkOYlFAg7utuP1CVrlhiMJ1ZaG5byD9r3KNwP4tnPMOqKyfxO0AdK/K
dg/diX3g3wtM2fiq14ZftBn45bSWKVndwRyfhN5tnYovAcTZqDqIwYH76a0ipNcAEpu8+xAEGAHE
VDaNEb3SGF+kZjuxb/BQwlUBv+3HJR96kL+E94RnAeXtjcUemMpLkrJdbobLTSbZbMNEPEGYZQah
sWO4uiZZFTb4HacRwRXvG3/oFFXQXWZdpYUzPa2DISCP9PQ2pLMXWFWxd42VxGA1jrlV0cjJEaoI
5Ycp7UVpCxxFfitVltJLBbIT/iamxvkVM4/EVM50vxlMh/vPmWmQz7iuh0Vf2ShD4ttKEbI/KUM7
oNwkQfqTpqzaAAo5NR0xpOtnGnUzpHmH0zU7wqHYKXcHQfe2yAJ2TygKVh+TeLvRAehEKkAF95B4
V8rlxQZwhKg+oMVgZ6ks0Gc67Oj2r00OtVpO9lD5f4BpPxRzXKbJ7aPLIVL1WSQq5s4ml/5cbivH
GQNH7sOjXWjQb2d7uy2VnidF7EJYI7CFlwhCCcffKNStOqdlhjWuQVnAjWRATqZBtpxLnJxt3zZf
VnSZ5lOfeEjIQNVKU0Oen7QiqNJqOsp6lEdY3aRdBc1yK+S2cZZVQVajzohjUIwBi/1szHr4Gvm3
Bp60EkEn/7ujxCHdbwOaProixDGtxchJJQQdFx0qj1IWGgv9K9LbKKbbK6xEtzVGsNgA2vcznP0T
DNzbR3drW41XH3Uo3e7/iUOTSTawJWR8Aj694GbEScN/zktuJzG7Z3dr0ABg3OhY7uFzB7h3iAc9
T9UOzpJATLR5lls3OKLvp6kwzRoIevSWfMA7OrM/JYA6wjYInRxt16cLsph4xXo7S781ro8VS0Lr
MYdoTK6k0iezNNy1T+ePWbljXKEU+wBdaeeMmJC6xGtcU6o7ydqyR/hex0f0JYTN7rrJjP/Wk0Yf
0FcNnn5QwPkjQBw4CjFbTNBO2ZEP35FhnNfxNfTlGGd6hDBQ7JTLKUhAgltYFhLu9gunIRqoOUg9
fbkTFOjMV3SYEbVfaRcPXr5u0/FoiHLvjXjVArIp6IYe9K0ZgCg07d+yDRjwhm5bNRo9kSIg90Bq
oKem9OzziNrExzTxQIf10YtlHcwvexwCp8ABcJfexx+ouD8HRB6GlMi4V6SAwUpynC0ZFdM96n9G
fL0gFfAaCWymC+YCWSJxGAPRHweE/7N4ncuPK/Ys5MbgclSPQ7oUX3Mu/PZcoTP0IDqo9R/5i+cq
Z0gpujIOGQtICh8N+W5yxpeME+fYPL8pr5TUsp0gt/8xhinlD5XTfgSKZlI4QndgtsgEaerdfWEj
FcSq5sIZlngS/KEJ9IV8FqfwRwyyZHmptAA7/ibSYotJ0Fuca9tQfoHDXxjELGKd7yPKlLQAZ4X8
TdKVLw8LmPLpEs4jJsfSO66rsRqf2CJihIYANKE003RDOOuQrRBPz1mtS9VCrYWU1D6FEltOe5xs
w/cur2oN+Eso5V+PXIubFwAQm4d0+ZfTxP5hTbvl0VkraVPZmxl/fAbzepHwPL5hRnqF8Kg7JhHc
7eFzr3uvUdhBf6G2RbMg+YnIHZ9BiWVmuNp42GH6EPdrW7C5AWqPNwfkZTg807WeA+EuXzMkqSgn
m//foDbXsLA+tNcjqAiexYXjPiVrpjpe7EkTEHtUZNQCIlNY3uJfky/ij1LUiiSCLuKE/MkM2ZB6
Mrt9cSrBDhvHxZVqqJYzJULIxN2eNEwy9PGuJ6gL6iCFhXRtS7zOw+xgpxhrzY2tUixBwC2V44fd
t9s0qTvGB+X48M2Di+yoVKh4SmSsKa1H+9STGemqSd6Yrz2EoQvqhNGOnsuy0fAYlQ3ej0mLMUEL
M65DoeYUytXxbNa85HMMIpcg2K6NCzthJxVnxqsQJ92Su2lbFNQZ7Rx6YcJZ2Ja83XYA0G6Xd0Yu
HkZA4+mrtercmiSu4evsX7GidKU9OdlvlrV4/O0ljDcwjghPswou9BUvRhWs5kV1CwKzGdMe9UC+
F4XxM5GcxJ458OzkwQgTMG/yK81wlD/EmcP299GGRACFUcutY+aZrWsYJ7sJ4qhIlyQCb+qPISaY
IYr9ApBxIbD0tv0boQFl//ahx8ovs7ytyTB5hcG6H2aKYpNJt2s0tGhKAYn03dIyecLL/eXdrEKv
Z68WdQRQo11n/Y7JWsWm1bXFfj8lC2Vlc7guzLdHKI93FPFviCLrkdlEAU0ViwjHyM+NZQtK4SpW
CiokcsONJz75Cw6pD5jIQEsbntRUeHhjLwRgE/0WvixvtgKn3m/bqBoTA4rPzCameJgCHebFvF/8
2QHlJZ70yYBmbWMSNT/MvsCo0orrmU63fJQIYCBbprnAuDM1DgVZpyr7Hi19zYwoHe5vK+1Dnsd7
uKtFMAZnZCcm5DoSBl5lYnR4Mx0yYrX4MVHdevhyVTiaiBhVhQoy8jrmFlvC5JM2/9o+PWLWr/Z4
iysgSWswXl44gwDP1BdC09rFaV34WKZxlYjVlZqeZK0sQgl7HP+bJNV+HA47Uo4ScbTL/GOCuEg7
42P/n5cW2cfVCWEAiyeSmuUwG50JsMwUvdiM5AIdX/GWUWuV512c8JSPGQFCK6tIpBdNzL9/De5z
DnVAFw6iCMfGiiIQUPpdJm69jhR88xA6kJaZv5IvVcijrr23htOz+alWR8jLqEhfUzaKpO6+W7IQ
9tqP8J5r4eIjKRAda5F+kvVsXOBYNhuqMX5Qd+44whuuQbz0bjg4cXulN3N/fXysZu58keEDOrAN
8G93dU6uRX/whoHPh0/5+7k9csTDB2/JqVL82ZVo5+xgLgEbJlSEkQVYekBwm8ixE3qlUOJ9Qe62
1b9kEVQXSJKAR8BImlscdkq8CbXhvpin1mm9zbcqQFaDlPrLaJY8To1yeEH09X8H37gTNiM0J2La
Y01LRtlqEVdPBB8tUvj/Z9YI3egMPW4X8CO4yT9phdASilbuDou0Qshe23MbrKqWHdmrzw2aL9WF
q2KyL+o9PN9gvnRbQc7PnDtRn6rIU4HGYVHof603sddGyi79D1OtlHdTKe13Rq1r971ypRWtqntY
seLajvrHyfTwHEWo5zkoRhUs5M7aoyJnPhR0Ahmou7Djz/eOyXbAzsxi2DbdXXe5ijMIptLCn56K
3Q+G603dpbjwvoQ7mMJaF/grhmUnqKA2KJdaFVlYS4aaAlkgoeiCIJ/flz7FUev33vo7VZVcTqf1
OEPXgEYLt9ouUVVvdSGEHIrhKCGtGWUiMZvDMT8eteNkl2bnHR5gz+eqvrA8XO0s0onjYbT1uCKh
sQwbeU8smzJ16yntfMjPg6LprxmlqKZhCkS5X0tO8YCdGB7mP8lTm7ffK/l0ZfcOGATppxHdDXqu
yvtZ9FkqXxcx7GVi+CT24UNruGVhC1gaRKJ35hN4pf029IJ3OS4GmmdxgPopvTZSllP7Y2eoYTxO
GWMB9LYSeiJs4PyzjSmGD2DtkYi3J6QYGgi4NSReKwWDNkjbn6HBqYcb+jtjfUp9uHWWHvstmMli
nqvXYqSxaccXmezXhJcUZttAV6n4bTPjk85qKuaWW7bheld12KuFjaFFCvV2elfcRrVulh4ONNeY
o9HY+idbcL1roEfr7hXpK4wDu7v7uq3WwqNs2pbw1XscPIkenUZETQpasVFBm26kAd0N3hIHYqch
ZMno1dmF3bOJMc9D/dDamdiNBcYlJ9YohcTLeo1Buh6PchzST6iJexoUYMktOPDrbUrIUxneLKB9
ForFEye49eQ9TNEsyjkhNDMh+iTgUkFIJ3mvgyt1t9WWeCjh6fZGMxQEdkR1ulTmS+zpGqOXjs2h
86MGMe00ALb0szF4kM+tPFO3B4ftH+6XsbbrmzNZCgpWssV1UsUjjsCGowb8f3tic5Kxf2libav1
8yqO6T5OljhUXqiT5q53BQSAL3BYDRkuYXuw7MUOGnI7cCsIzujj/8TwTvdr7pmIczafOQZ4caIe
h9xtCoHzNAO77cTQnRXIIR2NyQO5mxzIj6aJH57yMSmfAcOMdS/+9hnJSPNc8TUZHgndFB3SSPdt
I3qE5uhguvfUFMMivzctIM+ddpe69XBnkxJrRo8Xnq+5Zm4NgRQFWYg0I5KLIg+40B9TGWRtN4mi
sIe411fKP5s/uAhgor59ezj1DSEIXG+s5jMWQK3IgI/6+ABghxlEfX/3/y+ylkFWnjxobkLi7cWa
MyWskvrVAkM9fJm9qwPYfucjsjInG+AxS87asg37qSHI6Fa2MPONrmkzGb+eSPFtW2ZFvDPFub5g
Tq7McdZiYGvBJGHz+/zRulDoR5/EvYGgyV6y8Lj+45P4Ne+lrTKP2avK/4hVUYYg/siCLU4wH4PD
7CCKOrK88dgUOcYIBaCA1KwPecvOM4IjTBfyy2fpHl+OEg8XJJjGr2UpAkgZ5iKSI0GDCcp7ZLD3
rkcHn8+2Ux5iQlbb+G+poRZ9uVzUbzh2Xd1+ZS/0lnCSU0iLErx1DGlb9qE1/nOxg79FQ19OpkFG
qWYtUOCryjDKTqvRMcpa5Kpwx91KB057kY0eePRugNlmZnlKDP7MZBW9YE+FSXDP7jkWGhTZcd55
JhjlBd2kKjY+jsngfpHuvVi79vFHv2MBvntc0PlA/bJN/Zjs2sZqNrudEBB7zguQcDiIK0mo9Lzo
S4JJ4hFM8JCeX5hsxk+j2no2yqtB9w29d326ihnmAAMYHAYmmISplyDNXj3g63gqXAuunH82Ks03
D68w+KDTBkoRI7sfh00sMznuxv3rJP7pweLTYKO4EsPqt3WxRQ1szG6GEoH3wuLQz3Vf8Ii/awOc
duMfz7fp0dC4fv9r6BgRFFJPSkmuPDQ6Ncg/mTuSLqXVQBecfkEjBNTamkzB13Koht/g4B3zYAId
MeruZryqALk046pHoDzQGdW+/XdiL7+oOApXQ4EUB/K1FpwZuOlyFipken1aWiv6eD9aSA0ZkXLG
pCWSo6quRNB03r2kZPfHawOREeeJ9rtBRofIHIy7XT1ALRRylL/n067/uEYw4VQNMt81RZzEqbqt
fDSdGOMkwhEKZmCGk5xNZBRouoPlMoH5f1+kOOPhl1KpvtHbRj3si1hpiwzNHuIRuOGOHokQ9ak2
2o5PXRhzBD4Fz1WtWYph58pb++Y4o9bqCKtLVkanKT8zIaP8j0koD5o9iorCKDz3YDgzp3Cb3yIz
Ru9hCCAgfEPTYIfONtWbRnrB0gtoqqfbwGtC5rvl1j3VxawlpbBAIQUFCyi5dL/8TkB6ur381/KT
+/89C1ZyeSbHG8VzceJb+ZjI8fbzWgeNUNf2EzlKjIxAVz1e2+PhnmvmIdKvfBvuUkf1tnZGEmwz
Kc91c2Us8AVBD8HFvYhY33/+EgmC5gEh57yubMVXWcy0c8/VwumGIx2ls0xnJhml5yztxHsyHTfE
tm2Aes3zl3inDcVk8ZrobeS/up0hU2H1Vcsq+Fca5USgVS0aye81y5f5r6d6QllDcITWDQL9lumY
rrN78lWS5Gz+c9i5QEn4ftdFXHksgWVYPkL6TOn3CjJY3Riwhp/DGS8ka/Yz4d3HuJx+X34oEVmq
IQ2/E0GshlLU9nRr6y1qox0q9mtibe4b+FhEAM3W5xzB9u+XrTefL2RDCc02mi8ud0HyggKuGWvL
mFC3hPrl/kcZYY+1TIq8nv+dENPeHF/sFOZCSnsPnIxMb14/IbV10GGR8YARJOJ+arxY30ioOzmo
uYGDhkly0BRKrlcQQ/BuhuwuI8YmK5rRE65jiwlKaddjhXgGimIdvmM1Uu4cvK2AykKe/KIhGFEt
PmnU/U9caLaNnJm6BAHd/ad9DUBOa5L0gnu/TVYaxgUOQkTiJ5FVrLEdYFTKCxKh+D9Ovax5BS9M
g3bGMQMgsPvixD8aXcQEBWngV+Ta4/wvTzrVyNL1JJOvaUninps4928MOo5EN4mvora0tGQpVAUn
bUpDC4FBbhWoHrVBkLo1rH1Wzu6UernAWs0yZrBmOpFv+TJ0ORbezJ9yQsimWp3gtEiqPn/8reG3
gU9ld1uJNrM0DqhtEQTd+Wsv8IWnMdlkN1kKtO7xfEUGrmS/plmWnqnOubnnbXtH5buipoTMbhT5
2xUkrP4NLP3g65ABfDVe7LIJcb0gx0UNznDu2yX1nGRQtjo6VEObn2IjN23XpIQ2n4Jk24ptIxD1
iSVqDzzuffN9wp1rGFT1TwhfWxTZsQCWq8Dy4YTYLj5uTguv+43FR1z2QPg+9Jpt9J3ZyMzAG/jC
vE44hRNt+4yvHHS11nOHNeJ2Sl5fue4xILvf86hqFSXb2KLYEF/PU8Uap1GRy25cCCVdeoAUZ6y2
Nx+AwrpWAtvc0Cb1ba/lWV6xQFREUsREw3bfbsp1ZQCFYsp2Kxm+4sOCqZPqVXyTMNFJmNNh5OhN
2JjS2A+yCN7VMSMuXaz6Rcj5Z3+ywqdZJavgCByzl8K+RiV1dBFLB3vU9wy5Ie1VpIIYpgbqNJbK
H1+IEnlb03bjToxTOn7GVOwZmu5HTyAx6Oegbl1oBKWo3GQsrazYFsSNbyi0QSX/cRY971YKSlkH
Opt0lGoSw4tazctvnVE76BqpfLuPtkw0tNv99NceGvHuHSaPkOgRI/TNwxGT+uUrI763GclzAHCs
WJJxgeo0lT+xd8JLQlZ0fB4RjS/TDsUhKpdRO+RH2JQzS5FXaAG+OtZ4MQHSNtzxMu8eIFtmXWJm
62rWz9gbLfSRvQTHOfPQuCsiNrIDa+u1j7GL7uWme82PE+CYWdpPCwTtfU+DcnEG1F1QAzZqzEYP
jBtYMBmvvQolKzvTw9fqh1+gCmYfnBtGtcQ6ZG8Dkld/DFXjY3NBSwCVgSRkUGTUIiCZ8soEuAT4
TCn96iMdm3e4jk8mpAUW1yp7Rnrib/uF8Pn6qkqz2p+GCLX9x+DDPLfB7mvhtl01grS1a3JBOufy
5KE+xiSv/9mFwkHmaBvYJQQkODCaqQ1gkHI2XiFAkR2jShwNn17IirlV9MGZsv870OvD/B4pjK7d
0yWgPYYiUYnqPXmOVBnk8LTTEpvRnNQUkJ5AiDt2tlD2tR30Bv3KsOrY7PRRZRrj/d6a3L33a7J7
ZD/CYx/mPJ5AlGbM0GQFmL7FJkzF37rqdlTniwkCj+dyYD9pnj+ES1+N37+ExbjuVOWNh39VxjAq
qbH9QxmRiigK7VGyLpzk1MAxQFipi0QPOMGig2jp90jH2EbXwDLxe+zxIqloAoeYt1nUTQZxnHn3
IkbYN+5xbYTaDGEpGceVrKcU2UYxF5xzlWG8d+vi7sP4+1m53khbvXA/iu8bDGBk4bPLK2tsuRw2
FkmF6l7Z+e4EPVLzibSbqJX8Tky+nhfxW1FqC8a+Vx3Q8pr7hEVMjOC9mJ1yC5UXcTkeKfkZF2ta
JUUQozIY1/mZY+1GgDw5Y35eNp1akUWpbi/4RJCTToZBJCbBeMzinXUDlkBCHfmDo8Y9A1tbmUiD
5Il3khJkNNmaHY8F7AbUwqSw/RqjJn3fWNyCIN08zUWijgWAtkDyZU7FHKq8nry1uOWsXR5BpGN5
vhGMliII48gZte9F772QIZHxKj2CZ7kfldBfLR6Pt26odC/cHlRvaU5Z0D/UREUxoadNjeqTU9hD
moxr0EUthCya9iAvxsEt/2n2WHqCGnYzDkPrFoY2tPFcgpDYFGbNLjwERfAD4WvA9Q3rCBHJkAna
PjGyCA+43P3AbnfEb5oTfhH57fH9n6TAk4PrX5qavAvLBVRkUZr3thC/dovCZOiypxwFByde7ACk
rB60Nj2zVpGA5hAY6CnChr/NozIBqFRsj8YYFY0LYTwesYP4VkCcy1mYWhDfQBfi82yK6ShjU1Ca
VvKGUQ826y2BqKARpu8y533PUu05a19iq85HGsPDxKpiKsoeLUW4xEcs71rXIWwJcneZk1XOXGVK
Wl61kR0A+fzqnjWFpzYv/4FOMCASgwL8/VbrobVSX2Gno6h1UhWwgfZz4x4Qz8vuZOzrJsC7/RQB
z1PagLZ2AG6rsDjvTknVtKtWweUfw08p97qZyCXe7Y1/EY5WROKD4Psa+D9chYK0YCfOjaJx+MTT
yRTD3UG8ibN85GraNITvALHVv6tkGkz6d7KJmMwp9+THnJSkE72umazJ7bt1Z9vXj75YX7FA3Np7
a7fynLvxIfoKTG0L2jXYlVsVzT1h1cg7WupphFT3SSK6QLyEB2NQYr50anxJ4/zSwM1faoiv/6G8
ucZfpqpPrxSZMXN7VYE1uok8FyA3XCTBnEzA7k/meDct0aQz3H8HaofjctwfCCOBBDC7bRHNzNSq
mK/WpOr95aiewGuDJRA2LldwkZL647DIVVi1DwljhXM2Z7QDvOkPOTIkwoBpbLPtE9BT5GoWp7D8
JLGSq/Ugu8pJeececoaNRANBY0EQsQZMj8oNDDi+Cbxt/9BpkHbAKOdTACkH9VOoXkaxvY2PyUa1
TE13u8BrZO0PPFPALnJFj5qx2XgfktxT3UdYAYCe/5R68rOxOdbViE4se0L3H2Ku1wpQ+0v3am+j
mb9Zg1j5oIYiXXISNqQuQK5rpZv7PZmFyhqS+Eocnkox0/euVbgduffgaX5EffGb/zgHeY8/LIZu
NujLuETDkhRIQHxWHVzbLqS1NLz8GlLcKPpnNHfCJ6IkhVXTL7Y0QFck/1rGIMtB5W6ul1rpUX33
hu18/8ky2l0V5D6g3HF1h0B0zhTXeuYmhrB9B7hddhIjZObc1XyyKl+FvO4MNEdlJI5YxCw1Qa5n
qanj+cAx/By1MmANjllNPabDE6BncyrsXEFVQiAbNzWWqUR3Q/h1HeyNm94YDFFV92maGjDISxzn
gSvayRfOxGQDpz+Ju+BXMkYuz2aofM6LMHQj94CyQ1tO3+iEdaNys3pZHD6FHM5Xq+02AjJgvAac
AyRWvFzcr8JwpGUD/ZtWHzkwrz0F/wFFKuy01lYytt0ObAV6dotGBzED6NnRzHZlXuf1/Ahxodo+
Z9IQBIe/9dx0Ql/tjdnBy902ZFqXzzmMkIMKoUK1/UuL2qVIoGvbXfD8317NPKs2J6ncPoxJpGJ0
pA2vWukfhhDn+rQ6m8NXsxXBzT5sxAS1zz8a7t/uOp6m2oj03u/I/vs12n6wW/2ad3FpcsoG+waK
S/nKMnyRzeNrVdDigQxqORjQa9xhXL6ZJpRiK36lJSRqbsDbItMcglpxBrUuo4xetqaRZIowUbEf
XJwQYh9UI5zSfYQ6QAVmIsIvZFKM88EkaGotT3vQdBg4NEIqZyw6L/NZdr+SmWjQ+aBWKNo8Y8Ua
rEEkzeI9bQenBMfVAxU5PEvX1NWIChOZ4+YSdFsP+7yN2shiWuHAU23eYtZRMSbMQfZEHaFRc/FY
piLsIhbnyj51iBGL7WfRZNV9kMflwDim3Zmc7PRYnxGNeJ2GkPvHUdvM03kZ3FVOToZN5zgrfk9Z
DvgtZRmsVlGoQfu/UfEs+Vwe/alJCpclqNS5HmOTR6TD4wPTOC0VMVcRdYOjw8Xf6+Oj2FWHKTVS
0LjAYYpakSs2Nul5pPuE4lqDdsyW5k8gq99d42GXlpGOYbLVVQGxCCLH24zfLv06acKEJoesV4HT
WZ2KrYvYqdMe5S/c+47iFqpE8AOM2x6T9rnHDlamZp32X+l6Hbf2U92H2RCEaKrzjH0cz1IvteCv
VXoQPrYf2eQ/q4fWdMgWANVQb86P40gy9GZpjqmcTbM5rUATpNm2hJ6fUthHGx2B8nCDr+38X4aD
wsX4pjHQSNZIgc8rbf56l12gyzNFPnoX8AyHbE46bObMQ5I0CadOhi+feEpiEWE1A2UrAt1pH8o2
8paHO3StZaOd19rn5sOtovgBC43M0UNleh4k8OE8mBD9B36etrjcSxSxvGyOoVpvQprf94JKo4uH
WO0AoLByuFeAPyF4PdE+ehyya9BDWhU0EnzXlGmdWtnKgdbxI2aHTcru5IrdEynD4DSNllDH4bNu
9t08oI5yfJ+PCyerg/5R8ykwWw1vucImKPYCu6vFLu04z60kdN6Yq0SzjZOGf5ItrL1Yhc6hIZiO
2+CtejEEo2ABMey77Jhg62gLqN4cHNGColoTdAVmeT8D6LNxf0I3WkkpmmgEcdPDDBb4NSoR8iVR
4w3QgL+6uRVU0QdU+T0EMrCjgBdzplLTbB/qjn2j9DzhlWyMJtMSRpsXCog648on3AR9NeRFbrJr
db8bkHWeE0MP0GTtVR7DAdiOXONNYGUAgfGq8MI0+fJDJPZRTIAGKeXfHp4baJihWQNKJjMd1Hmc
YI2GFk4/sbiFtgBd3FIw0m3JqIQLtKdeRqinLLIzop2PfWLgyfjDoCQFNQKIge1OhGLRt8gWsg8I
VldoiuUyP9KxYQNN5Q1tMMCmvVZ55py02tVVQPpSI6N7VZ2zsPo6qEQnCU+4CK59hWG9rNMxvvIb
dNbY99JgRUdENayLpGUJ7Tu92M/1DgMCUaEsm4rX48++PatA3fwknNRW9/G0ydYbjGdXLSUOAFsE
YdLVZ49jphqhUlvZCCnszr1018O33/3ox+3VjdqdrNdCdXOZ4eGCcULdntlFqknG6Vg6CcZr2SSe
8fQQEfy8LRZt0P1RGoD2OG/1Qi9Fwnhpen4iN0tL+ziSiZdkG0PW6lrvSF1BYMxn/7n68vYZm5QC
hLKaMRC0Vv5OnWV5H40INpiTX5dGU/oSs0nxPdhJpSN8sd4L/G6cGLK349KHtGdF4IWD6vJmWmua
4Wv9YNjGKp48pSmvipeCK7NqPi2Lnoby1Gb+CAfNpGS5elWoMjD84uhdLrpQBnkHRp4RJOtfLrFl
Mc+NVNW9aM/RbnjOaeZmB6/bbl3hL9zt/SGLOCjEIVhNzy4bsCTWAIkUoiNSOcLPJbnEv170daac
w+dKo2pLNqggeLCM5msv5pNi8I2roWkRoi5ZpCPWW+sQ2hGuV3MLYreNbv7DQnz5woVwTU1BQZAx
eCA3rYJBchKc/KfmOm9/kku189SlyePhXbCYY6a6DoNpQKBB9hrvX4i7mZS5uCNGjELQRd0AUm5t
qbGnwOBdDWef9Xs6pYSuRj4qgVCp0i2gLfZyiiSnBrO22bm1MD/+94uJyBiY3iJtL4J78soc+M6S
EBu8lbZTBAPt0yCZAOTy+RXm6MRMdfTpBPpcvQAs/b+kDJG+Hwq9733+l22xKRfwFv4/tVZAXWbn
tdrVSb9CxpMN51GkqOD1B/XjH0HJTH+xKob0iPqWu4FySnHXI03MZMgrHmwEgTcsQ/DoHsYzpBr9
JsKvIa1cFG4javRx9Wbt6MYdb6zQZ6grqMiizWO6dMcT70SsiybkwmbXeQEcPvhDBuZdDS7MCmKW
9yYt8R6ZXZNa12S7d9/XExIJq3qPEB7JBIE3oqFnnoS3MXOa+r4kb15+3qtv11f/dwW6p6v9JLAk
sSMusQadOX4GfV9jsvX3u14fdrcfJxdt8JYboc9LVQLHBgs4MIkegLFVqmmIiNzM34x5HLQJ9Dmp
8WHXxS3Pc1h6/tVyskdQQvsoDGnuga5yJ8fQ76g17hWfPomGHSUDC6g3GYDQow84ZBaR5kfSvLM5
aAVbTX/CQEQQY8VKk3bDoehaaaFqsQuItGdTObx/9bXNJRlX2tT94wXIJMPFLz6IILvDd3HeiEJt
A2m6sBOjHgcinWc0rZkqGRU5ZJtk+EX7XYwCMp14BUPM/ivAAzFcMiISIZQiMsseFxKrnOXyNMCy
zKxnCWTQmCkJrXCrxPZhGEcX3aaPqpLoEz1sXdLFI0gC63UTRXeCc6TyftC5+OMBdtUczuvYfjwp
3clPIMdjM+NzLxIZwNcnv84dWZYzafTrHWiJx8shyXdd2cimQTSa/v8lgI49eIfEuTF0cIX1p7Hy
sEZB8UiodBSlffcZ6sz14gGOP05r8bQj+00TYODTjs/XURFUncPz4/zdReh8tzunF5cFnYOIkkj/
rfw0Duf/NQF6fvcgZX7fh5w4b1OgcBNCtNYUIn9Fw3OByBvE8RbomQwiQ7ysMlwXneIUAjH0cgM/
MT9SVLJJTEXW21Ztr0891V57YzZxUn+KMQf55LXhJmGZ0Ie89ZTFryCfDwJy2DXvQUfReph9YQhv
WapJK1xVrAb98SbK0XIJzcAVg0CpWSFxpiBL7aG3AvqKAZsocwYFLytq/9vjEQb/9DZwu3EiUkrA
UeOHVm8X5reIQiBgb25AlB01BRtfLjJk1cPc0fvMGUY+lD8aZUglbKLq4Bmy8gggm5vooqNtUSoJ
FFYsJy/y5eVVZNtNJrPIJFbNVLVc8GriRj404TRYxBihc7oX8iBtTcgKLKGLpwN3EYS5kYsdU6Hl
dBncu1ecBcEIm/GiLW/MkPfmPHLl7NVVRJJBU1ceqIcxUUwaXnneBm8TMCGLmPYrGYDH+HJC+v1Z
O8ryVun+afSlQ64RdnrtjR7F//zabJ8CQt2LIwwOAAKiyfwXyQUrd9JidnxxFFx251GzQ2Cf8ej1
GOiV2acP3fzG9pJbNdS2kyssUa3otGmQCrEO9idgEyhXs6Xv97OSA1nV2rbK3rGbVFd9K1Zq/PAq
+eBRN8wZQsKa7/TFQrsARCGPSRBYWCXj08Oz74FnMiZJvMhes2OWRWVCqe/KL2Guuly8My3/1fnF
gTIzeBSuQmu9fv4oAGCljgdIsmnLAaeGdGNduCjLMah3LPRc/exZVoUvXqFzzV+06HgWlE+1aDRd
qkJLaZiXhiAKx5U1UdO1+JPjL3eNHCAxMWMXhkbqoOEhIAJO6+50rKnLR3dygYbZsF0d5Ut1tpEj
v2Ha4mRHi90ysodCpm88t161t6SzOzQFfDZ3Y9HVzjgWTx/dZ6nBdXfCbDxYzzIM1lWnQcLMgbwF
tc1dhafxhjAL3UcvoMyqGttZXd7gyCpuKpMckF2rjJZh7wPcrHhhCi+gOBIDeheyl90/oRvGnYzt
i/RDaRB/CWhBCchqhBMghVkG1vVQ0QyHfjFU6plaxU6DqmNtslMiS5bhZt0T4mgIRkrBSh3vGi3o
TxbqM42Q7qXM+zP4ACr+8v8+JfDL5a/l6G2F5udW/yEPvy5Y++IfiEZmw0c6NqNmXucl0A+mPWqh
BrDiSJVMLdZVWAXWL4fBdmTzSvdMtbl4oxcYmoRy3QDDx7cz4LLkYMFYlcydz68VZKYuLmpBFZbq
0t06ZvnC5XuBpm5Qfwr/6CnAqLno3e4mqpZqKVCv4NmGX5x9E+VeSyH/pOimc9vRtn3Uhf1KugSR
+8e4hyBMfI7fWFUnrQ+nLKUND34LqvpcRjSm1P+wc9oajQgDirguDq+IQtbYVlOr7q0bbw905z8b
tiCJNDUyKY0ApKmexV958t6q18X9avohGVQ2touCdx+i+bz/uKrvVZHuWnkyA/MqKwP90FM0fsj4
0wQvqtgEIjzwP47RvXBD3sMMe15Ux3e8SPIgJLu4eWggjsTAAwtiEnDQ+8HdLDW2H3ZHZ3rigkyJ
EHx12C5yVzqkniLcQIql56rUxj0PT4l2lMDD2crpje8gV/fuANrxy0ugsT2tnGpO0aZ6UqYGAip0
Wgs3PtBCfn6lZYC36UJiFt0hqRNneZJevXGlFcy/Poz6E7EtFcRdEi2OLN68XT+MXfTqjKaFDfaN
bxuAvl3p5x15WKeIKe4w9/OCxJvenApXMDT/9q398t+VTEDUhjjfi5bohsDAFI4Ggr3jy4RAbfd+
RjtNjdsINF7UKv915IRFidwyim0ME5WQLvPz7ZFntXga/nobu1vJAbx/2xGlDVP8t2V1D8lzknJt
iPSCqF4uVHltybCDEPqcQ+eOWXid7sJTX04TIaLO2eXJY+vzUSxXvo6pTFakRRqmeREo2aulbWc/
BiZY44+9B76yBFjHCeHBfuR1zUgWgMtYNG9VVRJhWTQCmdU4ApdWUTteTjtpkuKI0q8MA2duOBK3
8BPCvQmY9OWGXAFuqPEfN2MQ8sj3r6XqwtUQXnkVMmhZK33oFAZsseHq+/bZxd2mPxxlh7Xl3p3O
5u2VgCpQax1dXO36E4fFrYY6w7+oAvFklylTtEC4W1TW6J8spTCu59aSD+rUfrNHOukslIK+F9NQ
dKZADbOMflVhG2Ym6jq6NiY8JbBFki4bSkMGCOEWGqm6avagG7FUyKB3teGkXcxIoMNNKC1h1+FL
Sxvo/AiV0sZqEbYV3PQIwV1JioQUAdcPkYR3LjqH2G01eOoy+MBeCRy42QpBm/JafO4P3FJ5Kxs8
9Ienfqm91j+t5Uk+YIJo6dhXwSS7Db2krfAMnMHXsByTxEZ23me5LaGvzu+qfRCBFZ/FeRlAcaDB
uewjoo1wbDjpVnOZ3cSQOKmZVfX+U4oth3ZMkmNDrp/SyJ9bzcdSCKL7rs2iKWJKYdJnbzhv3CK7
K0EoNjqXzPgZm4LA80CctlWpBQ0pGUgkNK5nWKfeU6Pln7g5byAYI/3Pmy6IJaRIntix9m3mlUmU
WqzbdoJGiHorIpzuPgx2lToDSPrX/v+QKcPt97yFwlAMwxhCE7Lp7Jh++x8XJ22RzbFQCYmfICW1
kcr0EpAnc/S0HCe3RpAzIod8pwhNH/kQFlQOdNAc19LTlBXSCfvHO/izlct7U1/Pdm+T33M8A5OW
bebFugsyoB6vRBNqltO6axkZU08QYWrUIZDp1dI+wz6uOnclNKLuQ823zj9hPNfWZNpNThTIwjyv
/1C839oZnQHWRZyH1pUpjq/S6Yy25otNpD+vNFGPETJXwvoVb2by0sjCRqVRo/yvWq8hMBx2+UpU
ms+hlvFuM1ZADBFgvdfZ8lQ2IXXOs+sH34/zREKFSgnIoBxEIcmlMuE7c8nLEENWsvoo8GS3evz2
Off+NJYYDOXANL5G0bJf7r0Q7xOlH1QNDyfbXv26TbD/SP1U6Hud8OrNNoHrUpPfWe3XsJma3COi
yWmAa/D7n75007XloZ9rAflnPwn7yMld2Jhi8PyWzrvGXTt4o9N+molqKGyZKTNC8f6IoOru9N3r
yrPA0B0hFVEIExyB47PMtX3ftPH3QOQ5nAZaU8PrFkoeg/dJep0BGwdx/niJkZ9HidxRcE6CLyES
cc9Q7LnVd671CruXObChrpmzdA2hXCRiCF5x/6/lpeNMDKjuSuTszsFkPjW+DSXcKtrIgSjiBFcd
6TcJaTWhQLyuCaH3tVNLXtJ1A6PBmUPDRgm7MvwECd3aWOfHhy/4vP03RwxBj83WXaZE/PVxt8lv
9NASy0hcoxd61Gb0Dy1Sq7Ir86DVk29s7jSs7du6EPQ8Qpuh5TWXtSzp6V7Cz809tbglZCovJsoF
099NjwzJtEXKRp1cyNtu4WJR7Cwt9QjyI+Yhl934ObUz8GpozLZtec1JJkC7JoTJ6L4tPwrsS2el
jPQBszVAKo1TI2PCrbGssnGD1zx5qgfishOrLCgsDcqQh55CvGBy8kApKlBSZqPxgCzwkaKJO5ts
fYwGKlesVpm3BL9WZD4Ree41IPM8Bf9iIWsUQL9qwN7wYbq+i49dGIHjd55gxe0Yw/ZEnze6sIws
ktjbMVwigtkY6ZnJFDa90o9Hn0W4CrEcOUEKOJdfDB7n7Epeobe5N1m6/KeFuq4/sJnqnlp9NSUn
NZqpsr1Ie8yAjtESVFx08dw3XOqHRevU5nuy62dN3JkWP1E9O97V+qlEFqYrjEyRrZDmlHhbgSFm
vj/+cElNOoEU2+o3I+X1sECuJrkMA6idLqUIi6ou5vYROolXVv021ZYASYNJErRefWPDmRbXgIs/
9DLOgxqycppaUBr/DrxvzO/sVpwKBqbb7pvl0+Usd2TYFfu+phFkPkwWg/Ben/k5DlUdNQ/HMuzS
G18ayIkX+ni3q3sYdFJHLLd1eM6ah92SHmNeM8AYIy24Xd/7yjy0+q/2JN0FtoT3iEvJACC4ScMQ
5Wvtjztoy62QUp72FmmfEo1+dqzP+PZ5enL5mNMaPjLbRZQFtHQOdS+UgaoPNBiyAyBbGpFGtBYE
tbr54wk6RAaB0wnPjJVbVK9dsYBEPMn1cO2/Khdk4f4cQgIOURSvPmFQ/2dqnLUKTCv7TQdqVR0s
W9RJiaw4IKHmlAIuXAz9a7sHAo4OAqQs64Wuild6l9oyH2XyZeZgGsGdoK5EatzsZEAL8tx/euDw
+gmCqjHFsYuFbIa/V9otJrAZHdu08qHncgKSOJBTGJxAdlECXOwNkUSIARr8JPehb8YlTIga+W26
IUUiUmsK3DbDjH8kZI0LAVomPBNC3cWI44I24COsTf8NZzVhqspUJ4+/nDkNvE+xCBnE6k1d9j+n
kx7fojjgvRSVM7wy62I1DaxF1vuALBjVqv+OrMPPabbAPkakOVcnzluUmilFD7RZDt5iMhuK5EIk
r5gZWjCyWTEDx+IGw891j5Ewj/5Z/EFwiRZtKVCODjtsuzHV/CfO85o1UDX0VAkwvrBu12a+0r4+
FRbIuQqLe2Xuqk6wpy2DaVWeWG5NXaKezfWGnNxjiRNzyTIQwaWu0VvSAU3PYMW25QBCiUe9pbVI
M3XUGmbrSqPEHUPPiB4+pqwxnHNai+LJRy/kDBdpEk+JSdgbrUO2NG+Q15wuQrb7ITZp6DkRAUnO
FIcDQayvhVUbzr8QFY4W/05Xz2EGvm+wvRY77Epeh9PiXhZ0Se+38NCkz2ch/xyMOT2D09XbQyFz
9I5txdAGKPw37/WpUvtMzMG+c1m6JItNNbE03Ut/fL85fpSfzx0N1F8AwyqnxMeG8CmCmSgWp+Nm
ZY2bDIncmq/mOdUQcyjnsnwx5PRrEhl+wqEXdb8brPc5jjOFAlIGOHb0DTS6AdYNynQF3XE4ETL1
QuqyVst7Yo7jyAKcUWTgtZWLTBmszZw+EkrFYwwA1TheGCPznRV7kAfZ+1f+QTUBUGQoHzewRii4
0sGytmj3SC0BR7kkxi6TYfru0EWI49DKWr5717zvAXV9oB8ypOBquCiP2k7cVl2tmFfkdyP5g7ch
BpF+wcBHd4ksoKLixrXLmkt9Fjr2eluydCxVQXgNlHSL0NwBH0HC8mhrSesnXD3NlZzBeBB61p2p
Y8dednbAoQopK5Q+bSJrGuguhoAayTHRqwzCZla9JjBHDYzb7WTUjr22Yvnygf6JDIZinyQnjtWz
+wE4kIhzcooOgi9lyTlyZeSC9md27mm4VmoOxldwcvmqlSejHp76HZViv/CAjij1/dFHvOrzrlHt
ZDmQw4ds1ikn8YjUJYt/+uTEe1wOubmnrGqGPHidrlHtfk+K/dGxMbjRtWQmVwDChAsWz2KYQkh6
lJ3DprJaqD6/u7IpBFPJpBp7HoZgm+ekTAhKMYqQL0zy3E8BKWgl/D6uclh4zJ8O4ptkWE/y+u+m
ysNgLhRc2XCvuENc7ixvUHYDFsuhN0l99DJ81MWMl4P8kc8wSqBjOO12QmPhYmuriasEVgx+PB25
CQA3XYQY7IuSelpc/YNw8txFld8YGeITH/4kiTX0rL967xx1q7lxCvzdyyEOadoX5zdjkE25kMGT
LYAFdRYuV3pkT1bYzOxV62+K+SilfteBDphPH/UB6fCmRaZmTq/RhK+DCS7EBqz/jPGyeZA/KkuC
dNbdbqcpUMOPfVlF+SF583VUfTE2Wvy8qG3Dk75fPDklRgv8Tazx+NgZLxM/GL8svZcOE7TQ7qBK
N2+zsmuYFuHINyff6WklHmD5us8oucbv3B+TFdJMb4IMEABdOJGJIg0+FF/kTSZmdjKSmEraXqHl
slwPKDq3GYCcO52rhX0Yig4zQkutJidQkTVlG53HKlOjHkDl/Xc2LsxPox8orUrLVzSTvQT23le8
WdqiMPIAbl9dmj9wW5mAUMAFvK85MMfs45S/ycE5sFYyC27ByYWqf5IDICWWsguA3hBTG9kaZ5ce
mIP981hDy5xF62PPk2GBeBVPdTUal99yGHlUz2q1d8U2wFAERMBK3lX2CAWgth8uaLtEgMYidznn
d4rShDGMmY+aq9iTjLhyDf7LMO6AlAlvGXR36NjqC7YJ2MG0Ca4A99aF9B85mppzjwru7cQs7NzJ
lnaHyEfhdhdYJpgNAoTw17+DzXpI6Asv5A6A308ySeX3lV1v3g48h47IOvENW7/MjI/P991nLigU
xCExXkTFyAazZLxAH/j2/K3wxM4E+rGPNgfSef7nQPBwgp6LGvPIt7qHuRjTPbAcKvuaidzHhoBG
shqGzaVCEKRt/eJIkpxeenybEP6ZDcpJgS+NzsX/7SYRAwHJEmjr26MaZwcS+QjBGcqZKb2fvzmU
ekO72PC5PbXtwccVwIIXtmnMhqbnrkEPrRIA6qxiT4zySIXkpqKir94MwA/cqLo88oLqQHs9rW2H
KX2J/2wGy1bNQI8WSCxMKQgBYIKlcusDkFwcnYonPLEzpk3W0LaK21I7CPwbtxMbDueh/TtO8PUP
C6+VzDG3akiP+gS+Wb54IZo6eHaZocp4oUsV34GZVNYbSCPlpGaBPntA+D775IdVfYZXzFm9MQdb
E1xMVukvJBdcQusfc/gw9u1CW2I/SY4k5QnCf/8bYw9PK08hQgtexR012WV+wHqyczPstekohWDX
R56tWMEGrjOKp1iYHcjzsyjMXmqkPl+7rXP2dYVslDMDGHbm3rueqGz5B0AE3wDknss8xyMSbtd0
bAjFSIr+eDnYVXdjSl56spRa3I5bSssatmRDDfrSX8osaER8fMS30PdU1OP7G/PIDRXCrFgJ4TUY
yULopW/6HdvdQsYqeQlVvKD71j8C7LD3CbByeZcbpDZZliITIpFHKKnLBrEeKAlmDx1k5p6MwYai
Etm4Z+39siaOgoAfNEelleWxpAPBaK/bH/8EAI7/hKwaMV7MA1qyl1BmpFRTCwFPGdI3+khigwcV
oS6adZgPCE8hpG2Yfjqn0IYAYWDnR5vS3D7HGdFvNVtYsmruaYf3lBPtBAVNJFbHTqqfrLGYpQim
2hUYbxpUbyiBUo6REoFNPsbvG4MtxpmdLBOxlg8ylDkx5lnjwF1JHoAq4Za4BdFqbFBscidEwB13
mFWkDVvYlibQNzDEUTmxdgScBJv2p4XhSOaYC3EG/QySfi2z2y248u2Z/jWKiQtElKYxfRa6mKT3
GPlyQD8PoMDin3E3AkBHY8RwvtT0jOz4JWTdRNG0G+XZBONV9tii6msUnTPLllcaH4acUUZFAPwq
IgxORQQIA/esqXbu/+Cye3SwyBFllkWYqcaAElGRJe54r8SmQl2pOPWopi3yde7SSVOgBZpatnLR
GTmhbYG4iYPbxW/lqgjKhGNsGq9IqaINHXpqwao4TEHwnyszAPFq+kc184xp7L5ddDeoV2mzJjku
K47kovtYafUGnYNB8eXNQyZxL/t3OxEMabOX+1Q9mSaJ2Edo15zxlfv9DDP/aaj64b2hd4ePP2TM
8lzJ1xE19E6XZix1PQtTQdLXa+PiRJwNw6fsqSkFQfY1HbTS4PMbK98VO7Gaw2Zz2a4r1tspqumk
0wEVZhUPT7ebhhP8ZXXbq/VHxGWm4UHWeWdU/01GRjQ/dafoHmhegFXPl0j1kZgUpWvbuqcMmKTz
G55ETgPAPn1ukcr9dMNr5LiBm+iDaENdqvzySHab3hYQyMZtCsf/taxXqDclV9vppF9+fvnpV+va
Ft82D1pUJF/AhRR4ZrsHy9uo2lU61oK/Ia0DZ+SmzxAHcCwWXdQrvCfSzN5fevu2zxjKG1O6XvSY
RDNwjGLuNIxBQPn4KHl00HHk0mNsF1RkRuzXuIbeho1WTzpeczlyN13Npgz87b3oBtDDsL09rljQ
wUnTl4iHe2aEkz7SfX36joHZgVyh009MA/t/EqSC9N83Ey0fZ/8TCUMVm4m3+DeBfBwSpvtf9m6P
WJwRNeogb/ritdbdbcsSbJ1/0cwhJ9xXhU7WF9YvBr0mqYZm2l9Tpd7ZecCeKg3RlJSvaxX8I+QX
ruOFS6N8SnR98h+ZgNdoU109Lt02KscchwBvpE/kRCRXBvIouAqPd1lUxQA+TxLluMkjxhSKORhu
nU6FbWPhVvctjNyfma/nsk69a1TfECNHCO195F0wRsAWYoHWy25gju+sFF3U9ckxfVuxgoHsboVZ
lxs7C6fuRNatbG3K2PUCiMbJEO37jiZyfYdJrvhPaa96TmTtPo0kyzRlKoF855QEnWMBmVtFWxq7
0Bzr6iAe6im9zWSToM9Q0ZK4dikQk3PNg39GWVbRH6DtPEPp6ES+L+UPn6ZTsifbCFFAF4tcfHV3
BEnX7/e+bpA2bPSc2HTt6qqccVlj5sDdMjLSFlbQPaOttnf/KCFZTeC2smECtpraziIwdSdx1VZJ
e5o3357RFGSsxkWg7vEfw0M6IYDrzoWII/3Qh2hYBVlSIhE1tgnC+Rge1q70PYjHf2ZCMd59Yd3L
BgitKttoq4eic/6XNeZJEYmHuBBH3dlivBlkdao344NHGlP57Ng7AW46g6IQy8wMv9LMghn+rL4c
aW1IqiUhM2FJzSWXqO4SpHyw9UlZgKlxLL0Q1/84ILL3YU/Wd7eADCKBtEutMkZLoNZ/EMq1CoTR
udhfe+USUj4YL7wm9juXrM1VDQBEaGZn3bE9sF7dl7Um8IgEwjepVdJ2W13OUnbPQb0Zn1Xt8Bl5
zJU1W1VHmLow3dmgzqPEALFeRatdgWPpEc1yISomZ7X11OuL8e6StRoWogiJgoSjX0l2ymciLbp9
6yYoYal42Fee44pBoP5PWbUW/lKIh4pRfiW0Pwf9FLWXSqaNEWWwtiyBdhjBkG/26y44MLm23AXL
98b9nIrK9TIOJWSgIo3cZQI5cGN7ipm0Kp7LO+WbrWoXnilgPN+HJ5TAaagu5VvXfop29XGeVJiu
zONg97nMlTg0J7yIqAUyxfAzq0QBncoD5ayuzTzlUuQrBDfbSZoTFmJlH8QWHS6svL4Ef7/h00Lw
xN9yqspG1tdPK6GiO9GEGPdsGkDYcAZMt4NBVBKB5qmQU9J+joLKgWPFZeZ/3PqCrFgc9bordKT0
CZ2+ctd/ghAnmDGAWFYmBDYzwcbu1zVJZKTjebxEluHK74JIrb7ifjKdNjEJdELiQ9jCk2Z1S65x
1noYmkNDoxCzAOtNG2g/D/m2mPJb5UwScZVZ/MepDsBKlNYMBD8Vj4Xu08bYTX63LSAEND3uInvo
KXGkp22sGv+pGFK0c4UkbY9IAtTlAnOxTIab+O2uh4k1Drt5IjZhAfS5LxRsWWX0+xaTJ3AdY0au
1by13lfbL1/XbMqcDOsGqHfyr2ptv+VPR7W8enijAwATBU/VUbTTioezn/iTJ1DeFZd8iwGbxsB7
TKYpkaOgz7mhaT1UVXZ1G05gzxe+euaePYnuyjWHGYbiHpvFk5qh2PcMfVPOT5JTXV6SGItVBzAP
9mGKkHdMX+nWu9dyEviDZ01Pe7f5znUU2LWjIBxfYVJ9f8Z87pV7JUMaLKXfJjk6RPgUp5omKxXi
BeKfxkw2/AW+P5AsKHAdIvOW/6OX7A+V1kRUeCGWrOeGO4YsMFwZQz21kft4xOZwPtqHl5xBm721
Dfc9pFRF8WAGuR6PPB4dAOyrxK/RgMJOH8mYzm3brY5HM4dNSTMgyCcAe7Z/9fmC19w19WxGWQYI
tFXhAR0y/0zRrrg7ylShg1mXgJKqeK/ldLRsdqNyX8uOlrfS/w4MhSLKDzs0YTHrYcykfnymdozo
9wPiKZWYUx7hahXsH7vHmnsqicmV8/NmAlTjQPxCUFRxwCHfPcpzqlF7KW12isgLNF795n8obn3M
3Hh97jtxmqWTBlG4oNjrHlXcu6qk86wViCkrSzXnSYMPhOz4AMd9MoknxMD2BsTJUmr/s7l+bA3o
zJvSQq0Lyx75f431JSzUL96Nj4iwL9y5NqM2abWF8q0YHZdbY6nLrUdSPpLtxWoNVE79A7kLj7W9
lv30NwJXxRDjbNvyfQf0LWcxu0E/At2P3xpTiAzkDLLO6dViuvGUFEnPBc+QJTbBWx639artl1pH
znYli2KzZ1AG30MdPGQ0eNOAK7zzGEbteBSi0H/dEtYun1VpZxA36eZp+mxhJR/odEKL5iYVK7/y
agMCEK8cm4/UF5yw8rtAtT9BwxH/imW5FeyI1SsVWAWGLQxHNVCs4+kJA/jud3ICKWx/QpodXALn
2V5NIF8u8yy+K2kQmAd72eDyQgpC14tF8fW3UO7aLGpLWydtblGILSGgggJbq6ggtRAlHIyG0+KV
WBMMIyozGyNtWwC2H8mKYYtr593o9dIRmOg7l5EQTd+k7DxCo6UrIt12gvDXrSfyMZERNzOBMWBi
jF9v+ZJExSIYn/kDh+UQEPEMlxTTzA4fhYBflwFV59wg2M7q1lrSji165kiwcK95oFu5R2H3CAZv
X3++3h9pgY2hBVcWvdqMtgVygig+Hf+c6jhy9hB5EbUzD+M6P5O4E6uArKJZr7yICrXo38spNGDa
/ehwLouScpveS3TLrfIaFZGr3bZLAZHWVes2oCltl0tDle0pIp4XoV0edGoXvl9gYtJnoAqkoEbz
a12/vMO8ncHWrrMs2o64H+6kJc4A6lFyBj8QMSy/486x4IScActmNZkMCj61RpzO7MbGdDI+i3rg
/5J6odDz4bnBuuGrapu8fMhRDl/OCRxHBQXlA5efL9hH2PgI4TC6QcOpvLZecYnm3gy54Sf/i0Ws
tJs/KP7zky8c8+ahWCWMB48vlZp9U3myEHgiu7S6qmjhS7Qg66KtYivoIsGDVRWynXR+jFSOjIz0
mDUlUax5pBmkfchPstSZGcwF+Hd6vm7AnYRrq9FJ8C6R+fH2zBuy3JaTI/5AX+LeUPV84pF4242j
87dHufaUdvHP3BsnyTC/+wWRdZ84hHqphZ3lsSvcmz3DOoIwZa/xVvsJwAekmxIhgp232jqd42iI
IrE21jtf/JV74T2koIbF7VG69cCHqyTtrrUh+FqlsZTC6NhmT473BgXCnLtFsrC5oJR0g8rTr6f9
Ryx3UpfhTpnRS2ziXAKJFXfgofbh1iwhjnMsx0L4bShuofatQIQ2B4h0lKNDAYGs3YOv5C9gMPZn
T5tCrnA1py7DtCkyE6R2Rlc8OAklvq/y8ATttTfdKh5zirBUAgu+4FSn0E9fZJWzaIDehFWpMjBG
qN2dbcNix8AIMXP+m2PtMn8RNvryOOvbMAlaBEnfge70brRkoSF1P2zNSmFlHwrYIPE0AQBSuoWq
I0l4PRY0+tmyVXlIFi+R9bLBvZj06tiBsUQlvfBWY0FnUlvmxiDbsmqR+/Jb9dyoeFN/VqgHVBKf
ohdn2lTZokw8w6vZNw38vhZB8D67r0SQADMBZ+uSiH9L48ivvSbY0TBBYiSzzC3px7zVeaKcZAor
ydlbwpkREY+yLd6ocSD/IsI8uN12RvL7Li3+ZC/K4LaqdW0pxxQKqlspmcIy89vMTqqR9RioBpDM
nkq6WkwhBhKIIS4SzMqybIVnUBBI7HAqRiaMcEnqho4ndPYmLbdYUfc4INYCF3rhV+G4dPDUdXeB
8rZRrkP1kZQdjiaLAMA4T7xYK3U6oJhuAQw1gj6dxGOy+2AOO9NTJYCEkUu3y16IgTQcShbaVJnA
EHC+7eMUw7c0XmWcI+PHIF1vwn05oi1HiRno6Xc/xdTYmwirRcxn1KXd6m1k9ZXNo9HEgLOWf09n
p5ZXeHij2YlmkXUAPR5IPiYBY7OqX3UuiaUuzqqmZh0562FNQHJaAQhVJqlVv7LMUkzkp0YJ6Nr9
/CUtHptWGaG9EDV9IF2esLL8xgjNZANLANcONf0CCnJRAiqDmcjzbZ0nCZzKx2sIWPMNb7o7ZYt5
0QI3CWSySiQSwCDTprU5orzz8swOlcfE73rrj5pBvzfjQMiLK3A1YT8FmF3OYCV8gGYk9BJmM/T4
WZ5TBhEDxI6W2bL9LDqgVL5cQbt744971ZrrcqAT8Z4UGmSkVBdtFVG3+m1YBmRmt7jtXa2JBNq4
bt5EQuMrkTpnUMr1kd/GeHdKXWlDR+uC8z7e+NEH3QHyWrIGr8F7BrLjcVgpz+Wdb9aNk48IhUzl
GQIweYKlwie1R99pYGjYfdLe8RjLSRAecFQj2SVZdZ8JPrPoxRyF1CbMny+Nc0qrNo/JCMsxpYbY
n/P2+t2Y/lQp5tCUuvxtLgppx2uDxXrLnjohbvNUZWPILAzK3OOHSyFsd5gAT9NRhxfuBrToOErk
XDxQmtW145/7UN0FhxCeVxVzLvyM8ym3i97wQ5jPoy6H1akdSiUlLMeumcBv90sCXK+o062Cy4eO
X0G6Xxj1sdoPtwKePqW8xVC1iWSVaLxf0S6BV5CO570OXTl1dFlfE8E26lg0jtrlHcXZkbSn1dDn
XlHEESWdKMlzKhixz4O4O5GX/yWVkpjSGdSP9IbOpKOyTIkMwwBi1fAOzcYZ48o70TyCie+oSND3
hTIFYeXJvToxanHRYp8R6V+U4PfT68NZv8a0m/CLOD6ImnPSqArwBy+4TBbpr37jTboSoc0IKOFL
wBzH94bdFb8ODirgWvnQ8L9l5W5BreV2KADetvVQP3tKtEtQmPWxloNKMlWgRT5l+YB/2vOPZ7Cp
n2ldj1uG5mkzeofbRAu+TRmsTQVI+MVXTJWgB6hLs30EhF2KrrgSZx0lcfZIv99VLz+qhotQwPnd
1xoPMXRv9kozTUOISYpChz3ulKOMnxRBj6ENXwQ1GxBC2p06bCkciDSHBeJ7e4L+kQtljdccF0dz
7MiAJwwQAasIJTrZBKWs04CdsPaUt01RLmoSE5jKz1gwY04k+6ANrivrt3LAX/bAqp8OxvGhYmqa
Vl1Uwekci+hM/Cue2yipryd8FEHTjhoLkXY1k5I9ozMAbpkJplgujrytkGLQYbON/SDq+jRoXagF
pvi+B90DLow26TZlC4euqcDUoySIfBHPs4cWhX77gXQ4vTyzAFxlGktvpkqSwOwmmD/XBaSQ0rcp
FDVTS5fjlm0TfWQgBQligywAToW7yc1ER7AZ0rHhN8eWeXDu1vEP+k/7PQgNOJOVnDg4YCz8BEo8
pBJRWayiHpnqWczmN/6C/FGYB7oLUCV46Hs3y6t9/h1Y8HAV+EeWqNZPxrDRVYn5O9tOGNmU3Ib5
W7s1mJdESjvs5cnbzVbZ9HPZk+IzZ3iq1KIbydkmMgZp9aKQZ8d+xx7X/fjnI6ehmC8RHNzeGHjV
Mj9mOgCat5UYkXyWPIHMsMn831DxSQynjLw5uM10rAEAQhpvqxsq4MA+1To8yU1zFsUiOKcHi3jB
mSL6LZvdGQlLciHu4rybQm8QE6FokKyQ+G8RgPeWVJEp0iogZxRNOWXniC8C3rSIByTKsDQ1pGiY
R07t9C+Bpa1ykKR/YCE7FovOBof9GSWzGloIIBe4XDS5tXqVEG1rFn36BpKIjsHPKGe8VIghhUP+
t5YIKsH+ISeBZLBfMoDZnDKCkREHqeyl3ajWvGY0jI8RQUTHblGoDUE26YcoZOcr78ADUCCWlxT9
OKivkWgJEm3sEilJxoF/Ten0s1YOoHBQchjP+8SHECOJZXbnWfgL1PB9iJTV/tSmERZ/RqopW39S
/otyygkfu2bPzRfzQfwtgah6vp4y3C1Ykm/fdCmnuTRw3/HW+7FoxDLI6BLr/C+qoksHa0QFd+Z5
oyutsHrRsd+iDY2sbq15gpvn1vqh1qJvZ9oJP+gQqZMM06eTz0xqysdbyaLAMcvoUTLobgO22MZN
onShcKAzIwAqRhh7meNbmaK0rHflgrjgeKedUnGdTyBTzExOy/jh7vEFet74SRE5rdu5FXMc3BF6
q1Ko/nDBJUkzdetKK9MdXgLqMsoYzewCSezMUludfWjzGGYbfnykuHaZn72nFN2TXSGadqdof5rj
tGTy3JrOIOTKEEfpOI6CLuT+zDCXc/sNnL/En6zz8Le/BUlZXZ0lLebyLdhmoNGlLAFGGkXSqa9n
0MeMo5wjY1vLRIhtUc/EUHFVloVTtTScvcabt/7DTupOuTUImSdF30dDpEsNkU5kIMwlHv41iRMd
+d9xEOnYvyqZApIYFmXzknnjAkmomSGG/Zewoyp2RGmEsNdNLLKGm4Eo5VMQkyGuENiTAA3ascNv
dHo377SNWkZHgK7ukZg6iBoMHnhyPn2Yh4/fTs6l5YuylTgdHmw1f11PN5B0e8x+jbQtm7ks9Y2x
nACgu3kFwfD9lGn8SK1TVNh12g0BMCpkEv5/7R7JYSVBoetdZNH8bsspCJbXz89U7HfdLbLwhxAx
Q0yOo0oYeckpEq5vrZ9y/efQbiHj/1+MpTRdwB8KQegOQA0uUI+eQRTPv6tkNhSwuZleU+l0oTwC
lf5TL5TS5j7N2Wa/W7GXJ2JZPJGq60YuNkjla2vMhzHHNrjZpqywUu5BIVi0cYih17TvZIc8UifY
gQqGYjKNYnJ5X7JKRqa8L3nSariiUWb2AS+lZ34sFMbQoei9g3XYn6pBBUbg86fI8FIO/ZgxhnCZ
fhX2k3QR2W0kUE/dN8rcuYdhhipCqkH4CbxcfmlQYhPRIsw9SdiAYxGd1g090y9aN4oRb8on5oZG
Vzc0qb2so9uL6PjohbBukex1cyd64ZMxM5PbGG7g2jj1zeGwuResCrbkZYFXOpH6LRQ/jhj1yfJ5
5kqVYtQwbBL90j+Qsqsa4CXMlBlwLHSAFY1fG1QbFqMy3gOSEoSUI1vBLlNCK2S1CcKL1mIjkg93
ykyM/XYygz9inyy88atBFdefYB83w2GkfytSty+2pYYNaCMXJkxLRNGbHOjy15QTGzuJQmIVZkt4
HNOTHiEgGfHyroeWv3+j9l46fyLMBHj7GN+Pln9ltz8u+yMU33TY4lQO6MUixEzgG83s+6WzZH4u
kNfkAW9mZJMYvceOgXysaTYkg8nAiXWlwV17goURTKwkfwdf/O7qnktbZJQ6FRr/G0+EwrCpBi7x
OmK6xCoY55ObzMeP14n+15ZsJ/NCRN8+cYYYF3wSsyCYbLk7gxhCPzPcwBqz3mh2o7yOL+9Q3QpT
COHoVk+NSpMwqiILeG4cKcHOoyfTNP6k1gApLtCiirVXBoOE9gk27AM7js0XYqr1fztKlgWvN3oY
c2rcM1XTpNXoSNbcX9j5+Q+Y6mJNUNyNXgHYCuKpq1DC0szDr2HnEziwasRMPgotniKW51wE0ysA
B3MtAsHetZTUtUQTv3yEf0b29RItyVU3J/U3Z2ph7HCjqRXk1kJ26An8Vd0SKgw8HPIVuV4K/NOY
6ZdhgwPsQYaiD9+fw291ccjUqsirLNPb0X7/pVjuWqagOA53IC4gC9pdCVw83+gnG+zeB0Frszxg
hwQdteUX5/3MS2l/vODJ9dIxMEWQTopeDyexPzXVbEspBwF5u+WC5esS86o8hVNpIwHCHoJFp/Ku
E5MDZFmwzYWYwkJatLoPFsefbY59YQ3Swd0C+Nifzt9eIHCwyisM8CTEVCHkA1kNnyyrt0UBykkJ
HJ1XOHvaUHQHIo3MyA4q1Qee47PH17zVUxbCA8NiY5hHRfFYFpgKNy2QfIXW5TooFpRplRny/C70
kA6Zogc94gqg4cqCZc3Fge9eC/YndWbNKmDatNw6qjx6tR/qav/BtUoqBqmP9ovMwLlcifHtqglr
XCtIBYnwBWk33OFgSJyrDVXfzptWj52i5knaelUdgIIHzmluVLcZszXiaJ0p7qwvnvjb1bDZw2q6
/anpBSYokV+/T/smwG8nt37PQmbCN9yRGe/HKOjXukm6lipfo8s1F36O6fMTyAM1K5j1kw+RYGjf
Qmza1/k2PGwBH9LdR7r0ADjG9juGpLvYwFdWyAbJl+pIxb0fzeuAeF2Ys4mydCmM53mpRZbxhQXI
cnxdr3RYn3aAQh1SsuydUvog8LXA3gQLuWZFZCG4ZA9XvS0z+lkZKFtq2fCoXhZZWe13cew7VHaI
89GwnsuYtecMG4AoK8ksqj3bfZDm2h3IKxTNWKgjRwjWPEowIYoMYzhsX1iT9KmfGokzGxnQEL4U
LAg07677mhtNCyJbXl2Xg4iwML18y/J86KTr10bqtfV12KnYaLjA6TPiGYVSs8e+Ec4FZaJdSpDx
TlKir7PYywN7WMFdohLyZigyeIhmFQNElG7Toj7fDTERIxQCra6ZVeFZ694Z07Sk1ZseJ6TQo4RO
c+rcvNcNwHM+V5P9yxCBppb027JXhhLk4hK83GhgRvWzNFTVtlOMR7vLUphwQOux4lv8/e3QgkGy
R1N/viyvwx64tgYasHJ+i6I4wgE8n710DdQjY1kdOLhibteM7RGfNJNgkTCNAsKgrtftUY1Qllym
JpEffwuw7geThT3nxAryoa0NY0vZBPAJQ7QWg5I/Pui8e67tg3uE39Gi67Ik8/Lk2PrdpL256Jyo
PrGhPMDXPTsNDpidhD41BOKE2XXpbBQW01X1GWhafpSZNlS9Xit16Fw31FDlFMOFZPJL1BRW2e1y
NcdDBijmHFhe6ROJV927vF7itQPIaVk+7yoJPoqAsYBWd7zdJRTrsyvrig54awxOYVUW1GSMtqPz
ZA3bsTxlDY0Ak9eRbhub+n+PlsrKl51a8pWFGfzw/8erGxeT1m6gprXvKvvJdap93NGXCDW8bYj0
hmEQcUtQKlJ+yco8v5Db7SnIVjqHM50qMv3k1gCaPZZ3YbU1LArmUFX0rQ8BsUx2sq7tIBvLyzSb
1YxSWoZeZzySehARH2T2hUHFaq2/woKurmKZBLkr07lmtVIPmrzNTjyRsHs+3NzHlCY2IE4Dv7wj
eJKw/lOnA9vj8MF2fn0b9CrxAI0C7Abbuxxt5/L4vBXA0akDoav8XTQF2gzOnBLgL2jdBBMhZugQ
mtabjoieQVTUznkdY2gp1R911iQ6EFhsh1jWvpR3YRe7VqUanFxUUsASj+n1+IbyOvxB/DwOuh8r
84LUkRp7yn959y9l3HFIepWUs4W1pcNTPenN++YpBcq5QNUnKrWM2LndOB34JcsvbD8pjhu79g+k
320uZ/accuNAc2xfYlhFWVc3wsVcgHrb/wYlAY5ITIbpEQ34wt92PCn8Cul8bAxgHmUrWnWieMci
PxPahFs2ur9RC9hc/5zAGzczAcip6xosOOWcc1xbX9B/DxiIidiivR1MT6S82Ao/yB5COX9es1ic
CKGx9eJI8wt4XPg6mlKXTYXfffZ07M+OnndYEZX8nXCqqxilp4Ymi1bqrE0Zsol5M6+KAP05MBUY
inZttUB/55cqeMru0GsH8CPzIWxFEsUG1KojThJ8p8a2sH/E7FjAienWc2CGrYBTIigOgxYgeKoz
NgnSsaOGXhpdzDOfkDVwVrpm6IaT5uMuVi8/c0HmBbP4PKKeOJf/+6lvBfC4mimpEFWpAHOlGVst
ZHe7KlDUeF7c7NwsdnM2YGZGe9jmKHJmEdSOpgX9mUOgNaS8oUyL2poNTepn7EX4vOXI0jvUBd37
uxF8MBETui/BlwZ6MXxElC5DeYOo9CUnbZOCH3YmxvxMrmaQix0DrUKkcAT/pctuV/zM8NGUfrNu
hPM1QzYsDR0grY4DPoniFL9SivJSECEd1q+dysMDJTRddm8hykXLrGmmSFqXIy1vmohQexoT+/Mm
5Uj8CY0lumgUq7GoSULN8g01/x0QArE6RSvi6Nhe4deWhI9VxfdGlbeFPpdSz0fr+WYZnlUasvP3
JGd9T2iLvettyjhuSoLu7dlo87yUVG8B2DOZc2FUruUbiW1f26bdJeryVn7Nh4DOlBrUVw9LehjB
hIac80Sfmbg/po6bUAHZNZp7moP2mc7AMDpo8sv1/oEDwlE2lSyTLmSxOL06Jz6+eZebnFffBo7R
1rLtJRwu8xWkl1R1N6Wm4rsUk1mUUpv5LI46MBiujjnI3R3mffxQYzKzDC4AxCz2OLyaGn3C4BCK
++keYVWkBxjba7hNyE1N+akWeuDHvplyzV64y02ueBnSTmidGnmvRT3xKtV6QnrQxPUZuDkful0z
qKBLP5tbaAv6LB+0SQSk20EotPTLqz/bY8jz9yfPgN0lAUCFKrgV+T9byZu5Pdg34Y3CDWl0jSic
Ph8S4Tsj/A4FK14Qq6IPa0rMJjFCtx0u/uTwGpIX9YqZtVFfctAr8Vidyix3aCqve/nrWSmwZlO+
LsXWs5exik5lqNbvyQ8kZj6lORkwrKV81CrD/WauySm0pcBWKTmEjOE2GHEcD/F+igHV8qsHu0BR
PxzsDibFB3D60je1X9q0qAB5S/eKlvwas7pbVwBTtuNBNIB5EBng6cmWKPGUFWEF8XMjAs59xfJH
uxL3FmL/lzl459NC4rDCEPSWhzpvrGivM2VqsqValDrUATq+CHZJREW6TWs1r4hKH0UIsYo7KC3X
gsY52nT9TLShhtZbuvN0fCUPnTRtMPFTcIMqfdOkdSlzhFm92VzBGS+LrClkDlY57S8NvSz8LAph
zbkdwlveIlBhHhdOWj3FIiiyVs06lzLwNMUxhCVkDwhbD8NA0Osn9RCxBPgLp0/HoopoewUIFHCR
2HgxevIKm+hSzHlryfCpQ1ruxddIGSdrpk3zPkSSibiMTyN8cBxIIpzdnXR24e0pCSNlu7QtrRWZ
qMwGToL63MZhPx2ZPg819F8uhr4j7ngWwY/M2e86QaoCeAkxjwH8G+PBHZTvLer4DhK5gfwZc8/v
rSCGXYPESQk00C8EuJ2UvfSpNMCuiDTi/NdCx6K1w8i1GpzrzQ+AhTVarHvwHX80F+n+/F/+oaAr
Ovp4ljEHU8n+mrRb3OdZHy3JGzjEYZjAuzmI8+yPX4jZYxmPmcO54FswSeZiYNWd6QFrD7RarLZh
MoRRpJlYWkG1YVVLYgGAk/a4S+MUcC/jlg13WLkLA95QCi7D5fI7oxgHm2Ouw6ucJi7wsKIEoU8w
FYutZloMikLimv4RHj0AaoYBV/lOUU22RRdF//ix90loFjvimUb6qb2Jz0Zu0ubEOmPP0zBgAfFB
rxlHyS5I1lV+n4Ch7ODfX+yhAiZ6CSn3m+B3x2XrQP08yKnBHi2K6UIFhn09cqbhLK2mtwzQg2YS
3e6CxZnYuU7jV1NjHYx9CMLNfJ5nB4eZ0/b4NwWj26t5RxjLuIHcGHBegTsh73CrrvjNnzkRvF3H
kysR/0aBvXN0osjqO8j1Qs2heTc8+uerEtUt6SBaJMR2v2aSRrwe94d2E9SjTEELgEpOD8DLq2Xg
IJycbGQNgEZ8ryqwb91JAwoRIKfj7kzKP3vQGpgCyalxZGSjA/1bvjryBBcOOZskWKV4AlXyJ6R5
z4yApi8qdZEzWnZbX+Za1h9a87FrGeXfQFzXwVeoORXEVelSsTmkjiA2D/w5IfoFJjhyMdEZzZgn
VNynoXJnqnjlp54VaLDzmuVxT2/MIB/jCl8NKPzt+CRTV1Kqlu6udCKRsHyQ4JbOzbx6hz/Jrdtv
bfBaVAZHU4pNyIwwVQ136JClnIJfqaZM71iYJmuiKWnAGRgjG6E6JQTNvanDz0vqP1xD5Lji6Czl
dFsiYr31OaJkYKjg0KXyAsK1dFSeikkyKeXioIF26fJ3NiiRgS1TXKZdbXk1Kg07dA7PE2bcSZb5
mcsqKwy7/NpJORXbg75qDli0FOT/OtkB5lnrR+reGNCHjRIkL8InrBJiIfpQXL1Vvw+LoMCRhkrp
KyabUDj2XcSAc7KSLRkesIoO+WjDf8wiCZN4VW1FgzVJfSK199iyd9Xkp3ypZkTHMq4OOW+dSLN9
P0YJ1Pkx+3s+bq/f6C8h9ALlJSUxSRSKO9plvHdoPrV4y9wtM2W62Y+7eFZS3xFtbN1w9tQRbChf
WZo80ORUJrvRRG+G+fl4/cpoIOyCs74Kf8TznfIFtToWNtP/Xo6QCR6o9uex/tRKd70o+QKf44uU
EEUdFM95xJCixrM+0DYBfEfsqgBz/9cikWnpqkgn+u4FXVxaIAZRfXiMDGcRFHvZe9S5AWGbok/w
hVzZShUHNe5fKRmk/HDqw+j9ylJLbgqIOGAw1/ai1GRSi67OjnvSkSlVAP6hUwdtyUsG4WHmVLpP
WzzeZ54FELhm2U9nSQZ1DgNSnqtA0HHF7PXqggUPTEWryNwrO29yjCuiWZT+mtBgtszsqI+i1GFG
1R5mF8jLh8uZEHGgKA6p8kwfMGx4PPnu1GRJlQ9/+2pmMCKlGr1tgSAYanoEOP+Dzpt54Rgj4CsP
6wcEPm7WVe/gmPalxDTSEAoH8bJOKo5DGNTP/vFuxWCgjjLkLtZx1CDWm/uP7qa9vFGr3/YYRFXd
16K3pU0m+XKjcKhpB5wO+IeyaQuRbdHxpgxkQSIzGT1BbbEDCARKnIrI3LJCQb6N7bUNtdVpodvE
oVvoOv/icZWDJW1L1ENSX/rplJMq8gGVue//oqAp/XBTNI9Xeb3PkShqSSLu3oQy4rOrlwpuzBC2
xA3Fj3MAKvRYunOaWnwcSSkYbHUAuUsN53b2O3yjT+hVPFe6sbGl2qKC6btQGH2UaJAlKBxrAvnl
Bougwq1Xl9jOHrycb7OJA/GOHPYkhYWAzc4aEDetYIowe9Zdkz729B5zUA34wP8UdYqWELuO7TCd
kb9nxipVa15+2lckV+6mg3IV3+1KQ5KlSEyMcdTy9CQphYHBm/NcBPvuM7If7+7m2nF2bGqj3VEm
tIc/g1fElzfvDAvFOm/YI/5L/8yKvXboUhkpEXwoRE9F/C0hjmGGOrGr84gYzYYdKhU18Nek+nuQ
wlwRKAcdpDzXdvzCGcJNhbZAB08NG9mDU1vtqOBE0j6zg6jiWZoBdXuIQgYcYM/f9CA872o9tVUN
OJjNnh2avK+CjrvWfzQYqV67+uFAgabhscMmxQ+I80Z3zRalU2tFTwKENNGdZr/w4kl9C6ZQBlvc
gAMn/ViQv/kzxIH4ylcRFu1CCtf145+4phsVbjelsxDg0MOt3sqfsyBpPSOB1nMrzMQo/LQd0Wkq
9rhTKsS4ijwXuDJNbS15xTuip/SO6t3JcT9V3N1wiYItX6wmQxYKxo12ExzlQiY+s4/8FGcCAry4
XBvml6WjS/TndwUbE30jK4R+Zck0DI0YQYHtzPWHhNvfw+SXC4ogQMx1qlQxicfcksgisHmkr0M5
+tyP+1pfnDM8opjVlvQa08DbPqOVP6Fs28TubyYEtbsNozbB5uj7CXtWxltGl08l81r3h4cKYoVU
lTr5tjnPcg2nW8gyk0m3K5CNGf6fYFIMZ+cYClskg0ND9mRvVHpQ1XhcoZHQyuWwYcXXavppO19v
zyH+WB0l0DQZGx9RWryVvIT420JlCLEw7Bds/6gK9ovciZjbA0UaWuO282y279Ca7NSHWIsTqpJB
ApCtlWDIRuTEbsp+9InsuTXOY4Y+uqNGxejW/UcpWMOTCVzSIOiHQWFoMjnhwSBOJDH8kC5UKAnA
lLp2f/VKT56+fN9NQ2Gnzdyu57Z7Wfw8HkhK9/NdeLeS7FlsRlyofLYLGYHYHy5jMW9kVroke2Kk
eDaqPDSJwSgCq1RzMgFlejPYyAtLfq2mOdLD0pYAmYD1P45FrxWagQ3bUUI3ihZ4gT2Yo4ALyD2J
aNWj+XXxfjLaNXimUs7RLjIpcSxKekzyi+qyYwgtRmkdY4d6x27TLkisOOQ9BlXNZjdGW8rYof1E
kY3bX2HxIyNfiDWEukfl1OE2CFgZM/YwF+r7WpwpjI1i1uMQk8mbVomrcCBVlyqPWVwWR/ouerKu
sh5h0d6CWcMkFfVVOZ8fItMZ0L7kExB/4klrwk8X72E8MrMzWnWjSt8408bnOuVtTtxc0fJamX4j
ZiNtcQj1vd8eJe7Fo/dbQ4jTNj7wc5HtuiqSaPrDYmoXE5sEEh5NUIYdvHWmKeqi/Ud0uNfpzNkY
MvZ0JJzHrj0CqqUg2JyYp7SaiTa+M8vu0qhN8RsHwksthMlYolfYmLkZJclsa4889nvaUWmKHB2n
TxAJJmWc6H/FAH4kjoxOIFc3Y+bKsK8Ou9lF8MdvJl0WUwg8VgRbF32nhk22HQAQiCuaT+TJJMGm
e+GiNYQH0F3BjbHDXnLXBiboKPTcK1uhMFC2XI/tZn5VqlA4WO9t1phidHBLuPAjL6pT7zEHp9Ol
DDL2qwdcgX9O1bQH86G3oQ5eXl+tzxcQbV/jXZvFbs/lv2eb/ypso4lFzuPE7LnYCti7f77ZiDA8
a0+SlOgADS6ufNXeF/m3lOTMg51+nVDLm6uaGfTyJ3GsqRp5myPpl3NS6v6bDo41xYxnvo7bUCqM
CQnI1YhcbeWYSru5WWeFizEHv5dMkaIuKAjas4LpawP4jMjhtx8WxfKPaudX+AwODsWHiDZu/4fE
sJF65/K8dTrMOPDWmnLRNGoqvtnIqmMAzkiHpsPnZB/Q9/+ZIzRyjAfv8ftm2He5+34Ko+j6gv9n
phUW7EVtzsNv2e5iulVZwqhaxIwniPLhvWnrK81vpOLdO4q8gcHfIVZNu0iOZPSrIRCax0zQOr2l
0y80myUbGsK3/HZSNZAfEzTq2015s34UktKMiqs537A7w2Qr/uS6dCLYWE0XU8qsZvWZm9xVJozy
PPewUFy1BlPtUU83Go0GNNpH7Ks/+aEQOHCY/h4O/gZc7TA9TKgdgmgxb1An7GbN4dPLs2dPXba2
/wsq1U9GeOO3nXTQ3O5nBszY+QlLHdYR2+nLmKCj0kYSPR6ej54toQLwIm0G4WRgqnhJW77qpuMV
CtX+mW93MoS+iHmr4dDNMe6swYOrI+eJu9jdClPdDC0CbHzfcz4oX6+0oSZKF+CWVKFMITsZl0Pd
Fk1zkjwpe+tEApw1wp2bWCQKS3w2JHNsX7j80Smk94okHFuCxZ+xS7iw2Wsk/M9TesvcegudkUE7
uImvplwMh8xYvyvwQtsW45/4+ZP67I9vLkrPeb5U3EQ17g6Wzo9wjQzukT35GAjfa/9hvPcmuY07
9zmhSz/lg66mec9YZyYet7wafRxj9J1VVI6Fpe4gifk16eLoZfJDpZKTv31NushF3CmJi2WLwVIV
ALGJo4KBoRXpAA2M9fs9ibFjfqRElqWFXLi5soaL5GH0Tv+1xs+8mwKldAGIt+J8GHcDg0HhmgXd
+TBoMSN3H+S11TNdXgYHPyJXtJRsGO4ksy2AjC/VbV1RcDNzD0+JBsN/02Xx6EoAXO45PDODBFOb
+ndVYDEXi2ZNzYHyG1qU1H0Qt73rxiS+iSDT69IDHsOBg69WvZYGNc+Jmk4XtIBl9c7auLyWy7Q9
5Hrcve0AZdQmoLWQD1dRcVGT6vpgYptbgDZqTS/TD16TYW2p0VQugf8dF3i3lqxzSoQSg3WVSJDP
McuOhuFoIhjMGiTDRj5kEx5DPmKaTDnFmY+2Gd+qhE96G6do+fe4c1jyo5teOlw77t5kOWN3qtEY
qKquZQGljorOAXAya3hbavqjVSH9WWe7Z6/MszFFFWISabOZ6P/YKiAHmwi1Exs+tJq3adJh9ZVb
MTWj/smhcPm9X0htC71bXvaWYV2NXkPSQipZ1iyFDwKwzMnsK0oLPL3FyH+nZZAvti+FkNwxokib
8MoaXV2iM+P1ZThr0IdsW3nDR2/wMS1+Tk+AaUnx6X7UCuovjFFkXi+j/irI2dBTPelFPdiz3fVY
TeJGzYsKJzfdKZD5e5kgcU01xM4Yro+cA0+Hwhdd4hLCVQdK2p6nHVEBfydbtiCTuf4P3hSvZAQw
JUPgjIjqjDYuWKCjthHrNpRyYRNnqsxgGq5wkKlHj3N5V/Ph1nUdjWyj4ETiME8XakusVnzET4ey
s5KtsyVuFu90qpJJ9YQDH4FowL/2zJkTd3WMyOouGSXoLTbFn7yr/T81xOvKpSz4IrHAgRtIgZMP
XsEQh3NjB/l2HQaMz3LAx2inFJBOMlyDCVWSp0WybLgfObx7jTsMgyW6qs/ptwTAveyLqRahnWT8
nVkOEab7a6Cz+VbsiBLXXL+kibzoOP1DIVxT5GAqsQbdM57n4byhkuKxw8uznBN69YI5KZNqDWw0
g4rmRpc5mgji0F+Io7fjjk95pcxEoSi+ml2TIbdhEu9DyC/gvMa/qTAwIiZsAtmnNQr5RF4mZ9O4
Gw8UIaFAUgNWpjdreS1U1PfIinppPFGQO3Lk/mD7VbW+1zz2SezcBMslED84n+uVVmM5YFbV4X/W
cz7AinVwxzKKmqwGJSuJAFM88LfmTWtx+fCUF+Pet9Ajq2AmhddMxtUfCsuurGHpS4VLLTGU09Gc
qVY+QA36DLSvAIiPtaZ9kOFb7wy99tK9aJW+mDWyn9rBq8yYRREvhAFIISySJX6jJzM9iDIwfww4
d12bzlZ8Rzby1LQmhycPmJscfzMwN4cbx3LAPCSaw91fSKIrCBBQSJQVrmzjZykP+q8xut3dEy6K
KatWxcgmu67PMqS1Ubvoeishe/Fa3GxOBnzWZVtHdhhbWc0rmoDA1FutZ+yWfdLEfW/TJSnxs1NF
PshMDXnjB2jewwNpFT70fWHJywY19DSoln7aVElJ7jJroHSlnOwUkgKn9luKjekIk5iMmYkoVc9A
hCGzAmZCLGS5wh2vd/+/50o9zA/pPQsqGKchWLeUY+Kz4Eql9uw8lLAplwgnrOL4szodPw450uVx
dUaTw93pEanlioEN1z1J3BkPs0XK0fUih/DLvDRPee9d3KuegEQEl6T7tyqm4WQhYSEml/FXaAEX
F0JGx1H+Tc9FaEm5aQsZUQROa2r0tuhYXRvdxx9APSRgEEHQD6NkBunbe5w2jYyi+LNgdeal2MD1
ZM8S5Jjt5giV/m9NeRnBnNQeoS21QZ7rwZrnpkaAAKZ59rf3ezjc4eJzTf6xRcY+Uy0b+DFtI9iw
wbAt1bhfslHK3PESgj1W0RHfJ28nNNeBdtKxFSun2jwC3lruuS8XHVCVLcMFLyMwDK6JIbSTtVMz
fJMwOKn7Ib4y+sy+vF+u9nlCWrgSy+OZYxU7fmRYYmv+vVHOMsmyYJUffPsNkWWzme9cVheO28q6
sCtfBkBBULgxIxLznIss4hPZHY3wB+n6Cb5sf0xO7hnTNRMTHzQxYa5T5480sv0ylkNBD5PjrbwQ
zqbXPY9mgaDBqzwexs45NrsYLvcu26Inj+hMlBdazoruLXifHYVDmqp0opHU8R2AC744eHB1hv2V
oWVi5sTTZYx/oDbpbsylSUSccRj14sPLarE9Pz+8jmtfsJJomsAyNwZtCfB3rPgpel5dJtqgRLvt
tNzF9NqLlxFjoMpk6+1ZNglFh8ZJtqn1Q94D8faMivGcjHmG3h2pxAnCrgLFDfaIPfkjf9IEuePT
SSeFuXjlTojys7miTMboCHOcnHkrUaZlsaXdA/tYVQUCiNrAS+/cm/GBw2WF8aIhe2f7ZYTuuP3D
OT8VkuquvUePJ4BpdTeE71ODkkOL4AKmmaVuhStcUM26LAbTh0ipPKOQYUDf1FTrM20BChMGGSNt
R+v7FkdwmCnBjib+wYApopsUn3g72KeMBYG1y7wO5wWMGoUSettdnc278k3COBNRq8Pc7OgGArZX
Rs1s44VhoFU1oJxndXUY3zgBrN0YH3vLhgw0hugwrju77iRB74/5dH7GMC7Xc2ANzByt4D1F0Y68
7u8RrZWpIWjFYBesJUkEBI98efvZnlUv0ZAlnpbP+jGyysr78qtYxuQb9xA6V40tSgs+C4/ieMvm
F5wBuoRgIWenOf2mqddPZBxu4NDoNlI1/cY7c4/Orbund0LNZN6BZe2uL/VnQVLt8YnI71F74KLm
ytwV5SJlGBto1dYisu8F6oAIw+CfKd6B4WnN9h7PdlJvxYWB+l6Uq5eMWuhRq8/EvkzApMKlc4sM
+ziCCeLQru1OHweV0JR6JOaLOk9YbcCS6rBCqdtbxhjVj8c7s2bLx+8odW3Dm28emQSdYURiO7ci
Joav/QoewEOs30+fCfFzZocZdivC1a+D5YI14pBLcBqipbz6TIdl/bOM4zW3l8JYtVslo5VOf/7F
/SIG8bLEX796a8suA0aMDQLEqNi43CJA52BcVeN9rdZTY5fmRlsovWlX9S/z1BeEAk46eYW9cxdU
yYcbPKVsMBa3gdzc3TRGH3WyCXkRMOgi1mnY5caOZylH8e8qd3hdrmnMi8ML5A/Pth6df7mQbL/D
2hJlsNm+ZHHzgNPfTNxRnPPIOdAcvmyRfRFgftTVzAmQQsY4wIuMDJURK4DvXxbuQ7sYqP23krwV
nZt0mLcXZfs+ph03LSCS06ohxxJnHowBU4E+jgFHLhkN4k2vwYwBujY3PpwC5lKMtvHl5kF9HIPJ
gt41CbmyuyiEXLXKiFKOaCmV9gfQluGABkvLqyFIYmham0hyMjFvqw1VXk8RvyJxI/tj4AKn58Qh
0QZO3aZovFDxFPHxRqv8iWremd8JqW7Xp8wWoo8D+aMXDvb4MH9lhw5lHOIKNL2mxExMNpPEz217
PDFIQMEhk9Mh21D2uK/rI/oc7YCxN/RPy5C5d7iRnEuROoRGJjxlqQlkh+9IWl+jJbibf2SOyHMG
fPkCNp0WjGvB1CuJLe3bthtZo68ge7flQd7tl3yQL/KFgkJ7gol91QHVcOgNjK80OgHyy5gXQVCw
I4myuOrG+6J6rxwFGqO8uJcyrmR9V1PznUbFub21ysIElwwxrVgbrJn3DPDX8u9xmSHNUU5O8sGQ
tK+jHrRh0ZNCCrsfYWhtXeLLFY3xbIL4Yb89OAPyZiKDwgaPJPL/9RjSY5ajTNFzluIkcsN994ko
7amRcrN/SPtzzmzrZbGR4ksAAzegN/FqYEfSeLpEVOfE/zei78Yz/nijZU2lf1ivkO0riH+GZ9mD
6Dtu86X0jdEB8wKufIYxWfq4jo8b7L1kf1uOKJMRzJ6MC8CTeXH/8fqEW16SZpDUy9YAmP4C+N04
8xzSAEHAsNVz+6IQzRZlLqttg1UXsHEiezh1QvHO58RSsgclWw4FTJ6oVpGBpHcbXqT3BhuHNP/S
G1nBB/Jd1q4lLAlh65vtiGqbCeeOd1ryAGI/syaeUgMbKM1XzIFKPYX9Ak6lW0osk5KtvLid5CpE
2gcW4H01LJqvykfgStH92S/qwWtr/9LoW04xy3B6T1NI6LAqGWPVNnvvojmtrupIjuIhhH4p6F6U
YyQWR9ttrwaY0hZh4tJzNzb1q/67oeJ9BOYOvYs05X3L+b4GWDZObvV7h+V3VrTVYtnBZOAYH7hQ
Qd+1GY+2+TIXXvFwcs9GecKOHOeJd0Um3Pz0kU+f82v8QrfFo5iiBC7X/4djfUn9GlOsANP4bU8h
ewG/42I0uRbsucMQxTKhI2bk9QUwUVnHiHYM3xIs71P7PWYZnEsHUJpowbs6CZtk2nSgt4N8MiXz
63+Xr9PTktJ1m1YRT7d2u50WBcO2mr4l4pZrofpCbQotxEJCNa56ObZEMTqMgu7xAguBL4GUTbt8
MkYSfqbo9FOh5rEQbGHMcXyZbRnq/KFec5M8zcmDSziECkvp8SQWNgyAeG4Yh8VRu+njotu3PGNs
TnYZZbNCQVriaYWl664ZEpzugMrfwGXdlXctB60KPYVg9QJerImJcSBeZMfqOFY427A6znsax9fg
Nu+hV/llRwXKfHgzXzkrp7xIArDCPr6ufCGYR0Zf1FbR54CxGAmJtGvNnR+GSdmafeX+mQYLbu8e
0zj0y+BSBucdueQumJDCV65mi0ixRYiGqGEtRg1MolpU9qBGS3NrZA6+qzxXE4DupRmWaIN4lNTn
t6UmlbB0R5efAA6y5fbOetkUN/kQcyRXURj6ijH12Vn471g9SNnq25Qp2IgAHmVnDjUoF7mn/gNd
mNcJZcQ8eU2YkFq4e9YXCaaKbwanXXfPuxllKgD/C5UP36EtalUH2RRcAmAtzGDwQzubDUTNedRS
aqs/JEqjNsW5mv9Kb+PJ8vN6V22kgfnlFlhnjYyj8X72p6Ub+Cd7brXaehQ096UWzRo+kf6tTPP3
LF4o7ildfHHaT6wq5fBrOtbKXLYRG4Se1gAPtIyk9t7Y4ZQ8LA+yBIR6+cNjvgMCYgp0nScZcDpf
T1sRpuJEPUrcDdabIRT+etSSVYvy0MhZxlZTQafhoKcI5D1XOsLsNsVzlXGO66GXcpPzvM2ktlMP
foDe42HaJnR3lxFslHow3xd7ld5v8Hn8cPFvLoBgczJ9Nt7O+MlLHAiF3af8NZj+SDJEjlJv3eO7
ORLKZLqC1IEFu1u9R9sRkfnkBBrsHzpOcpee4VxoWs8lI0xXO2H4wh7NBCROUrnCIBbkKdPhR7M0
yw/Vp5PeY2xVniFM9qW0qasPLtPwiigOTEczSDaSDZEipLg2dfBSOBfnobrbVuqMnOHRziOE+Yq+
z+rvV9lPecsy6xVvHG+CNQbu8L8VxlghpCDmD42ebEv0o0wo8pE3xDpVIsgfY9O48EbF/bYKy7lb
nb5Jpfgx+DKXIQl7XLLQSyxzvVvFwBEA3smvr9GWfaAZNZFw+Ea3TCKqNqxqRYoId5LK+g9Y/BhV
FS/vjPl8tbbXHdvNCFnDw2EKBN2r5VYDUPTzJvT1jRRU6VW3FtaV3cmmiYxnOdZv5AwVOzC6g/vY
oDuod3ciWnhQoq+L+Hn9QjFv0tF07rIuBSX/U4/npQK49iqYdUNHS58gRdkFZ4Zc6foKWmDsfcLi
7f95XnS1MWq7TYeV1AiMIssCRkSYDKYWxN1FF4HVypxXTGRC7zfyHwj9JXS4Jz5jHKwqBvhPg4yh
gvirhHPEwE3UZNTFmFknrUSaEdUy9jURAnO1Ore4MkdeM5+NTHS8nQFkCx2eUz1gjARPWjHTBZ5T
ExTki5gv4rPomZ2JjLn7tDDrcLiG5Gfa7pKPxhNSJSvFQkVxuOi9ncE2ylxB6o9koCfFmj2QN4HV
5lW3OWMIxEl8vp6nBy0bPzTJZIpVp7iDy60EZJqJ1S80nxO0nQVGwWzS2ElllSAru9/95hHQzop0
jcx0Yksw7LGNap0BntdBeqR2B1gXroC9sIrCbgbQ9dIgIDD+9oHibXe5ks3Qr6e1CiAIciTFR61a
9tg1pSOUbJZK2QYbt9Ryx289TqWYQECH7S6PYaB+zkxfx991MYu2vsueU5KI4+dXLRchXGG/lkzp
uuivZRtvZ3ry8d6SXepvQbUk8Vv8cs2SR7YpsGUTjAqZ1M+Ojbnq94ql6q3UdAtrxMjhPer5tJcT
lLJFVnPfa6o+pry0x9yilHiZZ7oJ0Qkjhcp/DAPE3SBjC8nUblsbyk2TH9WMuncd6ZKRKhYl2j3h
ibMDXN6MnAsC6tbzA3wVrifsXNpx8aOMkiqRG44spBfEH2WKXbztU8OeYkmdfCP1rgeTPHB7GC+1
ZVLoQf4z6BSApTaJ7hGcFf8LtHHjxB8xetiRVDIaLhNv76k8/dCt95upW85RnWKwcpNEgxTumFq0
NjQOuzRlcJ6uIJoYflwBhTlFCzc7H2eHtVcKzYCAMF0G4RMpK0AjB6wEHrwV3Q2JmKqxD91t3nvI
weR/Ar2Cp+nc4lAE8ZHXyPTg2PKInBR8wqFRHWkVSvZ6bI+j37QcOHS9o4a/B48ozgarSywHji2h
mrN4zQTHSmBaatrUfVwLvpsiDU2z6ClUaJubpxH5XMuxdsA4WpMXX1kQR19CcnZA4kzU8wbS1x9C
FLuq0yA0n1z8/lNIRUj2RO+lz1mi1pWSno043Kjfso6CBtgPFYiFDbTHtMTRao8q+ew13hFmWIW7
JVfbQfwsd3MUbScbUj1IaDND5NXkLDoSrCZZwdAfl1oX/fJNXLriZUTpllRibvSxudqsKQa7ZHgz
C78vuvk32TYeMdYEtjPboOzHgVhFExwoYHMg6dZ0wLoHv1orxHwK5JIDJ/uPu6fctJa8EIDIPo/c
M8jL8tlOSY6nNNOK1NgOKuxEsKL+3++1T/a0/yIwgkv79Cg4AnqoRM8PX6+h9H2W23mOGlNiRcOU
hXmSHrOk7/CGbc4k9McAzZ+HdaT0qgfVlBmp5xjQrCqv9+rAypO/Qu16zIJ/zXG7CUnI1MEMo+To
RGL8iiOSIlqS76UPmA4BuY0FaSopPAIrU1Xmpp022tCEUgWvhUoB56SFSEY0ZDRkaGyRFufipABZ
D5PxfxkTsSaBVsqeES7/Ovu64nUeflWScQotaqIvppHVp8rvF6+lqkRvhiFmBwRqUaxTNgx8Kqyo
X+5typBSl6KOK4TjLxVCYuVtRDSFS18Oa6xg8YsJoGuQpjDtM+z5mvHgKx+Ig4IX+XEXyvEJbgFS
Z1JpcWvaRFynpx4Ne5AGOolflC6cvYajkXhgC0KOVBAvIoykdVaq8DOcZS4LkxV7PM9GEbRo1f2T
oCUDDEdCs2GJBphLFX3qWHBPcWKnY0kWM0RPtIw+CAkN5fApiu0xVqF00XO7CkWsOKlrvqpYRPa1
LL3zV7fcX/Ixorg1AItl/mwDBUZIvpDWV0HEsNSqDT4myrx9mJwI3cDRnvVW4qxB/lH52opzOhsP
DZCGtc9hJWg29HoUMXdsjF0cS3SL3jLKw7vCDIJmSrQFVCuCwb0g8XpmgkZ4+nJqAyqoiT23Glyy
Otn0aWQoMTbHiq+BKFdvM9x6DoxEKPyNdSbs22vGoDuDtTiSJYAlUjyR+BchCBfJ3EffEAY6+IKY
jeInjrwViVHlKcp0XGSFDqcI7FUruPFfpvR3RnVcb6L01s0hbWYOQU2mIHSDJvxAYNC1Ump+7jY3
vV0bBzCdyjMldLdkIUgbSskQ5cQVu1YyylZGAsh0w89C1d2AtcnPHzzTSlMAedfH6Hubq6Wgi4Tp
VxnkDyRQCphmNjYGrWVLxqEo7fu7KUDs8SAypTjiUKKYNGL09IuIUgDak9sYb/Nra+k6RpdGK6eM
oXtoEl4Kf7zCJbIZsviXYnw0bcMJl4O3ypli7CH3mWknbR3M9t8sHeafXvgYxSbHWM9Qn2ILTpmi
1Y9dIb86j0+PRzieG/ZNoyeOkTilSHMTjsEi99y2oCyUollnjrL2G7YNa4jaOyWU0eSFoDw2/Z+X
aajvyOMse/F1+tCYLhD89N9X8hNUdJRVPv8ZHbqFmtPoSsL7GIihwRQOTnKb89yRvDsFe5hqJXW8
QgimRLt4aMN7DZ9FfKLNISmdm0F1E82uhkixGH73Kvcnosw0jgKg1fIW/VdQgIAlo+qA/qrTzMRR
SrQTpDk20EN3SU203JZDoNPIVDGIG/0OkN4rKFPOWmI7TGq4tXrX5Xttkj2zkRQaAzRWTwBUjrZA
KuaVCIWGokKQ5ME1p03bPuazcQmZHGVcDmRgL66QqCbv7Zro4WpCLBCrXSL0guWcu6j7nlyO9noG
cfknFyCYk2HwE+YpVTE9OYj5b4Ow4eaC6n4FlD1i6WcxP17YQlcjVrJJTOkOxQNMgZWeOeYzebyX
nREFvhS0ReWRWlYm1c9GhgxYNQmLrv3HQKFTMcMwStfZyX2Bc33Ayb//7ykpb2TrNWvKhnEH90Vp
vxiEm4xcqKBiUH51sC3PZ+yNvX50AfgGazjiD4iIZUIC6IeVtXzO7iBy3wu+B/BksNC9NWYUrjlK
MNMPCuj1V4rqVIHHqJzdP3e4J/RABHwYAcT3hIi1Md6j++ZwM+kbwSx6tYzjCiKc5p2sn7JUpDM3
YUdMYbGGOr3/H7XWHppYxLXUMvz3p6NirJIYsQ7a7B/GJVFhdjL76G7kgMXh9uZsOgJGLUnYcjpa
rtB3KrulAOGdHEVqDZN3664l7klZHTA3gEYVL4p+OM06Gnz8sg9eeQqQx+ik/s3P2EWm+AUChpv5
kIkbZ+bHl9v3HgE0bEF8BylSKruj3Fu/0Eavp6ODelBMufL2EyFCdQw689M4wo38bYPj9S8luTde
knkhuJuOfE21KTBwDILuCbJWBaJPuZ+i62U2WyvsecQ8rPVp0b+vPyNba9YXYVtSJyYoyzseEkRZ
DQA1oNgcILWPV1Qm6lXyHt/dtdawikyTWharZ9kcPmbETDP++J2rqpaMxkGgVxORNlvDL8E/xO5c
xRW0/goaPsA+cjDsjqzmFz0HGWpv1NlQd9jmqtMeStoLhl7Q27ub70Rl+i9tIuIWiolfjCIlqVaj
XMM1PoblL3qMcRrdYHVN17RlGHsM4vT5PQ8z2zO/k6qaWoc9PVxsuCqT3G6JVGcVSw5ocDVQs5Yn
OPoIH9o5WtXTArPfvSkgaSGLedUhf7ujxi3tyTlOwEKgE3cCNypgYHA2cWNHhVRXZzUwm4WMUzwv
f671jMvEl0JLGLnHUO+UL0zBfi6jm0l6YB0PqhaIaPoO049N9LIyIJ3k1YzxtMOOXeb5AZ8QB9mh
+aZ8D9L4i2J7s4PCHlHcf8va2S7knwODjB2mLpYGz5iAfoMdR0IaY17W9N9kYMg4OgbbgtH0vTuh
rg0NRbPPFZyGO8D4DXNTEZMCCfrzGabDfgCl6H9sYPpJlG/XvtTlekudtrOm8hozfctwGKEFThPo
H8UqCgpg5E4OMld6IaMRnIsTRilvc44QRaYAAlqVctYTLEMKSyBcPVm4U1II+ADinMMWwJg/C0VP
sxXnz83O68pNs/L6BQyErTVpGSyA0h/P8QOynul0dR9o4xk/cGTYZ1W9y8qf8I8+iACBpFf0W2cF
QjL4S8VxiBFISMvdxFetycquWxcHiobSlAByOX1bxTbVQcL9rHtHWMztkZSgCzbdDNTi4xd33vX5
l3C5uRjL6YuIew1qVAKxRTuQHYxHpBWItk9hT0KJz2bkOlTHIJZJaiAXX6RXSZgBc+eNpL6x9Yxx
aoNF3OpRvk55PtYGn0A81MG0Q1P8J2/iHDmCnMsm1Y2aHsjpNk3WKf1YBftsTjeoUME2OSuedsAj
sJnBxyBMZv/CEzbDt0J6virskcbH3J6FSzUf8sfKuCoOqe+mp61PIllEh0TpL4cJw+XtwN7laWHF
Y7EcH1StEYfpWJeM/a1avEXGpUl6KthTaDl3EBKrEQ4k3ZZsc+ggUm1mfOSYFlQdn3iyzdryRVzO
myedKblGmegMljgUDdNfFenZ+JGfB5wBRp5q2NPNaSFa+BQLhqFJM1YQIbBh+06d5gtDxjD0Qncq
MCPL65S/oNxRgPJpgSz/vNbzNr/xXtXCqxdOQPRwcjzu+lW/0OFfgzW6tFrr9AZEBxyYUXpP8aBO
g7GFxCA0zyqtQiuSNem03K4KjSxuaIKx/4fBlR5c8Mt3wasnsfehxxQlbwuIbdj8AFKf356g+NxR
bt5u/Bn8Mcj+UyLOCH91FoOzPUrqsIfSlnPAQF7kHoyA1bmkITUlFLAW26vIQVEF/o7Kuy7kXYGW
q0A7PJYkkXmtGO5UHOs5XMDw+Qxc7qWWkEGf/zGkawZvxLXkda7C4N517qMByBTnwtBUav+HKr9d
6FR8ZlVvigpO179MjvLsEdwA6PoGh7EO3YNoAcx9EpwUv7o3iRCWpUjoPObnwkkM1cWTWxga5gRb
tg+wVncYLAcit5EzORF2a2ofTftLZQnjpl7/L+M4StR9QYlGzHaSRqJBUh5vMlC4tSc/Zk47q0EX
rQSZsZgMkJmFYSlsFQRczCl692Gt8c+Ih8hHsNRSrhpeqNjFYOKu8IW23XWwBpA5juVKSgH83Nod
90NRunKptHba8LBiq1SgwR+joTx4RPzjufTC4/evQ9KA+BWS3zEGlIxH3qgtKUmgVHOY+9kveWe2
wRvpieJZPzXko0VmO4gIW2KZkmEuc1HlnundkvCIIf7dFm/lNH9FlzM14IOmJv579HKGg5fm6DKH
o7ZjwB0wXYRjBngeAJO+790/RcnKvHgRJwe982h16WA8qHMCLfqm+s1gaKLwIXO2zU1ZhXkd1m/9
SjhM6ZsoZRmmWWQ6cvyJAaGJMvtW2P8JTCA1+I6MhGy6ERosDPEv+rISriPKNuv9t9+HfRYVthUt
wBdgNPGIsCXSwzidZz/HeVB3CtZ72liN42QY1+wOoehNk3ydJUE81mP1eIqkesL0bpQ4CVnUM77y
R4C/0r5Noe+9Eg1YNcW6FYzbBIIxyohlhY2J98HEc0ka8vd4MRSvrIcSPxuydC0S4D3olJ6rBk04
GZOWLgZGmzR3xgzOfd2V+QscqLbWV+CxxEGfpEbts4k7GdPHUequz/HWWg0VOzXL1rRikwLQB4bt
ZOajJ3y/WlIx2HR6wXTkLbpLmqvzVDsqSf69kgtpZhQrFwjV7Q53O4t5Icw6u3mp4XZX2fhXc6ac
50o4L7CScdC5InKDH/rzZdkqWTduDKaIhS3Qp6kN/k9c4EVNeQGfcuzO8qzli47V8t+NwWEM85nE
czi1AoJFKUcPLJgBx6tAzFJipvMQQJ//JCSz4EStBVQhHRwpud4egf1YsDlmw7gjvIB22lm36sQc
4sg4vV5AEg3hYhVUb63fYBc6HEAouWwaiIEgnnaVJjbPW2UgtZWfaPFcyPue0NNSpmqJaOjyPXXE
AMnK8OeoWwEhxxZkVnlU1vjB5isyHobZiMfs99Xh7+WS2Pknsc3Zye5yvd3tg84QuQa7s4Nelvey
rU6OMH4foisWzU2IeCswrUpuZZeWMtKHr0kBR9M03fzmbWPUUaWk//FPwPxm5rF9+Irz2Z1Z759H
E6yBo20PjY14QvqvV/HyFLKbXPeKsdnaXNalWWsffzjYmmeoiQaeBxmlWHSce8IvACF1NQc1QIhF
wo2UPjypz/+ngmb0qcc2VEmlVG7HwptwbY70b/nIJ3P9cEYgyvbMQ2mbeEBvQa8Lq0db6Ch9T+1G
7LEX04CHtNocEbnfkdSUiUpYXdjMMZLIzddJfvTVRZrCIyYjgm0R02OGuAOUQLMWkOyQDoZ2wjSA
ZVTwpE83YY5wGhDXno8iDLjd51LkqK4dCiOF3ZJj6hc3rxWYWKTtMpcWX95P0bLXB4t96riKGbk1
rS1C49UGvbQbDhw88AuEXxfdrL/aJ7vr/Tmy4a20+xjTt4Ga5MlfvI/hKMQ25QMGWrLyTN2CaUvh
HHCw+66UdyJgiolP8Y9fNvVle+1wNaxHpAvrqMRPVGgM8HLWi2Q8Q3sN/vbA0q3myWTgCB0gdjMn
fGi9D76tiPhQgaRjPZN44TH2wuvF0kXebkyCLqhBtRXNRSb2oB7yLdfRi2SEi90v+9db6J6Pl1L4
bzCV/6mHx4V88B6oMNroCAdsZv2ZNAXaLG+WH6Jxtl6Z8NP9MbCtM46GwuWgC8kniN6RA35xzc/X
rCKcQmWxDJLugfS5HiyTIsRfgWyzL2gJv7OSDN2uAGQRrC58D2iY5e6k9k2PVgRq2FIaMxpdSw47
S2I0VcqITMEi7zKpM651XWkWgu8Jrfgv/r7/7UD3E+0rcgzJS0uZfIud5JezCHMlVhYZcxQQSWme
XhI9egQEp8DNRgIZixYwfGU0t/oeb5o7xaZzSCG3CSgmfBEOefJEJOV1x5o0AABR5VIMTJU6wwmM
m7yGswldvJDPltBIYvwffPJTIWOXGKBE2655B5B7B/rTqoUHRx8cDcTOcz4fjsKX72SRhfTo57dD
l2dNiMOwSsrKIT9Tod/CwqZuu6di+lQYFcGpjYUlYKo8yw1AEKhGc84Y87WJHdYGjGvIUpKiq+Xh
UdeEsTL7sMFI4u3OiEgsGZO0XO0gCgcEOBKwDgYWYY3BzbemKPAsWOmKJO9pfDVlv9wJIrwuLCUC
csjIBIpUyeRcjFfciHFA5TV4/bzFVmlpBouklYYcj6fzF4Z7QbjhJwlDbv6yz62fs3/WHByv2TVV
z94sBS6UZCNmQNFS0KI1WRsNHQxQ0r+FBW66R+V7pva7zsO9PtK2VaMmdV6jB/5uIxv+r3x7QkTr
/1GRwHPd8ufG/MFkW4PGTcBeZo4j2DqGpzgBh9uMpqT/VtNUUZ0426ZxuI8XpMaFrFy4MSq2/Y4x
FmGQfuPXmgT6tYpUs5UG7XlDTKTV2QClrJpKU5yLjLliBmHVWC55aXU3zWOUX1I6cL8JAanjB+D4
jjxzvkDRUvmRtwEoyZE7Su4ICYe+B50r3K+6Ejv3OS6xnkcjIJFSVqpf33sUdcZ33zeTvvHWWYAZ
0c7pkY2OEBTQ7aMpHrUF8uthaXkS2eGN79MEXb2SK8hAUHLEGFDNJ/x2Xoyl3CTwJSu9vtUCCKq6
XVn8WkCCDzFIb4BBCe2NSKb5Ke4PRneChNsCDyGVEwEIeOKq6HKlplT4XahQUcdxlU708UKtOq3T
Kzrw97dsvVAYVrIYeGBqgbrEsFrvqvz7IgmCCNcRj/lvWWq5wPzZhJvpuPWRHK5ZmjjTcmxgE0P4
EP9B06lcTsLK2nHQn5Nqqn6ekOGuI3XKOk95/Gho/LCcuR8pyBCMoLyyt7P21BuCvoDG7Aof79yM
KSHtnRPQUFVTbGDVvRA4pI69Ka8uzYrYqEje76nZsI8durqdByJlEPCiwIP/dapEfYtzUahf7o+P
axnn8euZNr7F4Y9txV9e0wmY6reWpedasrcvINZ0h2cT2Tw7Px+nJxYLT08A8RFaECRl5DEquaBD
Ha2WBvVGhJx+nF3NCLQ2bPU6HehPC7dku3LiKURo+pYuHotXowj77gauj0ske/ERmFyPCkGxOyta
kl1xJcOM8HivgxVY72ZeOe+7JrAIpcSEsdXBZ0M5z3fK4DLXuHrG+Va0Gkk6FyyQcnWamJYD3/Dj
SbkXaShKRTxOCv0D5FUTByo7DuD4X9HF1zZC0doe4PIBWi8U1HMvDgljPUmjS8ioJJTHvASXKhE8
4acXhpoREl5deByS3mzrmfImOnUYnw7a4pe2XBCCzoy1cdrMc+WQUgyCDq75nFooncwbtA0CupeU
HL2dzgDNVoZ6/hE8Hey9DQUwjAlDPrmpaAGZqOldgtRaUvoov+bU86SIJnZwQQryVv9XZa9wScNc
6dh8LDVORttIM/FKP0kG0rS8w/x6/zGECvkEGC+jSiO9c/LjmrD9mUUOnGzJnXQimXzjvZHjJk7J
S++0u0RQtWTIe4PHQpTWPGP9qSuDaFGXY5A31hqcT99YL+i3p4ymW1DvGiHOnozWxQ0ANFeYOCZE
Ro2VeKj63+azQFKfBhUUsJuMWN4Q/h4hZQyd2N1dy7KSi1lLd5M5GQ8S3s72pSEDdvMIMzgYHP+1
W9gQj0y5BkSTjYqn12M0MhDq7+N3cgRsPEsdcMgx+AxZQ5cd/Ihrx0hWMnSyYPfmoPo3jNXGCOsM
6ZpWF0Pb8q4OwPdW2aRA0XXgv3Cyd8kB6hf7GMNnJEjDj0Tl0xabJ2fYj7ZHnX8CeIq7AKk4BQd7
Ay/pJb7i14xq5xybVroS03yzbS7vy6m2+9azg4gXnXo7pCYCBCNZQcNYRFgPFD55y0Vdye/x2Nr0
QKHJKN+I8UhdsuHqsUjswUHyKfpGNf0v75D+XtA7l9BLEyDPlzV7IrOufP0sJc4J0tn4jqFVPiS4
17+oi5Ubojzq55Wv5kNky3CRxPjW8C9gLgE1Pxp3I4pjniIXBPxNfA2kSjzMVonfMbMzmKLndCAj
Qt7WU3j2dOoydcG5e3EB/bKJQe4XB5idgz6CA1vhvIRmnM3qTLQetOVr1CHUjnLJt1w2DqdrHqkO
dBk1smKwhAmC4Jezl/LaCE3/200Yn+WUYeeuLI9GFeSqg2cxp+mDuCbrUg+YvKPrL4UkZHNYT2Ex
PFvjR7hQMltVmxVDjxt5vkhG8AT/c8RslTYndALE/Gwx77OXyzzThzHDLGCkuOrgpft5b+P+9+Ci
KYfC9Cg1y9R61Tj+wlPAMWxGds2Sd2FrwVRIEiiJBSf2Vd4byzZkxLzzE+FXsbasvhylNH55MmGt
m5GeiAMZkwoUG4exzUttqpRp8/ExtMts/Gx630bSFDul3UGCtMxikR7cQBPQ5ppM6wZUM+tQwm54
+tGnouZDnCENdMinfS7kSGGQ5VSPnk8/QGnIHA/8a2sJI/6jb6cLKIhVJFtCsD+yME60guETCXd8
W1Srbi2YqJDRNP56if1BlPFiDk70ncrttcGdkmcoaVK4CEvcFBqAhtL/FOT0LL2Pp5VSk1VcEM3f
JUiydld0nhJrgUEvFDwg3xYDtmJUqtXm2sE+3c2LhLKn4MgosYGZm6aHdOIvP02sDsNdy54NeidD
P+3V7cPco5J0cYHwERjHoDwQmDW0n6YHFq7g9Pwk2NQQf/vm54p4cZfIVnV2g/rDRAyUxa18fL8N
EXyTOQk4/O1rV0sfnjNtN7RW2ERwpctFYcD1kPeafWwjWPFxWvwve6qNLANKiYJQDCr1BRYoS011
m0PjZUbKsoxxp6fiYxUJZtOfSNAdUOPq1YBpTRBMlvw+MbQFujidfUNI4OhiSi+DYt2NAWTLh1Tf
Uh7T5vTWJgApW08oE/llCWl907QxXdY/F19xeuN4duH9Hozc94HKnND6KYNWigZqnXex1l6fNBoA
5Ay9gpibQ0mHYyo831C+fCxu/5VVWaKeI1eiambYP90FrehVIzotBl9ANoZ0izko6BNDg+GpOs/E
Q3k1tRaC+taEKRAcPyZd4YnEBVSlcvk/V3W5DIU7NkqqzaFcvl1TK/NDfhFBptc3yKajyy5fUgle
kzgl99AhurepTSvzUu7FuUU1n1TZYi8L22duQsWVo9Sv9uK2UbDy/+EZp/AFmfT/5CEVKvGZ12DH
VXITw7FmHjx1SmAi9UA+rsn0UrNExJWFOAMvqPWtL0ZLb1CQyF20U0d5Tu1HeluYiuJLK4dCpIHn
n5NLWNqJO5TU+FfABhk95rOyZyv9g/RD0kKW0So/ewOlk65FjUotYdJKDNewapLiJkwbXu7QYiGJ
/To3UyQiqSVI49s9Q8hcB1eVay6HyyUOCu/9SoY38NVG352sSOQ9p8rW+hU4EkRVq8jfiIFMoGEv
Zlhcuvbj9M/QShDGnhBPs70QOdXRCMxLmDJrqdrgeLt3aSiH/kEYiJNzHk2gC5ObjJLAAWrOQadu
3LIHZMzRvwxMqFTqcKUMC6OKSiNMBNCVSE/l2Vp2YpisFAt0a9j3XSNvmrtGQdJ0Pbgo0zn8o4N2
VYViZxUKDJu35DHYln6V+NfKLUTNuX79nDwXA/yT9ID9FFowWcKy1mwj6uUt59XXGiBIoNfx33Jb
BkUy7uEprtDwHPPDVHdCl4w1xwmWn2NDslbE9M78td0vTEZz0l1QobdQDmELoJsJqDAPyyBo42g0
MJcLhqhE9b7L05AsA16t4a8bQomdezqJRiFcINuH8cW5IgH2Gip6y43SGRqLd2r9M7ea9/BGmOWS
ZqihlfRWI1nakOUAQohBnq4Q6QSwZJwA/glMGPf7Ovr637kH/dIsg+co8l7/ddbURe8Jy2BeZsFc
8IXSSwbZEuzqdL6NcQVHld2X+kADOSXYUWJNQD35sc65wzueKmFu2dpelBkQqHSaucOD56FfFjX2
3FsTNMZxV3O4OdN6uKyMX/L8W+eqO67MvASx7nbQM6bi+bYQqtNr+TbIhvuDjP1b8h9Rw3Azlr/1
JLf9xMd2Ded+am/WzmRsS2HMkRuVboeOfre5fk03Zbc5Inoo+GLVhFE/ew/Gjbw+wlErlZ6s7liV
vxQYojOyi+7iiLHFyx65XLAWVIpGX6Exch9OXpr+5kisrxbEiZWxxbCru7ciGoQZ/gs9qH0MghO+
iJfVrySAPMHQ1EtgQ/zUu5iFkHxDUZxO6+b/P96WznXK8bbL+xf1NsAtg2uly5UiSWP6E6LeIDyB
6X3+8OK8hJRkaXT8PsH1GuZ3Y57n7wPlwCFOWw13oraMDB2s3J7yT5OgPrK/6gCqZGBWVYDOPvXp
NOaChPZj9FtvmoeUF0cMyaVgOit6Lr45XQXodw2IdGdOwxkgij4tfxzRDepRjiI69psHMuartjZT
pDRf/S+pUrO9SkTiCz2zKwpEnTFO0XWf4+0GwAdkqwGMOTD5FD65XtK09VVIkVyhH1b3rfsKYP/I
cLhJ9b9UKyByTwO3xhudDtAWiZe08ve6RKY+wuCmIm1SgNwY7q2mPb7esjHl5mlSFdJMJamoX5pV
sOQvH+kR12fhB+E1/WXGr1lfSNxnblbyISqL2j76MLPZtVNrgwP+K+Ao6Ifod5Mesow3Cy1+eKuF
i3PuckCM0QuPIkkVfL69X0UbxEIpScyuKYGLb/5C5QfklauHbMRYQy2dwRQRHtj2MvOCKq9TbLcW
hlLjylNcccoq/pYkgy2tK9hTvMHgeb7ec8Ke2XDdQLhBqEulJF8x8m5e4qDbWryJm1AySX/KkwJJ
F88fzPllY76cM5Khh8DlC6Eq1h5Vnkp2rZBlmC8P5KTwWpZjpPiQN2gbrz/jZSPm1FoJllVOPbIH
jhmqkBGKCCeVZyk9Pkh3kERfuoRwWhIN5ig8V8LE9BdllMvmEN+78JFHbd1FTQBHecSi3SUouFOF
eL6cS1kqKC+PZdJMkx3LFPIH4yXXg8UXKQrSdIozBYyuI6w8Qrb47SZAQ6Hryr1SwjL0DcXBaNVH
1RyhXS7kXmHOoTHmIaA0sLVm9op8qqu8L4sqLzvav57GJ507jA3/5NMK9nQyHJ+2i82aENrq4IRn
lDc9xoMrEJ9/KOpaProJ7OXjkxGsFoRSv4QR/1XHnx8Nn07U/GEP+1Fz4fqXL3QuU053+Eq2XusS
yh8sZsMDTuLtHRxrCMOL+IcejxOyfJLiqhQjt/1uFSlayz96/EXHXZlWqKWr8n3YNnwhbHYzt9UZ
S4pRN7aC1ZG6vT78N+y8XCiCWN2t4q5LrHGZ3nCzXPgRPmG5fT9ToTd+xk+JwX4yvGrmJMNijm0v
X0ji0pTgAEvfwe2JHHxL29hyEzC2qsIbupJe95VsMwjl1kpj0cttA2JN//V5YJJ77xIYT7EiX8b2
priway33Pq5QZuPokLoNN2ZtcnrHD86k6svB6E5zrf6eE6xt2fXlfpTjEASwkNkZ7djOyLYw2aim
MCgpEKN77JH9LsM+Mu9GjcavIC69in63mTj6jTjkyaEHuYXikGc/saaCnWlS+LOcMebKtSmxqO9r
hw0VsoKfi+gy5VM/fiWbp/OcdHe17bPRBBLiTDH2QaN8zmZBNZ1Hg+o5+iKLT/pxMACb5Jcmhscw
lSBUQMDNe3bKF5ofBQXCqZNMyqZEAm3MZZBhu8v+XJBj3g0+e5ActXClDKzRKsUcg8MBcfF+/rJl
obAaXw5Spm/aLYhy3w/QKu0goXkJs1Udc7ulzkmStaQnYLzNc4V4XOqVjbgepo04PbFON3/ruSos
dvZIiT1iTFmV2WCP6tLc+eCcGIVC+6gdTPGZ5lAtdl5xgsT4UedYmWo68AByLJwr2ch1vOMfq7yJ
SLT00MkZ1hlRCbOQmHMlqN4hu4W3mOKT3UCQG1LNMZKmpZ4tINfdgvsbFIR/dwnuzt8qoPAt1+R8
TFVM2E1rCo4kdrSh8KWWSCdo02gCLnuFhJL5okv2qnfBVyFd461fSRnMGccXPP2tqtiCxubXdiR0
IlDXugYEs06OlU1gf5SxGjFjfmzRY7mBGDWGUA2GRQbteLbr5RhkbtZAWaYVx6BesdftcJqHdE1k
9ra8UyL/7BHsA8jcfCUDTU9tqNKgesgmNl5WYsk3UrcHrNfvenjQy2RZ5UG5ywTbCukjxpmmKa/N
cSGmDpEk7wMOvYmLlTfWla9de13CtFZKT5l/9PuTugVoSf29EArFCrooopnKXSp1pyEKBpjldIu8
mTWQvWulUB8qbXkGTZOOoim/0a3qvCDSC4FzfNg0uVr7wd5JCMnzPfh653qV10mlTXT3Pj9UTRUM
GCph82/qp9MYX0ofcj8Ng8FpGBhOd3rnM46vw0+p+qzdLY/iCkm7DltjRnGsQHI1GiFsJCK5r03n
a/imrCInGTA691DCC0hgFijOSWyAsTcaWIyghX+u73ofBkP6v1r0ZvY3w4uFOOaEcEL68OJu4b3i
3snrKE2U2Axh7+2v9aJXmSlmb29rBpagFr3hcLwclNPbRju7cMsqVjg1oXxJcl8Vc1RoIEHdsE91
wnMJIQy/XlyjgtKe1Cvow66nKy4eLpXpCQtK6mEudfIUNNsbBrM8deM5DlPWXrRv9BYC6ZQOBXKx
n1WT0O8CP5cb4nK8UtPwDbCrkIM03bb3xnUBWPSVWckoUgnlatx9Pi2G401UfvB+WjENX5q+OjsS
h3T0WNQ4gynKHkmCS1vpIzsxXXkkrNUbOt/Nm4pnSJ+XnJIpjIVWZg46LvdkXCA5oewQOa7X8Nmx
/HDeUbK+PWKSrjbVCVoWd4EGQSDL0x1mCriuYX21+1zeBtiu9NHqVJra22CG0im7zMF1sx53g1pt
3q6p0xc1IRjm8ZBCAUCqQQmAv+xLT3LpM0CJNm4h8VkmHrwI5AoJ3bOnCAnNelKCbDmBf3fFYNlo
doeB70j7/RHnshXddca8PwyVPvinZuxlxuYTpUdt/64vRIe468B9EaC4JNI+ucJI5yiDzpZ9AqrB
h8i8dlTAo+0ZorxSJfAAoIg7fJjCqD1Nn+spX8KNkdVAq3XKz0EXlE97ZkSeU78/10Ica84Y4Aat
m0GTjDPlr5+bZpqSiGZuqLhD4tlirP2rMR9/A5bU/5VWqyPkD5Q1fgOCiIL+a9kGn4gpWpH7fG2f
4/9yALSlLNmSH4/EYrxRJnKPk+HkPcjQQZkoR6DEm6Irg2g/SJEGg8ewExfeq8Mt1gMNCea7B+R7
ltCzcwAeclaqNr4wUt7ihQP0yGSb+FJUQUNBNn1UI52o+DX5XZ5L9/eAwLJQH6GCMjAWeYCnc7n7
GBP4BLt1zPTM3Unktogn9CWNItHGNf8K8aoFgIs/82gUR6drvQJm4xoSvUDppW4KCJ7GhAxub/Jl
q0fjYmoB4UbhVXFqN6s3SDHvTuVvbOaFm+CnyrT0LUef+Z+m0lYThYUCf4UiFGGdSi71GK/Zfej9
OQ4uYv5xbQKUJs4KpRPcI+vhPMr6v4+Mm7XfPfL+6sa+b4goO9epjW1kcfdLxnWnbVj1kKb0DiXd
Ylw6903rdg6IcolF14oIr0wqQ622KgQuIn8S5z/FKyIjkdtdWurN/1UdjP22fFHHWnF8NM//Hw0g
Tkx+WQZYxqNO9AiscQr0x4WlLg7AhLmtPEGLRDK5ZLXHmJMs954gTJfYBVyWdiX0UyDDhSq2MROI
m4F0LQS2R3cs/ixhf+4KaOWodKsZKYUwLwbmhL0HJiQsE9t4YMNDGSU/LoYaZ5mH3EXy/zIuiUCv
7B+6GLwfFs8nenrydKFPAubFLVZ0ooet9z/Ni+kLAPEvwx7BCBQPFdr8+2siqZw92Xr2A9pk6Vpk
YfI2qY9qhZJXQCPiFI28No3E06Mbh5Yy5c5mq9LTPVbUkgTWYs5toareiuniFl2W5/DZK700L07P
qWobE5AhSAT+Z18UTCly2NAqVPTr2hE3YylA+hOAz+mpp/7ESnpiH29cC7+BHWaFfOTmnh9nYXzC
/L4unlP2aLoLGKHu/bHtkdIbJVQ63rNkBEhiUF7rf+GayyS72twazwhtoeTrQW0TSjuSAyeoFXMD
iEimyIE1PpvlNQKhF/CO7YYRE6FPhU5yxCyUd59ZWfZyTyJRdiB8qSW+wrtYhaj+/kSnRpUB/zqb
5CazBKApl8YzHEId+FlDKvECQBHPKzMqMcwYbbcHgT7iO8841962R+Ru8Dbx2c0EJCdiHWVR2Mmx
7JPV5/iGKM/w8xX1XaX+oG7m5KaIG72NCGfCyy/AkwTjIzbtnPw0OSX1gHFI2XLhjkfiEO+KuLAQ
gVXujAdoaJd4B9zQEdjclgSWGaxavaUMC5KBrIg+cyXdLNR2Xcp41vMuwQLa3/Gou53ggBLf6txQ
x35r1ZhB2jjUcKeUEH9p76XasNTqt4NH0UFRl6lYU237Goxyt8MJTRS5dlkZfPfXhE5gmpMuS8hm
QJlrkPdIX77M+kaZ1dFGCvTkxOgsmmbCYS14KG7BWRpnLUeBzPjl9h5KVYdkQ0KX7KVnahBFSEOW
+ME/tLwYqr6/Qd09P4c5ulYkQViP6qoXWMpGfCj0V9wNQZiRzAll+MtcxKrbuTbakBnkIJitj9Os
0ybcpoOFuSkBgVVI9e3ci4ttSBkVfZ3PCuQsCAkH80fUm/lFTL9HsfUYjJT/qrnmRVKbI0fMpL2M
HzCCU3zKldpKfQy0vXKaIdnzYWmiqPww6m9dsVjhIihNalOvHsXuKTaSSshiQ83ftYVjC7keq0Kb
D3gcwE40qPaek4PXt3igxglTjz0JYI+HIx/8t43uhMCHMbJar3Xc4WWBKD7F/mKuHv47vVjzkt2k
zPxByJFkRKI7YYvYsOa3VxC82zgjKmAmMSRABJU98ynHqI0JVuzFV/RqVd3tsVALX1Mm1aZ766QF
XB+podTqIRSnxA6cQXX9O+zJQ6qdEHWo/1wxCBcdyOpTFo7p2hcyA7++CIthCKgslWj3Blf5tGuG
mRHUP4YG4wP7/ZHv1VATbiBgnfxfR+X9HX4+v8JDi/6HM7rv8iWfCi8JX100M+kAzqQsMcMZSpdr
zVZHIavCHQvbJe1pdn3yTHUfJN9F/LdQvacKEBzVjKXn0W2ywOEfXsJT/m0+CChZ+5/FUfyfDHjr
510n4zQJlxo9sFw/EpaCO67lUxbZO3QEEhjPjVvscSGb+NzekSYcj/mIAZLm4a+KaBYRH3/VAeQe
nqi8/to0xQ0sYPwQyi7hoetCcNP3zpat2la4aeZwUpZ9PkpTJAT9jfEtpFH6Hf0dBI3yph/k9xw7
hp/7wgkg2ze761g/ps6GPmfCqGzBPBmZlfSZUvxfFJzYi5DZM+6532GPj46nsoPnkoHRCDBD4apJ
DehzWV4D65DhCpRTWHwxYD8INx4NrC9nCvkmpiKjVruHuZt9YYPSPZeT1a1DctfWXPFIEnm/An1M
JB6LXVHH3EXg0xvwrA839tOxiO0MGrhq99rbPFPFFRn1ZaE+vkb8lNC1ojDQQu/dozxc40B8qLeg
JUkVY/Rq5vVOUG8kt2zIluMdiO/a0ccYrwK0aFpPkdiuR5ptcwhOfyI/QOvhpxUoWLwKnUmNaFQ5
OoDRR0iJbE/CBi32bZsXdt4vJLCUXjoK1iuy+imGuxzNy2rJeYKzreDERAX3EqhGvwu08/PBCItw
3vI3V8CZmSKyXjMGC6lx5L8BeHUtkmH1dF10gY5cPFffg8tfMAe8uY7F2XUfhX2ZydAmB9d3ena4
IT8Ckrmwc/VjxwQff+4xbtjA43Z/FsSSclpnTRUsAJvbYQASwVBmsk6wSnkoWO/eCZSjhuz66l7f
DvqSBDjdrjqnq3fxSoQAfqYlDRPREIsDrG77YxSR0QsneGfia+qu+JCxwinZ+sWflkbwbOVxIRs7
N/DwsxfgUCZksMDsiTIk0goq/Ve/4BVPf39X51gHcjxUh1/OJZo7kh9EXd3VUtFIMEvJuYcjz3WK
s15uNBCy3AYG7YwhhrrrpNkacCbLqYsYIngG0Y1N3K13OU7fXfeuBk2A62YWd8fzDT86XE6SAY4w
YUVUOj/QCq0Bqgsld3JIHAFCjFVWdJR886dNFd0bl6m8534mH7pPu0VoNZDef4aI5wYK2UA2PqQb
D4vl/1+DlfftL8Vs6n9mu6QOel3MoQR0LqM8scEloM4TH8Znp25rQZdvRQHExCzDygHl5XCINfqF
mSFnwprKcN4CAqdPkNZ6tUFJsGnt3gOnfKiY2f4pdpqByjHEs5tyug5WEGJQgXn72iE+zeSwyn/g
rgP8KSpxhvbruLLJmKSIe/H0G/VwF0l/qiTRm+yZi07V9yxCOU/aY6/wuuGrbSbT8w1Yo7U8Ccmg
us6au5TZHwM+4Tfn0/75UG+iK2rBCFd68lmeV4mzH1+pnhRG7Ndoi1DyWxKFtUTTso5TEoJA0eRM
GPquleMUvF2YXVCUVGo8g632jmts5d0fEZhLNKPaF4nNg7sykOB5zC4SbwIBy7XaJdEAqqXXkneu
mb+l7cywtRkbesyoOhGPE/icLNNm4d21nHUy/nagBnwQGjAbygi8z/8H6PG7nLdQqCioCC6UP1fV
oOIDXpMcmCFVL5z+qc7dQijLCEOJJXvMMBal6BYt6KPxeb0BiAxddoXVFgrXTfRTVZmRlKzy9Y9J
j2uI9cWNKpMpFlkwplVAECOvyveh3yWoFdXGwB+xrSLvw3IUa8kkVW2Dzq7NKU8lRkNacdMfhdVR
71naHEGrXGh4Pf74SehDhiDxGfmJntm3EbmEdHmttPZSZh17b8FPuWglI3QMX5uMuDmanmJgd/3f
K+8KJYTvDUDwOv3M9YurFZTp+zYwhS27L8bYG1Pd2kLdndovQ7hF50SC1SMaOJr/myVd/eSl9tzB
dNcoSuNkLcSS5oaWeIWzklZux5/wa7opfo0vL+JxyLPSdjtKMhGUqBmxx8jhsZGaoq8hMtHfyImt
N09+duiopg9NhIG/3xbnlzv+qW2/gegfhE+rOLTRCEBvJtIbwIW1O7SrObdKDR2JJKhyd8p5XSAj
B6CBXRIW60bqc/BMZO3nATA18Ay5LcsKXMP0NVUW64zA9OL770+nY7xOHvvvdvmi7NrPolu5V/xy
WVewl6iaZqKfeiDCVIQNM6bSxWm1gV3qIQDraE9qj+3TVeb695QwiBkPPK+z8OFOPt2V+RlFnURG
mD0+1/fyUYrbfUvHVOTdFNIdPel0h33k7izVMSiMoMaAH5aLLMOIbAuGzTICoSzUcWgK+jKIyX02
z2XnTNw5n9OERx7CrlsEujDbCQxv/MXNl2AKz+Ww1W+bA/Wdx/BM76EKEPSt1hIk5qls0lJTlqSW
ucYtRWj3jpVMYcbt/Q6UBPvXZG+zt74JkZOPmsuOnakiX7ZU5dMtoxfjmCefWNVWJ80/20uxOPXF
WgFa59YEz8lUxFMRpJyY+pEJm9Wn6qASV5SmCy8ZZTVprFcbkSjzAg10bdSKO/mFW8sdFziNGWho
hau8k0rfG/UDXOHEpTDXrn6rY9Xq91H1ajYbvOikr8Rwp+3xodzihP0Pg/97q8BAw4v+jUKBcgHD
3q34Kbhr7+6PswgJDJsGH9ieC7ABGd9kzj/Tser+FtFYA8dMoyoHmQQRiOt6VBUPve8jQDCUn9uz
F7LSow8GKW/kBwUBix/swb6252Q6WeX/gKmxudmcrdcHzSRORDNxTE6mxP7S7hSUV4t/HA4vHhpd
Rb+3ZyXLtXHw1ZNDxFX/+sZoZ/DOaKB9UhFR1LDXj1QS2uauXj5sbreEuWzpjAhOcQMmrCIc9ZWl
JzOSUc5IvT5Y9p1CAbtLAqoOMcGujCsVZIA2DKZQoYEf6+olkUPbkJ876CTWhmkXW5OwE5IeJshZ
eZ/ZPIeBay/5reReElhQmPw9ZwKy/h06iORV6Fy9p8XTgDyKUDiRBcpvgxQgZLkS+vxi2uUZBv8q
ZF+36R+XkdwnkOdxHh4p5O3gzcZRDsFHBUuVqdVF0uc1K4nKFjETXAAaEvrXjl62vq9zVisgMw7A
DY7HKwgZZbI7zIB1Ps+xX2MiYxwKQEfDNEz+8xVf9Xk5DoN0CwAnXNgmm1nzqOo8rOhPZ44FV8bf
Ds9n8sJiUHcoyVFOLkSuMcCpSUlOLxvYkCkJcAvW8/t5uCO+ncb6n/YWvLLlJUMutmQaYGeDsRCa
wH2s5NKRlEXnxzqwLxo/HZ4BaeaAPxOum0pXPfYKhDELTFmyPucBtFwJDQdYIOSm49wx0eYnxZ/k
DDYj1XW9pTmSOiFBxs9bZ4roOQOdFYq84HiJEz2az7wZpytq5IfHp8DzXj65eGar2s2ozh9m5lFf
pwt0X/QhmMjuG6c/Q9wPuKd/uw1ELOsXxl2emEIPih1xTYZmkvrV6weZBiKfplOXWI7z9XBA4BuS
Uuhfph33swU+VawjSdGTuSc0HnSesOJfUzXiAWJ/FMgc8Cy/JFuqGCK7KRoCp1kt43YwltVLzOzj
qXgbz7hGrDUJpjit6vnLQoeN+7UJlfbxtry7ONcIiEOCXWNWZEnw7VPKLUyLZn7JwLZ11BRj52Ky
HCK9fMUNydm7/yZF3ZbcrKgF4SwhriBkxQ0sGfARr4rOr33cQbmHt+puzOhOXSfYre83EMS5NXwG
FrKFkJ24UulRp9bibUhTHpEM/yExxOD8UwkeSZjV4Kt+ptD7TlEqTeB1MaBFcm41bmlI4YRNDx/1
Dn7IuWG1MEAQTHNilipKujOWIf5/Wpf1lduYZrQZLtWzWrpNIDxdf2eb3Z++iW0/Eb/evd/yKn5S
VEcrbVYg+VylC9dRqGTzOi20qhfv6XXjAFEdRT5wpFTqSLRKKUsYi8VGxoUvPFBDFp5sCKl4kMR6
+GUa+SdI+FUO9DJr1OtJRC74IrtruOQ1gDB+Q1lr3Rj3+XMZtf2WHFotSfodw6455PlPimXKn8gK
UkAuuecttk0DHq8IKT97Z2y6gNM4RRpady2UZ6vQ8LJCtAFXx6rHp50My7RA2naXBwNjTQHF0pFK
uvmbHYX/hURt7T7wDbexw7K+j533Lhpyy8/HOl4Kbbg7beVH9q3dHqcRrI82s2bhIy/mjviP45ih
VlJGeYY4WaZdZQWk2oeMn4g9mrcM2v0Vjetj8iJbN7fP0TTgGbkDu0IBp2qNr58iR2a9ijLaEJAO
Y+CQgS1mB+D2/Lisu/zRQ5mvkPo9bNTNIxB7w3YPkuE+0Z2YelwGbkIIoHHfoDSlKL0sXGlXHcM6
X5BoB9spbmudMevu0zwW9HdDSbMmzXXH6x8HaWCFwb8xiow4wZG4nUNNUc1vdXJkMq2eRvThkrw8
PZ9GqEv2w8BDaccc+hDFvrOCuILz9dboZj0OYSnh1bioD+x5b/bLkuUDjNNrqPU9dlD1QqGAfxzc
8yCdHDp26Ydbr4Bqlj4vwdl0DihkxpnjPAwXhuWLdQMa98f5Ko+yUHxLBAwOvb/Uc2nj+JYr15sO
m2GhQoc5eLCuSzpLE5Fpb3hNylddJyW1k8YtkO5cCpvCBjG9xLa/ioUDhM420UG22z8KcbO6J1OH
RYVKLxIsiRiqKg51IFYx6TQJ6dFmXO3azoIWtE3cvVK2fTqBhi36SJlBof3ZfBNW35GwHT3MfACa
pJeqGzt7t9osERYoT7Kelx5X9V2csealdbdpWJ9Vp8KWEnCcxS47y7pmBfjeIDSaWUxxJM7p9QgT
P+xvhRjYNtIECLSjKs6be/9fIm7oKtufsR2pWxki+H0i1UIAufdA+de9zslnKiUZrZf778hd/H5a
a98J80872Zd/mUeQJXGKbohEHaTRHlMlKgOymLjC2PDVzI9CnNqXEIluB04cKwHzD7Y6Kk1owCH2
HEEHmhePtPXRdGoiVeFbTSO1mmdfePX67w02cIFEDW/iOxfvm5aurrJju5Jw21P/BJoNVQQ9P3OF
80mnMR1fheOoq81QMXiGKjkSerIHTsifQ6EtawvTMh/uW9gy+/fyXJcBOBrnNjanpE9QWaXMTUm5
QiXZyusQIlgKvdEKK67+PEDUjBMQ6ViwSPNoHZ1Fj4up1rEjeipNs4XauAH0Pkz+inhVbYq3eV3c
1UK58N3ZTYVDo7TcQoEb8yT3ouc9uc8ZDR6q0XFlYDCsALSaOYS2aAeslKekkeij1TtLLVYXEWZJ
dnRWQWwReFUnNjaK7jimtTprV+mwpkrWXl/BniiHzAZ7xCPuuxL4ymHibhOHRmBgkDX/llFL5xhM
ppqdPqjJzRqtFoUrr9qJgP45kW3lcr+60DQyB6BAlwETUU5VyENVwIjMdMhW7u7qcOpALVhIx/YW
YrB5pFcvTvdAS5VPlT6eaZV4wtmbunoJUUxRVZFNwOkm1OJZB0H2XyP+tnObjLrbEuxitlXGiW6i
UKkHL6UTvLt9U0g/BCt4wW8RP/ShnPlTmKml0J5NOwLaYgZISVkDGsAgJhJRNuBEC5S9HUwO9eM2
qhSbzAJROv57V1vv0bwSlCc2uBcl5sGhUGcbcdzg0nA1f1JmC62oUuzqRIbbsNnSWp3xfqUdVQMx
4Fgk4CZBbQnNgnKcP5WYQwbEQboZD8haUeP715IS1+swD6Gp2bgkIJk68ojO1k6kGcYTVXGkpE+d
1GmgNxVLP0R9W5ACr41LieRqIsfoTZXtmvW3/tzG3BsgZnI5YwqW2KvPnyIdUgCh9XLhiTYVVpbv
8aGjJ2LXKNChTaEQrFtAFp8nLRCrps7zEGbgCHq+EUq01tm/hjtOEmO1mMjJCx0qDImicAmatpAu
Omm4TRqiYnxmLQlkIpsnN03bi8aQJ54Xh6CpwVYzrtTz7oAtCp2/0/YOr2D87CIVttAbYzhSU2Bp
TtbCi99dGl/TWPXDeFDS+VhwR90xfc+d293m92D1fEWo5FZIKQ3xEAczY3efMCTqvi4swcU+fD4c
ugA4o4y5y3wk8sieXdMQFiIVFIWP876iOaeFl4Tkbq640TUnTAkjBOR5bxhrOhdV93bT5/76IBKu
xTcbiu4JtIFPYXxVabeQFBO/Zb6XEQitcooNSRHZYBRQV3JJmKq1tT1hn+SE7Z1XLsvbVCunKIrM
4dODqUJuk9IHe+mKyHzjagvvKYsx6CImSXAD6c/cWXRTkm3PTkf1udsIIM1kIpxjIULZPQtopfwK
yC9to5rqa7DJ+sFYPkj3Qwha3PvhNAdsCK465YtUxQZd3BWV5buvLrsRS0gH1ZGwfRCRT29Xa3bQ
vKz4KuHuLypHVstXug1JmtPYFovQhpESCJh5njKn44XVpVSCbirIVZjMpd047/b5sEDgZBoXFIi1
K8kyKlQwlmmkrfLdQl4Wwv4qO6Af7yjusT491UXTjISNQCWkvnww37xx7HvWOs65qQuEyLDpQUf/
O+x7QnRuKc/7ZbF/4uNcdreIBDC5Xw26iVxeAWZ0L57RQs4KWRNAHssFTOAsWQpzsgnFtkWPOtKd
UVD9oByIi4eaxlkc+DB4Nbkz8gpCsLMnO371e5Cm4IJHYANMkzQ9/rr5RIUFRyw3dybYysMs/oup
z506k/x6EZ09m4BslzopJYmhq1d7+fIF3JyGV0ri3+GNEKfLbDguTjukX2s4XvWz39meGxhk5s5Q
I2IPe7at9fSH2lUr3/ECEylql1J1KOeSo53HQl9Z2ynsTYRXhL0XgngU3z90B0lsmV+bgIUQcpLF
KbX80i49tiF5AODNnQW0KIqDnE43NtGodBCuKVyu/aAVtEP0a+W+bqZs3Ot0mW6RFG33q6h1klgR
myFo6oMMW+l7+Sh3siGJi9s7i+gnV0FHeY+IU7/he3HDHvIoknOsG9vkl7Sr8B448t8BHWOEDrH3
C4TLOkzPKWINeaYqhabdKkipwu59cW7tmpavO0c6XgpPDdoedXF/Utjugg2GB422qyXNjdFZdUd4
T8jt7iwxjs48E1eGkceHbVFKWtMicrOaaTNse4x42xSNNNtuLeZZxBUozYghCST3w81xWI1vsb7R
dv4AINvL0dxwq3qDnIW/eCAQkXvBrEGDWtr13LPZKas/wqSw+Xsuqe+aFMzqy6Y0yx/ro3coWhD5
8Win5XIXdbDOgZbKTBHjFvuob5FMmwZXRD65cgFYsqA82v2tc+Z8SlVqeV1sf0s9lM0+/KJpSqag
WaGQ/2pG6oxzjvWoKwdcA2b8HKCwWz5YY1QncEghrGWumSP8OdhIvVtFRtbB3JcsGCTPT6iPvX7o
S+dMN3ddN0l0ontx/X/genFBPbQusc5iBS1bZvrzxOI2c0VA78R4GG12p78iaOSjaJKP2U1Utys8
5Rfd32HUjfngjtxjstAKLDKfj/7bq6iaOD5GeInN35tpoB3BYKnfJpi1VZWEfUfXmL+fSR/f0U0j
a8XC4Q6em43FOfVAEifQvPkJ5iisQha3jwZvLtk73EGdUlyHeQXskNX9D4470bKS9CJC+2Fw9FCh
QK++7vcKTHrOmeMfBRfTBWTqic3JHVJW1A1gEQfC/d3f3rgOaBVYJ1r0KdQyoKSwCuZecuDVVoVi
tlrA1wFh7JWTAP/S6kf3DsxSQi3y6JI0raYLRW7rZQ+BreKXkP/eH89njn2ki0cO3/WILieMMUD3
3cNYLse+kjY7FdwzdWf5qOVPxN3asp+qXn4FLclUiWiVv+i0fawCvXtvBovgXxHGftu9WnRB55sU
zJ94r1oQzP0GyRFuRMkU9I0PV2pdY98XgeVBEPy2NPLrYoKVxZhSzuRj30EncItopDyonOrzT8jq
glapBi9cmIVM1RhbtRFMqpu9QSfqwFYiFnmz7oItOzIp9Rn+gBt2Udyq0JX5nxNCo2te7YQFDtZp
HDTKNDEiY/sURtBOnhAeaATuP17ZLQjp8GbkEhJxFQrFWUi9ljQ0BI65oXJkra7xH0Dk2xQ85xJN
elfzIGtK+3uojKHShIRNf/o7KxUta0Da94Ngz3AlOb50huuiB1VvBCkL8jUmE/WsSgkTAzHU2Ioh
BTLtR6eB2jyAV1RFTt6slI0jAC6VV0lNuOsQT4LqvBBd+XCd1yqVs4a57a4njkOhse06/IiAnN+Z
LL0yIwqXUMV3t7qEK3+zf8ILRdhNIb1YdIciSEBMfp1vMVwhn4cQd6e6Oe3feeRSoCibGC22Gm5K
TUw/bOvn+pZhpJ1k7Nq2CqmTzh6Mr8+nPz6lhSOwfqVlSR+HBrZIu0ourvn9rd0yEmvSit8fHw8q
icQlGfvZn4M5i8p0Km8bkSEZ80tYSnpoDKlI6qUxsjLudYLfD1qUsexaq7w+5Xln74pllNrLcETf
B2bIk4Rw9sqf78YyXxw36EMIOWuF48e98bPpqi2vlKJcu1O05Cp/HUSQRaMDBYsyQUNqdgNUC6Lb
x4Wb0PCn8JEHL+HDUYMbFLD14nzIPWwchLIIwxwU8HrAM8PSoMfYfOBQSewd5lRn7s3l3/8xVBAF
QkjHllwIe44X2LFTMy4CkVfoz/OZb/MTLFomqqK53N/8pWiXo67hlcx87VK6LwK2n2vweorNhBtc
48M7bt97mwGEMvoncNXquBuC3qddL3R2Qzhybv+dRWN8CEJubgeuiqqKFmtCO1k4K0cxHzuFdRd1
mKE6rgzKui/uMiuFqd670bMLuZAxODaW5eg8u/5KoedN/l4B4XqZBXnhNOAlWaTcQBbd18sXjfUr
d3q8uFKB3bDn5Pq+nbkGrLuJmj41unnhm7NGcv/VP+8iJqmjgBR2fyhZPrxWyQ+bPHchNglK7+fB
eHMfdZoEj+GaM5XwH/z5ZZg8jbrbyW6uihA23dPCj0oKwVri8YA5oH0duq4zojM1j23DXX0GQ1Ki
6kNo7cN4VGIdqHnUAeleP8zSc6HbMpGb+puz8AD3jYFoCbViwE0DZ8INLpmyKM6+zbDkDlhMWgLb
5lbUP6IvkUverA9+xhZhwlV7uF2ajnz4ys7p0hRMGygkiIq2c+Yk6AnAHEtzD4j/KkzvILHtcMZK
Mkp82EGPsjs1PHrT9iS7RHoHpC4qeOTVzUBnMAyj8+kDYxN6u2p2uEzTkqLbGU2OR0EVB1hfV8T2
ib/2n0WF7BIbPy2QuHqA5FdNAnH2Fcs6VTeTsxc91k2a0Jx841NsuXEjV4/TIxmt2CnI18Co1vm5
Ktl4sYcXa71VTGnPn5me9uL8arVXr95NLln6xrnj483xfTwFtSa4As/g83f3wZ7jP9MwG2pIkVMR
Yu1eLifQDF6eZe4Uh/u89W6QawvBCQYCi7UVVzll32bEmRLhkVqPixXoPg1YdDB6QC9AaTrP6mrI
WKzVlTIdCAXlRbxr+AgEq1kJczNW7DvyVOOgc9HuGFE2g/n7yJoyeaiDecJ7zOdY4wRL1pVumjkv
Iu44ZW/bITqlm2jg7OsCBBAJO7HYEZtnVTnPRORteHIe47BQnov1UoGhI1XsGpNP7YtIRyd4QBbE
6WXRA/I5Zwy5pWiX/tHj6rvkO2aFaMWNSX4oQ2dcA5rmoGE96RK7J0mjXQ0SwVW28kE9gW4Xa54u
A1bLRjP8AOvRZY4dbY3hhKREvC/4L2ClWUrYB5xxQPj6nysZvjj6rpcrDUzi0jhR/3Ytt341TBmr
YuqU4oNHQgfqABT5ytAUI75EuVrHrxEb4dGiJuSOeBgZh6aZvcAUGWj92MOz4H9M/QiEi/43SAIX
mVFjEIJjQOohxrOcGyWggY2USxLVprjFzTv4FYShWPbE1ek+/e24K2VWnM9mLaJ1rlkdh0gQ8hEg
nJ6m0tryG802dzWpkz+/fUAdU7r/ERvnhmlC5CU+0uI66WzL10qByUGVPTHh3cnu/+TfymRY2rHz
Q0/leh+i11NjVhgW/sqB/xMH3ySEQ57CHmMjXat13eI3T0FJo1cFzkk+dr7oXedgWO02NGXDQjsE
tc7LZQBNtZTT8AdLwqoWCbfwzb7D+F31IIukZ3eoXmoNnz/94RzFK2y1L+DclWiAWGOwzn6kpzq8
vY9rNKIHixonq7xFJJknn4K031+Zg3sj2S9aXwiUbrsQ/o+6zbS7XfeAoTWICV5/CFYOW1zYI3fU
87MbpRweX29+30h7YXD0fDCg1vMRUkZ+Wmx48X86gOba1nj6E24FTbTvreX+ENlWp/BfGoA6yqBU
uUSIzSyIm4SPPyzlsEBKfxXacUg7joPxe5iCwmXC3+n3Ik72ka/+bVDB9I5a8TiW1l4TFgWiiKwU
EYwscgOfjoYpaMhighHpwrDPBpozP2mojYz4IJdQ2fK1jx+yHZezc7BKcYHuOeV2zK7VONRiJi3y
nxCmXwS4+u1EhIkejKizWT1xRnrSmClk/M4TvSsNb1GyiHltDPJ/pk3K2z8cCrQ1y2gQPnm2zU/7
9NIcOG3qqIn8JrQJ4HKvu0U6l4X95CI/rtngKz8EYMVYPm3TB2APWmp4QZUF2qtjOyMBQhddlJU4
JsPMASM+/A+afXAKfhsgdrEN5OLggBbIOmAt55hkWVxTCKilsuVj2CJmefUGxXAitO99nDmWgrMY
2P/dSqoiroonbl9prnm9GR6U1h5jr6gVFd4fvmRtNqGMMseg5y7/BvYUko1TqLdjUU/VjAX7qkph
YZNlRJjgCy0ZzG4FsTcdl7BlkjoyufgMFS86cTRNYeBBL5dpPZtd+nkCCe/DwPO7VzjFoW5h5FVp
X3rH9IPuHXMT9qQ78MD40qLaqKexa4NyA8d8VWr2A1vJKxrZphCryZVHPVG1tRdGaVtNqLBO6M7R
ht2VfIrau8Gyh35SXYFiAvQAP08wnaiYCS4lhIRNulphYL6Q8BqnsqUYZZR9tj+AW3hBtNu3zDAR
EIaOGyDGal3JzMdvj+PUxPeZNHpiziiDyZofbmzOL7xktp6GkBcVDcKjRUVODzzmpxTRLJzMxmqJ
AqPNq1FtFnzr7OPq1itpmr2j9gHYvPJ3AyqlvLD7BVNLshkjHhBBH2+XstLdZ+Wl6E4DhkS8lklV
D94R8wrlvC21GUHTqCFif4rHGpqjcMLCtI4YQCtZjaTCZ+DdehMGkHNhQ8rfYXST9PdhpYbXT/M9
HRU4I2eSeiPu5K2jxy/mki+kef87rrJJ6Z1SSE0iS7WOL6kRDri+CvTN42nt/M/TNbH8BQEIr6xw
rBnhTFd8NeoaNenIy8xyuQD3HAjmEFTpKV20XMW1wgvRIPLwNTxfNTAeEi3DA1KaGaPLb+2FwAOQ
5r94wyR3z8SV0PfERhlGFx3Qo3uqFZgshSryimsyNNOKWWMWnHwaAyAH3586tuLO2s0audr/ZsN/
kom+MOK+aIOnjJXd9LWwQM0CdT5DrT42Vk22l/hXjZrJr9vJyG6+Zb05hKGzmMSl/d9oGIe6yhYQ
KMi4HBWm5f9a3EnPU40QC0LuVS1sn0qnxGlRHy+ThDZTsTqVs0vl2QE2ItuiomUFIw3AJp+9wtxL
YTfYj1OAAQDnUn4x0/OpOWu1MTlqYjWCgQLMRhDve6fo0V+XuUTNsqgQhh86lA0rYYGWym3GltYW
C25WxNjE6KWwZj7IcBE05LzS+zS1tReZ5+Y8dhlyFuVaujahdy3YeLl8v3uDW6Ugfwm1Ctzh7Qpf
6hz1tBJuxdtU8FviNrfL2JRiz8vaokdaHn/MU5bu5GHXg178UCM6QzjCH0ba85z0rGA8p1Wg0R1d
08Z3epn6656uUxPhacwUlADCDUfRRxna6qfP4fmPAW5ErdqpU5w4knjWLu5b81VuLw7z5cUsXsmF
xwUEpekwGYIqkDOCc9yK+NrMIREq8uDjBY197heYuMOJB1zTf5vXbO3J+iYn1xg0qtZrFu86jfzF
QvG8QplyuZXoWhJgpp11Kr51lZQVQ5PopFBetArrc6A64hBsMAgUF+cug5wr6eGsj7MMfiVXSxih
KkMODZ1vIn2sQSGlG30PflDUeiatrehDkAFwXpMyCBOox+tAaBnr30tWc4AvlFGNYDNFlqqtyCfB
kaKmJLxZxKARVkYLyTpo2uapFKbjT6jUkLPRzWiM0r0OzZ4qeH0a0eGEfh0sVF/9702CFxI1W24w
JIcgVkTAJ5jRZP7hPG8KPLcSGyt12mKvfCtFPt2VMmliENlEfohYxLSBNoTwZ13eRr/2/9hx6V3d
KlnByOSnNkzAWCFsXzKioi2sxOV+NKVeDrFQ4Wl2E22CG70Kj3uvqiwF4hicqrAZAubHonQu1iVT
l4l32oMdMVHcwg3a86avPq1X1dnGMxlS06IoSaMeQPgbGxDtcEtylcHvtSoC7ZDCLTMUgy8EFBvt
piIDWtdmAjldYjjTr0HTFIDJtwGXuqVXDGZK6MEfu3roNcficMgjzTYa0+TonwTDEpvDyWL96zhF
3CpFP4oNPE1EWuV14wRbwe3eAF+IpHi8PIzqm4yaUOXDFH4PEax2FL2l+lNad6kPDX0+37aa2XW/
ErFpkLjkrNp0UoNXKce7h4J0B3UgWVpkPFXwh7RzXtQLkw8YTSNSGdNqO+qku1QRdIqRoEM7kQ+1
/V3+nqbzK0bGS1i/nEzZQ3JYNrjsc6WBo3PadWGycCVms7QeNxGdftNctZTD60LnU5JrqiovXm93
rFUE+E4lngjr2UkYwA++MxSnx6rTjPgu3gcvS5ZaYYk0CrgWzDXMQpyTHeQgx74v6DYFummgBftX
e1Jjkf2qZzZaktcaYjUxG6OT/APgrLKAbmHTeER/R1WqFAuyMYl1zhJWJFmyUNwLHYdHC883Ah6g
xCW8ZXTBDsoTiF3xb/K4o6RiCpDCVEdb4Bcl3ePCQyXytfsorF/SHOumKguE+j1g+KtKFb5+LIaT
SA9qNbo9ZG1h7d/iM5XHCMaDGYeuZll0Rl8rpYhJT2BTQVQ3rYlTIyAqjvRighy73szanTMY9I06
jFvTUX7nCl3w+p85SKmNqV7qiUGDgzZz69YPW0sbuSwUWO9KNy6xJQRj/fFRVLnmbBm0rDcqRRfU
kd0oILD/Dokyx7Lz1hbVXUmui5oUUCPrelcmbvOskYKYsoaJ0jWFacLcUV+ts7zAh8NSmrkgHnUO
Wq4aVwiRYFcjCU+qzzyH6u5La98q38BDO8OfEEDl6AEmbJAm4dB0/+9FFjgCfjTLJvPIeIyvTwBr
+boj/6F+M6jTfb1dbUL/PQgA8EB25IuULHXcmq1v69K1ND2PXheY+3m+WTSCd9HQFCo3+cn0/F/Q
oinLzIyIoPUUWw/gWH0EVAaMvV8jYMy/nXDYwLAjFYh8Utr+IQgI4VvUrpmFgvLBCBJY9VD2sLOH
ZNQhF9B7TjRr53iy1X5WZpmb2Ke8ZMMymqKOYuF8QGHVaaDQqPWTaOEyGjv1pOf923aQ89Fc4T8i
s40NT8dAn4jz2gMp6MEGjyj5FN/cM5lxeuMXo8RFt2KW34COwqXMy2KXR6ug5xw3bwhKFlG5PL9E
HMGOGwWO76r9aEfPxm19/8XFFrFcB8XsvixNpC0JuSLYr94XwCO7DH7dLcqgHnALIPLOV1UgxTso
oP52rjW6devDfk8gQWspCNZdDRp/b25zSPevGWZiV3K/xV2JKcRJrgCS8Y589ZpGWYSGv3l8pgYi
4pffhVsW3+6OCb4ChRddXyxzartmrSKo+5+UqZyJD7IQEFLf2PKNodwVi3IMO0VA9wHx231vfzQW
9GRiAfFZOY+ZEJgTHR97ncAybFnaI0b7n40XXUJHrkid4sFwMSbvZjbw4rvmuV+y9RxSEeb3vPsX
W1ofhAMjSrE9+TbEW39vXrPAlXHXU8oKbrUA2Sdgu1SZrkVzzEzKUlCRj7h554RF9XjgU3HKRvCF
x7zPSIlEmA27wKdNO9kbhkHj+iR0Bgd5EV4NnnqKv+VzpsM5RArylXjbjJg6UFK96BMR1op4BVT7
LBr0K2T1DWc4YZIrfH0eMloiXWWxRPTjUgl2/UZqkxBdsTkFFWqd1TY5w6SvDpAUyyi4BAbVrWLp
zvKjreY9t4AXZ6fp7UJQcRNAGRDiNM3o8RVsFM8VPjGza1QDPEWk1NZo0/gcL+i1mo5NSk3fYKxU
SHCO3VtwaCchaImI1rZNU//ZMf4GJgjii5oDlbIB4nW/R0aB7K5iGt98zmMPpyXIE73nij/Glq3i
hhCz6ULo+HzS00KZ6zbkc8ZAjbzGirpf2k8wEOADL+p2qWRjZQVr1Ph5it37lr5bkNJ3CHcMp3dd
2xstfw57pT7PDPOaqN0iCDRV2YoDSCg+RS9o03bBmktaKwkKUSNZ3Z5LZecjCspWyArfiWnjaWli
X2l70MP8Gh1kY2pfBjgC5ATzxKRblOP/hwPWRMHfdSTtYL6WFn3h2MpK3EYWbgbFZE/15QX9Qtw7
m09hIrOjBTayNW0F6RCrGtGXzgET2O7dU7/fJ/GPAvN8wObp4bZyLUE4Nk1d7ZBdl9bNzB0KeqDo
+GpRBo98fPFr2tsIeOmHtimTa9ypXY3T6SB2m7gfYbIxa8szmuICMXP6mhdVXFvUq6W6+iVtLNnl
QWuoy8FLeLFzCd66nmrJHn925yiL14E2mny+hh2CY4eaTR1avQE12YZQC7KEZJQgiOMzLyKIJVPk
0WZ/8P+8icFp4GKzZuztapmI5Un/KXUxtqwqCjAvWM4V+ITPmWE+hqTX3FPBK+wFvJN/jQrleGXx
ol23aaE1UlKjbxOYpKAjtMYLUy4+EKH6Io/TIv6UKcpHq9W+8SuZwo662ljJkcg5i7QvosEHk5y+
54YQAkPo8HDeHvGUOvrZQTSCOVJN8lzMoOz37oyOpf88aMIylb9Vt1sB8uRqEmrz9b2nzThMxIXC
h2Asjb3CfPIxLj8WJ2g8zO2tyJu0ijoNoZtfV3W8v6hN86AXaIgQDC18aWIBe6ZTUdQzsbqKEXN4
MC1G3U+lVir2T39SvqEGgRhIHE6coP4zWu6pcZSVsuYCgihn6Yh11X/3yLzM3cF5YadEyPCiZLjL
Nb8jdeHyzDQ5oJzFs8lc69ytRfhloQ4RRbUA3lDAHfmYXtVaM3VNkLxzExwsiU+afyQpEQRlRyBG
IDBCPXVOEmLYUJ9vUVWPlSPRHyezhAe2qb4OTp4hNziWzip3IIn/ZfwcF40WxlZsBQjr28RxpZBi
HU6ST0kr0K92DZd5KS/Xt4uQBnOpI51ksJO/56zvCtNC2yV/79MsOCQhRFyUM+ELBEfaDGCIPazm
QGnUJBp/KlR1z08y1ktbPb1T1ot+9DNrPU2awBp5nPoSmZumE5k2jQ6dlOBTpvJZFgoU/FEGjdXU
y6PWoMu/6A8RuvbY/7zo01uA9xTcaoyeApPKtX+TdDZ2wgotLfR1UcbdqiedZvba/u8+zY8jQQO8
jwA44P9nsg3k2DKpeqcLSTpEAsnE96QAjbXEIN6NRYJ+9W/VBgXAqp6jXrfVRUQXluMqqPUoQDMB
JfWylkAwEug5GrLnurq6ZVyTAc/sYXLcze0QTEzurcwN3swkJ9wwgEYOiWXkFPyy351tahqlgNJU
7Lv+vW9Lqrhm7GY2j15OtizeJlHjrkF6FwTJlPks5QZ8Z1mL7kH0kJFCr6cmtWyAcfjyUgbdCIVA
wxiZUR/eHrFQVGC8Fih0ofHvXwunC4EoiF7fuoP3aNImwEUGV3BH10Rkyz4tFlTpCOoBaCWp3aEH
yecQZT3zP1V2NGbX5ogZUs1AyC+bFwkEpDh2yUUiQuEOePBrlE5Z9KEcX7msXd+7OESwbp35tzmX
D8Fr+ll2HHN2CX8kdigGoWZXN3sbTDIOMNb0/Taf82Ex4zfHNFPnjHI9VgGsFlmET/1gKhpYgpGC
ujWFMY5v8F9chjYDf4GeaOdxA69KryBz/kPXaFsBnF63g1lKg9wgnOdYVw2gP82iZdF8aDB95Ua3
sMbmK5WFthmghAsU77yEPLJYpsKOjPNVUeyltKPv884TV+0vLJ1ELqJQf1azFGbCxSkq5mg1vaKa
yn4IGgX4LKlgkqjF0CLzjy/dm53QtKMluAQ+Xadfjxwz9gPJD6fQ5mCg2XyPINLvieZfczve88fN
+FdoMWKYz+csjgz/FXa5hispaqTyqA3KwwdeVhhTXAUe1V0EwBMmA6RIsPcvAid0CP1pmarthq/o
tnJZJA6dC7qphiyr3zFJV57KkHHIR1mFSBYWo1jnJ88aQ4+QHb+gu6Uo5zUhPle0RWgQGxjTZkNI
UIUVibYiKr2IcI0kLPO3E/NFjyHQyFr0+XOR9gU6mZUg4Us6qv30UWDYzJiyqPHMSTHwQYJoJejp
mOhHpg4pHEJh6MQPkmg3lT3F1WPvaiOFd2g7CTXAtTfDLnTgzH4Xg77UU7leVnRknbj7JAS/89YP
R7UOFo54cjyfWj7aZB9M2f/xjfGICnjuy6HwIzB/NsqOZsyAfMYKb4r870WWQHBTOwuSSmSmc1qV
B9ZswUM/QsPdf7BSABLBYh8DKdBO5s5p1AqUEK0BerhfB+zFhQJWXr77OTTc5OaRrEzJqheSg0ui
c8+ilhIDrG0vbxm/Z0YfVJsIe3c1aQlYqvptjbrmTv6ro4HAAM0Jsjjmad19VbMKzD3anp2+MH1u
ogpHUkcrPYYU5LM1lt9rfOpLNx1Aq8ka2QDydXH4YCk7gtws0xZcdW9x8/bc+9BypD9nzB0fUAJe
eIv745PClZwWc8w33aDe6TRfTTpjMYSNwuHd60z2BeWUfka2BSJ9YVIrIjuXeKEma4OsQ8sM4SJ7
4gPUbiP0MKKK5pU1dHqfXJ6HfdiHT9XY02nzkqGfJTl8ojl8sxqTwOh4lbzysIyI97aR6tUTVHGa
mxTC8nhOksOe62X44M8KCm+KnNgk7vj02JwTExKKv6Nzc0myWeD3+7qSZWpKB6nQuhgTi4OwxXxT
8e91xHX+aK0MMHctpbOefifILDmzp8lb21aQ+0Szi/OJCM9UF1kDSGqTZ5aB+7dqHJ77PvagHc/j
aPVKkTW7INUOmEs1G9V469lOabWOakuAmArXVf58GhQ/5H3EJ4nXR4KS5pSZx0XhabwCFMBrVPRQ
fdqfbbZOuhp6SlIATw405KAjKSNrJ3q/YgKs26jocYWXqaTX03fEKIo4BGCc1Ng4UMrbwwncGpdS
iBCnRF1rbL/zXJj9EuOushqp0vntB1Ifwrm2hWnsnJJA7fiMx0O45LYkq0au92YUrpKlYhHc4COA
sfZ8oW24vs3huMxmFOdmuI9qHoSubQPAo2+KMxE6qDfGFK+gnflIet34dvzQer9lkf+q9KDijaYX
Hf4xqg8TqjGXfiudEA0BQOWevlQopAzwT3SFc1S8DPP6/7ZBROaMLVdu9rscSg131L4qFnvImu4I
20CeXhbFyXhG4WzZYboVkSSHvErsmIZj4KnkRM8M7qA+v/d6xhQ9okynypwWU72Ss2YcmN5Ec09G
T47ThmGMYvAjkgyEr70VSen0qMdMfapVdJrmFcXa6Mkxf2Hl88gP/HsvAV8wnhYJYPUWZUO2Z9/v
NIcJGKpFCn1owJuRVKtz9zoOskBn2dkNgDh0hsCRg07aEXaP3OBxXYHC5zsIk6USbWFSp6W9qknp
YxPUJ9/JwilMx8lg5gAneYEi409aGPFQF4l/Fum8cp4dOjcttdcfRlOmeHoFrgprtLYtJcnzmg6P
UWsjtkzqn/VKbYEX8BQJXgMOLubO6F7jMdPgH4+Bg5Mza9O6ThMPkDXrkJqQU4LfdpvdUgMRb1dN
cThssROcT2MjccgzLELedLT33/gYL5uWMchefM/dNjCxwT+KmCgvZQqo1FlXuSffm1CUFswfbxzI
MAI5HvrxcASVVlpeZMFeOaQBJyrJEv6QHAnC4NnEIqnSAuk1uglcgzBPQDzz9qFWKov5ffm8MlUD
m7vNq7as59aAjSi8Oq0hrB2zzQXCQ8dyeOV619ghbT2i5j97e7vI+F0ecwwK941Wr7w/FCXoF0HS
SRBGC9AL3FN7JC2bKFnGPHxW01IzrC9AX2SxVP++Y5RkZRMVpfnD4llHFJg9Q1yeFuXMyWjxMYmL
KR1wCITEOJhptym1ix25Ap+6TGbpqMNhbtJNDvUJGgvmqRyzwN2tTVbR+ohBZ3qdiRBpEzKB3mul
rpkyk0v7fi06gTA2OgQOaPYQ23mqrGPDQ8Jp0z9ZOKLH5c3KP0eeg9mhYAO9UYK/YRKXNqPWYsoc
4vn6DUqhQ/RUpz7UgKxR3HRv9lM/Uq/gi1sGgiiEKPv93p/QelTrR+PigGdHHdGKqO9Ty8marb4n
eUprp5SCEAsXeUTJfoLOVSJ9Yn0Yf3HkiMExhh/+K/glwk6gNZ7zYFhlkPXAk08z/KVzggVcwtO8
ADeKoBZakljxHF3NuwY2/9KdjdUbDNol3AoEbLRpKiBOGqgNCQZJ9G/AZOfENm9ipAtNWnZ91wgU
6LrQ/VLrKaaW/OcTovQfsVAzEmkLtvWy2ObT4Fkz0PpcVxCAGsddPbUjh0z6PsHeBitl/7h762VS
qNuYJJ+P2IvK0nESo0jSqvTqI//yjfLGsUaAAp54D0Ak49sRJYsX3cjsXwoLkdFQQETG2InNhops
UDnZjYFEAh2U1KpDC8bWJbU3LfCkdITXQUUgj5eTGvk74Z/NybI85BPRr2AsJ9usse4bhM+71KTz
ziq2Xahdg9QAxxr8apjtWX0uQHeAR2YtOHcBpHcB1o9IxGvMdbRgazcc2ABOLWyDetnKXYy91SZg
zMu658WQa/QzyN24GmtZsQDlb0y3vnFRf7SqCsJctrTrMT9ElPlLMHQEDtLmE0JSE9xKymgh/AcP
RNfVIeBtB3893rU4r/tpIjPjtT5XWJHYRWvd+XzrwPCo9jXjCl2ElCuEk7vPpf0V+S64552qEFhr
rcL/Nn+kz5K8b4Q0SBWjmgL02cfrUXim0G0LTbLMvQfNKXencljJ/6v5KigYFjDwNHY7f2Buffhy
F4FN7Ms9AWiKX8Ee+2Pm1SFgMWisEtSLN1wbjSOm5atYoavcmZsP4Y7v/caSf8P/oO7USmdrcBKa
+FD9c45GkZYO6qYPj1egIMxRsEbaGqkTKbNhfaDZqjp6WtuVh2mNY7mp1Xvdy/N3HwKj3uDu/7RV
2UN6d04ypi+iUfI7VuXL/mJF9A69F1tYvFuyu9JdNTTXVjsthkI72kfwQQDrwI/oWZ8RRYt0xLem
T0Y+jXa+ReBLDzI+zvjnGQ7UAxJaRl2lLpbHiOhtQRlk+0GoFpkDrkPcVKEsrTS1jrqzBodzxtbV
ilezPO+20D/av2SloaLE9GRK3rBsPFINPR7gtn2wG+I0Cd+uo54wHTcblSUcjTzTCFxunwaf/qt/
VrqpBaxCRwbAxyhiE2rEmV+QvR3Q5/PKs83dtS6Mrj9kYpXZfDHA83Nl6yfPxOCYz/4GhH1kHHvF
uWMSwVhJh99gVJc0bHuAm09Cl6du8t6MVHaJG/JXIneJdzjjDgHP8q7gHDu5b0AKhSjbDLmbJusR
2ES04KAtN7jqUUwfq5gvmKqm3czoV6f6ZweU93xZYTEKt66ibxrnUcK6FMtv2SLDz/tHrGZIzXVA
ZDGraHKh6w1l1DP4J/6LE2qP4br8k/wzvfSX3wCi72PvnnQUD12LKzFhTscykWKXseTqDdJthLJ+
CRDv6WPB1QkupUFkoOo1SAgRnDqXZG5rs/DlLJowIeie/MQhQ+wX4ItZMojxrNp+KjuBdS7qMChF
sV9nmGZsu08rcdekl9LkprxcH7BToOlQGzSId/ofyWncQZ7PPSBnpByW/OVNS8KkA3Z7VmlfIBDb
BZGPtiYBr4zNplU1/zKGcQietHmrstn0WBUX43ASmlGLDtM3R2vPhiQIdBSGgD+nuxqnIFCNgeqo
EAeD+h1H9ttjY13PTzsVvfNbrE942lvfx81sOBnxPdApEoxpKkLM29m7cnNw1gnx+kC+nu8YLsfw
MD56x36FjckVyI+WaqwJJaBsf4EvjQB5eC1wBllgp2214yHG00QTh9/ZOjjDd/7EocoHJ1NatH0U
mCZqfgsL0CekcV/2SFs3F/fYsjHbvFY6TeY/plEiFTh44di0SlA74FC5ai1qwsdtx+PQhxDz9oQe
Ej/MUvepACP/NjUAidXKKtEUl5AvJG933sb0coIDQV16wKaj1IYFMXEc2/XhqhCBnRx/jC/ahnvy
UPbwzZ+zk0BNn7Q6XUn93LgqbYS15uD66e5oRNpYQ4VkE1lfIZGj5JUciFpasOIju1atMIsq5jyK
yFJHJYCcTO5Rbfn/gaL8RgfZ97Sf0dPysrmnRRk2psk6RFTQJ483ZL8pqdGPPONC12sOlEXGfKuf
M51/Zx6JjYR7M2WEkLN4CAY5pyDEEeahwEeZOkI3Roz1WXoHh4xOJfy4yz6gQ6FRLbKdGHVRZSAU
l8BVSprPisCbPpWIm1XWmw2LVtUO/FMQ/AZh2ZLZ5uMaJJ+/3wpYhNoxBAZZVa1wPWYxpUXJMV9B
IIbDf/uRoAvMpewUiVW+RbTrjc/szFDV0QxsjTSe7aweRPIcugPj6OTtZ9fRRMNEE+scrf2h8Er6
MMXZCtYAb3XLMV9f5MGDsM18ZOokk93XSeI9pe+IIu2tUnMcydND2iV9bmzCiibqPmp7rpl7LPSw
v3pugmQR5eCI5v9LjPySP+tKOyDQkWAfjWQScp0Ne7wFbq1hHujh9ZqJuXktkxJd4SPgXozXyod1
CE0PeOAzl5ZsWr1Nlx+ODT7zd0Pa7H2wm8YwL2HUPMPiiBnG07FhVIoYb0frmrTSo7y4lt/P6+t0
kbBlkfPm/KsxfWmkm0m62nvaevUO0RusyxncTjGmCcNiVhEFF3D58+aRLluupUv8MN/uHN/c6Z/v
uFyMKrc5SRDQgAvqKvOlbij0hi/oHzrtB/ffleT6gb4yZrSs4ZwNmrKAy4eQRdWp5aZeVf3G8ceQ
ctNaq7YBgDPkKZE0rgWxKttgAM3ayKQrwtTKsNxXstKdDy6uDWlNH1SGbizM4fL1mQAhLFT6qy+X
k0OpTmCtAvSoQo81+CJTyN254qohsGvc9Q9RzfAo+OBqYqYWONT+BDAfpkyNuNqoNsbeU/poKZ7g
BrKoAJV7HIhG+ypGCnP1ythzWHsVwGv1KVYkLc2THakq7S0N5NO303MAYkPjvyPmNExyK30Ey773
tpkjOyj3qHOfiRf2pm8Ke9Vuzho0TOx1aBbZPyOeqA/YbTrgmcPNWidqkp6YfbYwTd3dS5w0WiNB
w8YcFAGK8rNI25O1gvmVzHD/n9ylqFwN/UnyAIFSOkEtJFqagJtyWliquO0LqP+izi6ei/DBMUcQ
JQ6yuzZG0snmVmj3nCFl6EHHcMnDUf0kLY7PlILNd8ct8ifMd+HTXNA+I9AWBy/baTbki05EU49K
Jd2+yteJuqkCwwAP2MSJkuoOOLU39jL8CYQqZc3BoWANc5qn50P0vyBBdLmzgXIZG7RhHNjT0nXx
bsCcP0PyxQlp4YLFXE6EuxbSlBn7pzTFuADb62ZdRCOjYh3ahiZpU2zG3usccPAJZLTAU2nVnNya
rU1xwLX1gpOo0C0aVKtuQ4mnhs2ECNdgMOqOTZ/Zo8sWpt00K7HnWkvIfp80rCL+6SpRAJJUC5M3
tvKOKHkAHKN/7Q4WCUFeKcnDZ9pCRceZA3chXxhVFj9HetrIN+SvdU2PyzpkIb+g5VFPCBysEXSg
/X9C2/6MoWTd6Hky+EBBaoO4bSt3MyHeOZiR1VB0AjBvMJt+7MWwUEDXYqmVas93JmbGgMgWKzGv
KIPRVsLn3+pTNIGJdHoaBC7hciI8UIeT94MVdu7B7ZzRFAE+4VCCG1HMmZ+D0twOTf77WYWPUP2b
PTGDeymiZamw+2QpfbiPVZN58ykBpNltY9c6Pi/Fo7OqlbV4kFwgOPX9mLFd50CMiTe3W1EBdJWm
2fLil/2OYcRvKW3iemwTIe9BSLY8VNc7GoKCEHKBQl1oybyZCvSgh1HJH3F38Pc9zjjEp4xSz1e6
CrXyrUC+JUlTGEjPWA0LqEqmf6vXMJxjQvVeWEjBIolRVdqKYACjOkVCA9z8Ajw5rmn25tqLB/Sb
yD0xM6GFR4YN24rvvOWiVNncQJFoc6GzJ9HfdzCDSYHJC9VJmKyZ8vT0WG7WLfMI5RLzNQCZciNW
hSRncH2V6QkpqIjDpmDi7PSzz+v6E565/VlR2NtOpg5Vl4dEU7bM0QSOZv3T7/uwVTzQkV8r8PM2
ePUZoR3opYhDycqr6yUiuiKZbC5Gao633fB3LDfDPGmRZUsnRJry62BnQyIrXi9xjOI/O1d33LaR
KwyvjOVbqrwZeZXTGDpXfTbclpk339PnmlgwUYaAfvGAp4IKZaN/lvy4h/JMez3nX54TF56j9jAT
nNXWireKcccTyUMINCeXbO1AtSeisWJ5yaF5EYjA8d2xKcyZTT4WkoHzejhhLhHu8VUrhMAD0/0d
dxkIwxZnyqEhYLDjJ5AfTZ+xYoz+t3TOS5jJurpq+utjKNbgKsTgs/dFccBA/Tk/NDiFsTtybWv6
DPF7jwoJw5HvsE5LLeFhtE2tayOswSE7kRll08H/xtK8C+aIVNsehyQbe7WnZBRYM4+skYClUPCx
BHDZaBKj2Sn3ISWk1uO2zWRu+UGZl9itmNwFo1/na3ASHhdLET2sRKFp1dhMDTOC1oxtEZTcYmCJ
/dwzQFczSn9L+GyAoxRh/3VQjaw2A3y+29v0EbhMAkVcXnPBkQK3ydIzbu0NUdnmNfrVrk6uY60v
bzeNxNZwRXFB5A2/tK8ZWA9HwIsKBABWNUkJw/dgdfRrlyFLWHBf7VsDNhk10cCGGxiC8SXDIq/s
604eNTmnrUILynpTd++gsq6oLRtwr1XNZT6ueNiihcX5FoSBbHsSwvG8DEHd3FdVIq+Ec9o8zAOX
BLrt5RayDOy9nConvz01hNYSQ+dh5uk/rPC+62eQvLUFB8Qm6eZaa/CC2WILuxDGZiNiTyLbYitu
WbUtdP9PVbyuGKae8UjnW8R9xQWG6K4krzXbhABLfNL13YFUmZF06Oz2MzvUnjmABIWYKZp2wM+0
23I3HIB6di50lraOZ5CVYt3OCgPLUBuRJfmY8zhf0pcsQ1drcRkkGn6fOY9v1j7h0VJmrQdLC04j
q46EQciEHRRCVF3PecbO2Bx6M7HB28gmGBa0jqyXJrkZGgQmERtMnK44Nc2KcJyuKnW0YGb/PbIE
jjH28Z0KfWOqxrUgeo+LuvWQWstH6mmt/H0rxPnRd2cFsTmU6gfLcxyohpWBWcwOpbFLTWRk8Ntm
SoP/CR+1MrkCGTSdqoB3OMKxZufk7DJiApW+HIFEQC4GEpnt1HUbmCq4+kluubeUOR37JQ1GpycT
nB85ILqydpZrnTqxWY5zT4R1TsInxm+JsduVdq7iqQa+1nBkZmk7cfJJAPmhMzIq5aFZ9QJZxi2L
FJ13JM057nJVjfnZZLry5K2yO2lSr2RSdVPVTib9+TTlnj+lSCXZEyj3HYkp+EgvGJZte+1NvlBi
rYHzWxxshLnzSc33x3q+9JsIwFivZ5JqWrUUSF8tTXY6gIma9jgvOkELxFBb4yKTzSylTo5ADLMV
bq0RP057ywKoKHW0m6lHLXa4cqgNH2Sf/gSIWbfLchl/BFhACgEOlORkKzpinyMiuLtjde8clAhz
beAJ174VIobZfPfIdZYbPIBi/6brD3J7hB792osUuOWfgjIpohW9cn74kCn8OyegAgDy9p+Myg6B
56BExO3gzNfGGxCPPW3TpJUpVeYUgDKQ/1LmoDcA4EdIu/uzueulUcK+cat7aLJzdkSnScjFRO83
7takKKJVXwHnwhmFvXd2WMevMLyG4ybskTun3vPc4VsJ+/Iids3M5BR5K6QY8l/Qs66GPbxRYHfu
TXDAt2wVSBfT7PPkS1+b09SJZkceCYVVFsAn0E+UxCZ621Xg0wHBtHwPHtbqso+/S30vYpVaa1CI
SNvy+RLpVcw6+NbRFZeAkPTYCYoSM6qGNhoq1RUss7LRzwDVNAHPzaQ6YPjjdhtJP39pNMpgXvuC
UD3W0iHxP70r/B+BN0K7rNZ0WxrCBI56JZE6ivrnj60ToI4Rch8QKw5/cq2hTOlBY+2zm4DybjIW
KuSTqBZrhysdyLvGBKhxjQXGaCHh6Ahqe99+8m+1w69pNB0ka/XoMvBCgP8RrVMpgo9+URVt1FjA
l/HslJ2rkqLW8QQyYMX8jprBBfjinWqHE/au/qO9HPv2UAL2h/Fs75hr08Uvv+Bnph6J80PnGSU0
HrW36i+HJyIf7HwOi390MGODaCfhLYdMsEO2EYKj27SqvQvEfJHuPu79f/pRN6TdhZlSL5pgmq5K
kEE2+2Nl5z1tVI+aKDJ8M3nD5AFzzu+pxdI2INgXpEKlB1HkatEPkXQtskE6lvDw+nZrbCaNDJ31
kmGGuXewdxgMdgKFPHo6rcVgXJaOU45pBdffzordgjR1E8CprcIPysAo2etbtLfZwVKgDFeI6d9x
VFK47mLDz7N2T7wEE0jbqiN3azmwqS4ZJe+hza4LOOzrAoSlTFobIG1Ltnag60qpY/A2nVUpFD3R
x0SLDKIEbEVn1yB1dkDuyNmjDdoNvDBCMqOor4hUqT5WPwi0pUK3ceBXTMyld2G+uaWtn3bzKGAT
BSkUYcAyNIMLRdyLmlLbgvzK47JFaePxXd42a48Nx/LHGR96vgtXUJPrtS2nooNlSHcIoLbQ+T52
+PA+4JUj0F1EgWcGV56USgMKOD1kJVrUICxazecqJuSXwhGAEseBJ0yuZGO4GD8+68wnZuOXWna8
ojbU2SNRGysd0vLdLircv+49h4zgYfUDWx6OI8ywCdrAtuK69pjhuzEO4q16Xn3U+k59Tj4J1OGp
vAM2eTk0uvzcyzlaqpKh8j+bC8VyZHB3FuQCn96Mxl/5Y+9tpL+SDCLhTkeipL/I3XNL+c1YpEX4
MbtynssW0r+hNwXB+vGpcTlw0YbDM82abrDCT8TZmOKsE5pI+hpTaEh6D+qMfp+kLdpWZa3ou1Qe
MFBcbBdTBMcoVMTDfqOubjUgVTHLtdwI+VdQ74FyyVmRxEbQWPMhBJEWyJqSq76FXRbm3ZwTG2S3
Frnt5l+g7YRuQ09Dimpa3/N4ji/AVUHcjcc85OsdP4AE5duH0xExyTJc2KFTWNGy3QYPbIZDCdjj
UPPO2hRz3lCGbso2Sp7Iu48iAqAfdKWHd7LRCtnrwz2CIA0+UfOGN/MFW5tKZL5wn6CWjseSrNAl
cgvfsS6ADIvdnkZvt++32N4lbx3J/vINY4PJ6jNwa2LyF5f239N6JOmxNOVxnONJlpECW4TtoKhS
h8BwvbjwXTXuI2iomdD3qb+Qo0ijnUvPhdS0uvjgevX3eYRr9VgMMDJh9eY9sW35LPQLsDGnGoAZ
AR4GEkuGUuy9ezEftJA3s9B+egS7x2aIhWIKPpGRS1XUIzTLJ4MhJEpNJZjJFzHO29uH/7d0q4hF
uLWBdoYSfN0uuY+3J/wU2cikjM1QYi32Ucj/OnepXBwLBw3G+FANjPqWZxsp66tidkZR/ZoQ9ji1
n4fjBlDT+aH98OIZvYDKT2BWKFMYrvnE3Xm/CWLk/sV9fFOi4SpBrpWwJP9SBsb83F73pzViFQhu
PiFneqg56yX04CqGqp1IDHaAF/im1PwUstIkECSaX1cmYwWi3+rU1jGugYbFKY7eicaUZD50vUMh
pS+lTqpHfGwwI8tOsWBiFYFMCJ53+xI9h1/Zn2QZ1dWuv5Ry2ap8LJBXrrdujZzUUtqa2fhCComC
6gkRhLUrMChvz8i4giTf7WrJpPv6yqbkBaB7t/V+CfSa/BXWKjILUKCM22uf7rX0y5Ktbkgr0Ah/
5kSpi7Pu1E7prVDeOCoFTdUs8NBMdIYIF94fokXMs86kOqAgt0mZsbESIgVh6I4w2hUMz2kieiPg
Lc0Czx8fM7BtVfOID0jTFlfB4/gfeF6It3GggchfNRS/assI3Hj70d/O3q6kHPfzZJ+FnLo9yOyK
WtjS0w8jQA1f5pYECQrKv8CgnhE0Fj9pW4UmlbNjxgl4PSM4M4K+0isniow1w2Tbc9nFV8/KaZX7
2XgLDomojGOiCk1gY7yADa6FDblGkgUCzFFL3jDcMOzheNM4f4usu/SbyONL0byJpQ1DEBwKGKOJ
S42ZaLDxk3DY2ox3A3MaqjgX8139NljHMA6Dq++cEq8+lWo9WouQ5ll+MM0itqVzkbj1JyGTOZoC
TkGCxy4k9KL+UVdQhsw7+MxKP8CQ+Dw1/rMDlpxWbvZ3H1dlXWbNa15nb3lJuoO2uSL5bppiiXL7
QCnq9n4oSs4esL6Jyw/Q05Ai3ev7V4JiiYf56YZq2cFZXNiLxVqNCeJ/zEfVoWyLzzJ9mtB5986S
451yyjJgjTv4zAiBgbar8dDlcOqq2rmzj/C3bfRdiqm+hkP6eDSCp4YBXJlBE6Ms7mvJk2zqaRj/
mTl8qjxN6vEuEskRDSSP+x6hanrcDplchljejYyucIzUZHTY2hXCFRUA4Fgds/8R+uqqhTYLWtHR
HGKo493pw9ec9ivTiv29K9Hj2jo/JzlU3gUnhcbakcCNN1Mq7THo0pnqbzRdFU01XakgM1lsJj3+
6Q5EzxbPVIndgOoadV/HkM5Mafb/18lsRtjnIqYyRlh358fOcrBW7a30aAuf8tCEQGfDDDPuyrej
l2DKOIwoSN8Qsolinp4VwC+9vwNub2zosK1UZfj/6CiQI2YqOtNpv0glBNybW5NJgI8EReunzd7U
1F06KDufQQiphEs5eZNnFltlKRRrt7qZSwZ6SGZWIpzJ4dJ9k4CKFheZUa+rNgu0mKF+pKAX9Qix
TfJPR0H+6oA4RNP+2HZby1lCv7XPYNLtdbiv0zmO4/DeIuur/YUlvsHM6MQSIvEyM6FjFWm5QyFU
dChXS7dvdPYWD0qSTmxML9gAHhdf1purwNUqWlvqjIuJ7z2YPQ9Q5Re4CFiFtZldcIjh1+iBrdP2
Sfgwt/3Yq04VaflLMzjLzOB1/TfY1Awa+a8PGzN062IuliiCJvKbxcEOOu9/Wj49OkW9mY3DbyrV
oppHUMclVOpVmZh1JV8twUeJ5Ee1BrrQ7tKYbbvf1jC1BzFCaykDJZLPpR9kpb8g9Z1kzACwdyB1
Yx3z+2zAr52fxSlD9codMOEt25+RcoU+MgBz90zA51WnHUsLP0nlvwfvxSjkqPjQKZran2+oPckJ
RVwb+aFo1b2iMk7RWQuFwU8/jUUH0tSkYLrrGwf73XIOJ8j6PmzMYkSdXzkTmsxoOr3wDPSFJX16
c8Y9LpJmwJlEEswpe4w0MftawuHpotAcyUCYqcy1BdedgclQq7C6mL1WGtvDT7F79c1iLZAFq8xT
6oyqvyLRck1tlj23NzsdTU+4I7gfzwmD/z6aD/BncswXVLrRyGHFJujl/DphDmm8Nmd8BQlZwTMv
lQLv5hSTYdEuneYuJWeM6nQl8Dmtc8RrdVzX8aq8TbQkLp2EuLLB6KeaAYxRidq4pdgujlM9FtLc
hztKFAcIDHYVoTRWaaHVrYSCX6y9NBDDyQs9KcoRl7DylpoAItNET5xzer8A4jKW1t5EtjoAw4x2
eFH+5oZ4okdLJ1dCWLBEbuTifmUHdjQpydJfQcRfzxCm5Lr0WgF7iiUd4UhsJqZ6m0oz6c3KB5L8
XBUYnUIl8JXc54hoMqbkWfwW9wdivDlnEc2wIfXoIDHfgHcqmxrCQ1HuJmtxEnbR9C89Mv4gGWx2
v38YkCorPGLq+LxakdM03NkDLBnNNmIB2qGKNrm6cohvR7k+7uhjdf3QTj+359zw3+Ad6oU3iBP/
TGBZ++/wc+ozrxf/3d2lqHOqtiuP54iosB83UwnLyXmnmKWONNkk9AiHOV7CNlVIH0XpS1IR/sL0
/GA2W61s/tVsGO83rq0D8NuvCCMi5Zw7Po2wneX9vIuQIVzYNVAufpnkyBY974GuS5G29lqWauCx
xD3rRjrF0t4LTl/87g/bwfUopAbMI7/YAfgiRXC0IZGrgOg7V/VFXNX6HWPH8fUJ867ls9KkLwjV
Ph3gVjTWF+NAOyVMYao7Ue0TfMrBpkmnJz6c9oRzh1lJufHGJbFZRfvABsKKFdZcPIJzxhwHU7OP
cmIiNqQ2VICo0JssRmsy71FfpAxSYildcwJlP6qLp1N7YyQHFiZn1TnRz3b7+gQoyrRRIaFvHIcq
ohhJ/ebDOHisb+WpQm/FN0nv4QKojqjQfFRdqcIq5nBhhi4mQZ3QGgkHK+IhhsYebzbsJIVt86+7
cgc3LCciUsXuNlAn/D58gKAe7H4ivHKsejL8V/M48QJ0b02cKESO5bzwI2QqyNp0pe9SXeFzlETL
FlSyktHq4aeafM52bK9UuDOYoJZhsPUqYi7blYzsUFbvGni3yCcSlJvzQjOnJ4vgFIslqT85iobn
Bm7U5ALLsNv2dpURXrQPwVI2PVFzGyx4FDBVua2y7vr/dJIgfeRV77V3fxF6Z0/z9wqmlbjWMD0D
fmWEWmIZUDYqWmpW6qJbXYYqTV5+Uvc7CyaD4iOdqd8sOg+2GVGK6rVaDvULIFBlgZUNH0PvPxUB
kdaq197NVZ+duY7y9wN6p0awSyIhlSjXrdpfo/dMTMnYrxnh0VUeNTBDNaOurUF28b7YoHnriSlw
32Twfrr7nVWj5mAE0OL8wW9oXdxrGGXNNpB66kfIeOf8bARqQ1kl9n7apPps76q+21L9BgmDXSCz
lCulPZSo3kotGxOjCoUwRNkOBNUKEKV2nh5WpE/DE+7CtaDkOBFo+6hH/1zRUGeaKkEiymFX42ah
LQT3zcHOwUHUss23+sDeE3kTOz0fiyerKJtlzHziw0vTDT7KocJl4CQDowG/qD8SRLnCAOiWLEwe
Daaa8mj6kuAuikyrrtIXHugPKw5sVEzbgrCa4kMEQRtvXZnApXq1yveU31i2KOgGFiaTg4BTdbnT
NTL3bqyxpONG/n4Py9Nf1gvObGsdzy0UUvUZMdtwDa780h/NrLypF3o4IkwnMBhpqLwQLpmtNYC8
u7pSUumEH4/JWf3IKBbyiEV39AKzzsprrZEqiGOOU4LS1VuM2u6mff1MZ4FRjUdh2D8C+4cjLT+7
iYC50pON+Nkgn0L4sUJr07cF89uhEWy0Wvx9VcKcJwhNV973kLOfT5dATuhMGGSJ00PwPcvdRmq7
TLn0JvUg0s4UCcsZ7Udq+vNcQwYn/xgboxBJ579sV6eHc1wpMNjIIBtIWPjI0X4ABwJneb/7Z6QC
xdr/BmDid5cOUPazyU0XSKEuucysyQUGIbf14OKipRGcmIerKW2kUO3FWFUj4K4+qyEB1RTrrf7V
FNbXHcQvgz6ogtFtMhqzZLF7RqFmEFkFxD2uqLePTHazrvdlWC4Bn19HBQsbp0he/Cm/mKLtdp+I
ISt6pKwNnnNhz6Cbm0oekQBcQLS4ZZjqzXbphRRHefMRUzLCrMs7+nPAwu55Mc53pTouUL/Up+xC
+pr9M6qBK3V326irJhkxgbLslHX+lz+tYhwEQP73t3w952syHITBWiLREQ4eoNUztPWw92xYHi86
DJVBOQTx7gcSgO3cCmikLY0bUt9wMfLdvq3m65WrpJzTiq84IqLH8x/IJuesYpDjVhE0VdZ9uTgy
D1FHsFyCdINSWLfP8DtTi1C6YCkwECBNcb0F2HKpmicnh8UCqFqrTfrhRDGT4oO6lRmA5yphTy8/
xNE13OwR7ZS4oR8qLQjmRokRffWaZA+uLp8AQhdKJ+MHbTEasqX+rmFPrkhIhYjJAnojsxdA2vuv
RJfeUG0P6GypTqzmKB20EsPCCVTxGuwh/Q9YXcPDw0vKOdJj6jX3xu81BQ/l9rI8ceoS3p+FBTji
EYhy78FNGSICluXcSJV+rNvF1rbr1QStdRplI9/uGEv7aXPGkJmB+wXQttnjnkn0ISi0KSKGUK/x
XA3sUKkEy5cXDEWQ6scLNaBfT8fx4VZvGlDvte93+IHtd1+n7JuiPnzJGgzf0vTBjCROklceckif
H+TrPWCFJ+pkp2bp93ERXKYA2uEkBRFFDXsHjUkM9/V8Vc+UuVtnOhnCLDWpRsJfxcIbGcYoy9bm
F/M1p4k82f4h3SWkf1rU3JXCIWKMwXlyH4Dm+Uo3cAHAdzoJasx0xNiozcE2RGXMoLgwR7SckMKU
qQC5aQpAIJLc0VAOrVrC1eSro/mAHx3XBLp0jaqYI0GQeKEMLn2H+cXg69qHBh9jnlCFPe+iYfh+
7zTmz6/1B41iNRYZE7Hq+4e3xjEPJJAk5RgiNS0VprsgK7urrJmvLHJcsESwkNdCl5O6ljsv6/g7
lR8q7WoRVjPMzt/Jr0rEUkThJQjbXkpgIMxov6syuZRq88Vdtui8+Ic4+P4EOuYcEen3oTrbqBl1
E9iggbtOhtw6MYR1esXLyKpGx21rknBkX+FIKtwv1b5cltHjnH219T4d72Xbm6EBOMmo92vXwjC4
7550xNrSVtrCHdY5mCLES60svzM6fqBVUlqFRSUS1e5okeTstcUiOVhYkOcaUmggmIVj4QttvvxT
crXQv+3+FDZj3HQchEIlBNnUgT4verW7ThT6WP5SbH8pyLQv3bhOx3ClGqvVB7gcFZlGgESirDPF
F5e/WMWi/bVDOFIStcX8ySS/EIW8VznvpwQD8U825yU0QBtBDUrYbYKtY+IBw2lu2U8HpLSogp0D
tV7LZEXn0nwn0pIHC6wCWv4VY3oxoKuuD6oniYDxpK2bZdxPE1MB5w6dJSEeq+W3C8GIlzYF+ZwP
72tRAoGvSQU5mT3jA1w8/7zC+0+sw1Hc23KMXlBBv7PI4hURmxBIiT8E1i6jQeFoEaCoIRnim6W7
ohgeuQbF+M1YCVqw40CoFt6JZKT7LHUa0q0AHJlgSRwiLT1hm+egGWo1ClFjDhrPanLTD9kcVhtK
S8P+uhhSlwWlgkeO9wlrdyNpFRIAK2dY7/lyJjjQD9zlrw1Iw4DqHdcTLArVS8//d6gZsu+9PKWX
JVpE3b7kJpfSFTlDgh08ettUg+dCYDj9wis8FEkXl1nMHNIlGit6t7lUqxr2Ur8K/9FEqhD6WpKi
PjUs8iBVCOCrdvGWE7ecvuXrNuIWCH9qG6K+HnVfy7VUn8haZxg8txY6gu7M+s0NwCY6kNecc7/o
yjz9A8vf5cjIeNS45SYqO7rkHBoH/Ua38BaiAPTu3Mu/2TLwIGHExM0FBRAwzAfbcY/hxPqKXXhx
s+dGCZBHvEMpuIL4u/Uhkd3x0xeFPD5vbAa+s05vlLJSa5JVTS7HhysQcwyoSZvXYp6SXrdJX4s9
gzdlY9kG5D1EX/B4O0JuOGoqTP62Dn3LibI/7faqd08BchDZ82/HhsLlFsxe1gZM3rmnL4DvWos9
4QDUnEqUuD7uClpEOTjk/03zsH/p3uotWJNrTYTZgJ5TxgojMwqiYezAZsr9nsh4ffnq+quG2Ofs
uejyZF2Tlrz201cFzwhELld6y2JRwjm5NdWUYhVKeqmSCf7DFSE31CK76dDtFTdyqQ55QdlqW7Of
dDSJQWD5jlaIzBe5G5iOUYGZzmyz5MAtIs56upKjCK55owCFBFO4s7hTzbD8s5sjp8NeVXJ78YU3
kXYsEZSMpVQ2q0XZLpBK4kxoDZrXAzFHCyyqAnRy7yh4xa8d2a9462/0jmgGmVijMKC/CzYkBeRe
RpHxomBf9Jfo68vLPyvDZmzAnSeP4ToyBNVydxrp8Br7cQSRBFo61AJqg5WxvMiAcFUPUIkH70lE
6pht8/73eJnNrj07s+0L9zTmM7kzHkAnk9FIdTME16K25mebFfJKXj03Oxa/vnwe0OcyAFfCXxrg
ivL8gu/H89pevR7zVPxp76NIN/uiRXdb9KDmIEAcc+5ZzH+ZroY/syIstTsm/Fu16GnlSxjVUssZ
BBiLzbecDx2bv2y8TVMJr2HmQ9w/U0ucEEb9a7OmSBkouBgitWHBMA2V1thwFUJ32NHhPZH1EWs6
bGLh3ZNhlDYcwDnZTVi7YOZuHEJ2HUVVPOV//8CCkXo7EkhKugpuLeJdZK9sxaYaDmMcrEhycEfi
dOY00/z0sT/XAZ+kG6eYUEXtZOXQR0ZLDp1iEj1rTA5/pVlg7k602YN2R84DJaWTXsbyD89Z4ces
/JVqI84EXlp9BmSqm6Yy26JAK0xSH6GCbkNRaHZOipuGel4DKEGp/5ChAljtgmPgkQxy5Jy4t461
SMIenfLsaEdaUe1YKKdjk9DYIY9y2Cy+LUpcUoTf01mU1UAPsBeifT8DElOwRQ4jo5GlS1xaWJ1l
eaDOyEfyqstGu+SgFBTWFMK7s7GQx3DWeDr+Gz0OoT3JACo9uuR3zXd0/HKDtcmLlP8vx1/q5Vuv
yI6KpfPiMq/Xh5ARI0Xbeab8cm3dmN7137eeNOgIFz6ePSd6Z8W4ArGtcdIu/JCxs8ugCZZA/jJ5
v6XqLbbuw68q4zC47msrQUbF7K0CHdDtLloCvFD1wlHdXdAw6XhF8xY2atl9YPbTOwMTPwYhr9jU
vtBLUhKEn0LqjJrdl/G636LHLY/YJLwZP+j0vxKDt/NCpLi7hbStqBXfeLp8vhcVGIJDGW4VMtxm
aVFs2UlAcAWB1suDWcVWgYGVAT5zuuxoNxW5d3RuSpCm9fdpiF1yaOT3QEHjaulOqY1xdFkeKr9o
+l0HnEbX4QUNWp7ui/wCR/K7b7yz9v3C6QWpkyqxglk7USE3X2uugO4RN6LB5JYRjdiSah7JOE/X
1cuOHwb3q76f8r5BDEDnyahVWm5orN7V7o1nTAWrXjCnCgUYT1myI/ViWF3SYNLmaV6MTqM7Gn6n
RTOU/RBLNXQpC0XrBuBrUPLGNDUntsYInX1DZRKkaEkIFewW5riqIhVMhatHk6CuzE5VzFEbqfXg
s9azNRAaI1LAsF95pn0x03Lyc9HdCHTEFk/iIPzwZ6/rgaBxDh03ZxrcLG7+MEoRm7VqF7Ckz6cZ
dfVf6dRsxJuAjtdCes5cTD+n4D+SDzqt3fPH0LMqG/svEMZOfJPTZl9WFg0VihFdAUuvFn5titF/
ZonjBovVpLCTT0I98RN4/oMQPpRp/dBbXxK2TeS5yyHD5OszdEdlfujQ3jEgZ64U4oWnMGiWC0Zj
EOmP9vrPFvLddzWJ5fbg35EF967OG/kphNSGYie7Z6OtTeKjImn6HKB9BJ4CeXamtzFG2GjMH+Dg
GvFwYLHli4GU1paGq9Z0lIKMj4TRxn4pDmAnzeyJfHin0Zm5RoUEFYUgt7S92xwMEMN8h33o54ru
VEHbVFvZ9rxXLMCYZy2B4mswetnH45QzWCN0YqDrfIu0OS5Qlp9b7pYig45hdAAxAYAEPzrvXFzc
OQ113EMMkp77ZZcF5Y2IsZ7CR/cBhcD/DEY4ZFDzI6MO4gkNrUehVQ0YBfiYQ6De9AQoi05Qm+bs
1UdvygyMqFMiVxQAI2Qs0cdntPI1aJkcnmuPjrdXnibGqFxzVbXTpyPzetU1AzSqk6JRzlbfOt01
eL78JSBL1gi5bTVIHGLuYQ2AiQk4wxtcuER1TVpwe721MVwjqyZMuNmComlboo0Ocu31SedBih0y
+W1M5uZ2anCLEj0gIt8uZ883DOGz4nfjT1NFUqRVNCppQeg8xfyEqAcwYnNLmwJFh0emM/qBJ4yK
yGhecKjshhnsEeVPztJ0e1zNQJ1V3MMwhd1x7NpQkCTuv9lu76FP0hYltX04v57BgmlNF0HZ5LaM
icMONtEpEMw+nSJjKjoLhIky9N9Xk/d6RZmXOR4Rm2a/NhXuxIIb49OEfB2H2QiVdDSo5WAkAKYU
n5k/VMTyljlf0SQsd9cvzsZMTAyXXaqHJRQXWpAHRKOvOk63ytY8uguKALdmmOm2BiubVmQFOXfb
VeLnIMXqUv/ThL0mP8w9yG5kmZO66rmFtMp4VsY5zkPd/NMX0OZzemhjdfSjd3H0PepAFtkw5ml8
F8qpNedPXbnIs0SZok7nLDZvzhTuK37mO2Lg/6ThDebRtv09oEy4ByvhzMRkK9P9zxmQ3EN7YA1v
OtV2gacY4A32OldRvb4CJeCbwnt2KElKJNqgCi4ifIkqx26EkAkOjsd6QpZsx9krusaz7iJoR32m
bA3cwra9XGbjjt9gc2zovF80rwLFJsaGbU/oGZlFNW2CpySQBfpkxKNaL9sCJpkGHMiw53vl6kma
66Btj6bLED2K428meG8IJ8uZs8OBGVfDmTXlU6Gm2xHKYXTPg8iKuHrLuDQZ1+k285q5SE3OECvq
z8mQ9GTemxEEjRIVQDeh5aXvqQCAlojTNUuoOpl+sdfC4TFo6NWd3lMJWw4DMdeq2PF8bb3TmlJX
6LSY4/k/mUWt/yovTiMVmBp2M8P4Bw2Rf7fGka6V7j67lWUHMjDxud2p5PkNXCFLZSV6cjgQOgti
FZnED2LHVEfpaQGmno6rTKp/YSPLdFzU7sBr4myy4ncEtmB5HLNAJyb2ViyQYnGx+9dQmCBTNYEz
hhJDkcVzzBRGqZyo05J+URqYNpYuQBlpHTO3qZUFnf0ufp8IL9EO9sGSsaJBQPjeLq0ciJkDQ/dU
Ugsx0rGOFZ/us6U40xVYRe/jrTxYj71wbRZghSDjxlWuulwKnXOT7Yb3WPS6SBeHrdxc056gNPWD
PcD3sYog40z9Fk6WltFXqlubC+GmF+/OQR6JjsJ6aEvNOtaD65QHkNHMUwj1mXkg7YnZqeVqf9nt
lg+GgADl3tPUqvJHWPxWonUeEjlU/Tkue5abU7mZb4fJUaHkPqHBKZri4M8ss9EZYt2mUpqsI35X
oLiLiU7xPIdJ03F4IY6rZ+Vk+LpH6asZUkQ4IeiHU0gaW7lw+tDoMTkY1FQPE1WIOJmSoqXe8ny0
77ljU33NhF7oFSaCEXKlosxm5cVpiyZdiyrhyy+F21f/zwdQuYkRY/ua3m9GlntsEsO9uM5ujHnO
RHGvQSrj/qfrSwdr1caBGFm4sn2wSwHZzJHR6UVRWkrvoCDttZo8l1/ABEl6FbqZYPEBDYYOCYEx
LKdBW192vsLmxWm39D1qedT+WPljWsVtztyGMZ/0ih+LbWkJV3vscYnZhU3cqdwnLE5Kfk/tQBpg
QKLcn2ruzQEpgPRRVTa42sZCTl5bHRA9996sMjMDdPLv7o24HOfNIK3JCGcXXOkBh9BxGQi715GX
jMvhTtLjVpXh18ipz5Us3CxgKDidtvdneDQIOE9QImMz2LB5IJekbPdgweJGXv6GYsWOH91XEe/7
xWpzpAiccBf76SBo2Ph1Cb+GDai4m+6C8RE/ANynY5+PDQ2GT2FeLZvKKF5S6PngKcSmedx5BTb2
BERw2L74PCwwwR8yO6A2ATVI4fJUp6sVq69RVddmiRqBe11HacDMaWAPWR2BxL49RlfYBW0iATj0
hop1ik91YotXsOL0O/UHe4PuZHOHK1JkfPG9fAFQnEKpl3th2JLsu/NjpJyGjcug8SjoiWQWT7Zf
vNlR8a/X9iNQac9cc1auKS49+1A8W4CZC9ejg/vC/K47Y15QYARI4rcKr7eNaRsGvLp5V8RLzGmv
+w2pyGgq/XYTdq5gR6L6lVUj0A41gQ2kRr/xnjQgFCsff+LEcM4ckl3zFEsBsXmfZBp7Mg0CqLJW
YACbLvoXd1N9ZzipSJW5SI8MjXKqbYZ+STQIHne01yLmwKqc1UKI8SxOxSP0ejoMt1D0ghc2xk93
HC8MrRTGOo44u0oWK7Fy7R/uLK5ljh2H4Yr1V5dOhGOHn79nMhuZ1jOaEyxHWP2+HlryUQiX/Myz
F+cSPFloVCRNDhnGA67tj90DC9Txmc1RYcY55KAgX8SLACmvMxKBWuWyoRt2zgpK95BU41sBGGUa
D/TNylq3MDmv6HrzLZGPDbQbvPcLYgm+h554b2EyG+81bEAkXmKG5o55dtz/2/tpjWSo1Li72oZX
Ij4hZvyovX0MqkExmfw0fALusc7Tg2nA9nETP2i1mfovi0RjAHyB/g3BQNquIuu5YqairT+B1h4G
DEZIoXRBGzTgfbW5Q2itmy+X9/mAYSNjiEZBY2UnRjLfY391ZKzVAobJMor0itcFnVbYWU4itdni
rKATlOoULEMczD/ybCuS4vygOVhfeM/9yW5WdNV5CyHoqHHHATh0Bw6m6dmzTNJddCEKMg4mxTWO
MlN6RLjoJZSIHa2TX7gBL6Qo1flKoZ4VxLMRaDEaQGaPBVkNVXAu6ENQsjOfhHz70tcsrPUBzgPV
P35VQY6/8YqV+DKgJZjzWi+gx+ORLqBRw6GCifXZGScexkkwZF5msxhCQHW/arQ1iCzYyyEd6l8S
yqiN6BJh8fkedzr2EhKLqvGs/+HguhveMjk2WKyRIZv5RFKzw3SD6nEQDXDjn7RPPbvdnZN7vumJ
sZMowZXm25YhiptjxkhEaWgRGHI1BsmrxAumZ4TPW1JmWCD8vnaeilu1pR2F4gI1y3APItrdaPO7
IQWDrAR6yHZ+pMd1SGHp79FCR8XFueUEX7jvPQGR310S/AXR36d6opTEuW/hbkyUW3HetiTcySeu
omtfXIlGm5CkrHXhgsFdROdMQjUj1t2kzVM+ELaHJ5o8AOJkQrGIzoMcwik2ONrFM5GNRvF/BHgB
kxiSuJ56V+VvRJ8WPCOFdtiSe+KhVz9P6BSxkf7YRJsC+ns/N46eRSZdv/aZJwd2KRRYea69XYaK
jw748z1Q5nHhJ6I6C5Oph3KfYltvzGEp7baJjhrlJInPbagcMndPkgZuMuZdGoz0Nsm+cWhGrMTg
QY4SFTV1BvcLK2pd02nHU38msIqh30NPEqjqaMFxxBSQAy4rxeAZwhavB/hBZqKs023TW6Cji0Pm
iRukHiCSlbH473bkSHb1c1kLN5OqEMRpbBVsrAIrEveJXIXGWB6b+PmJcwYdLzjniKDz8W5LqeeV
sXVuuoKuJNpZtZWTpS3Oe2FZyvsDFxdO7Kz8HULtPvvx4HkpAu1Yrb3kG6OEiExYDA3GuGeAOqFL
075OTQULTqa22WbQVuSRGmsYH2BVCCYkqNNvF8qAdu7pt/5BjSRBCticH+Y2Dc4MNN1XRhq/aKEh
8rQ1r79a7KExkjszt0RC1SnBRS6BjnQtfwiLSPc15v7voxvzMXF/ZzR6zOzofqiwZELMUEWIDzpY
kOHCXM9kQDDmzk04o41CepzNXRa+/TV0jd3yfJLqN++FDILbDztKVygez9Oz55wxG2mITE2jZyDH
2uGyp+4dbjYp31AWXCAvew5Q+g3r2b1NWiq5hGqINAaRMB9+KxsfGA1OyiDLppjvw5QG1WjgkgDz
Af/b1bX9rmqw/zyAgyf6M+lrogaU9oSsaQZYS6JgxaIQ8K3JkSoHFCcj8hnwhOskvIPwHY4huC3O
lN1BgooOJipmCzL0OxrCc8RF4Wp+nCKSP+o74qvSUXhVZcmAACqWyzg72bJD73CaHUH7qUoauFP5
OG5JYudcgxF672z15MQXk06nJMZF3IHmFU1FtfolFfoG5W4VCSdITC4WXxmeQHN+BoPdum1LPukY
JIRcAGNV9/VY7Qg6nmKMOrdhGHzCcq2vFs6ex9POHSwbSHlP7LTLtsqs+dM7KYtor8H435DrFfKf
9T3mC8dksHBuawzpaGJHEZ8/ZpzDs19YC8y7m2EmB4LFB6dCCdAVuSC8Sacf/7nGXjYKA560BUYB
5pp5b412+A0IJ5g+JnuhkHIavy+gOt+X4VCNt7sZk7UqkFkHXvuMrL2cZ+rED9KaW6+BHwP00e+3
kjWhMlnhS2aWqeiEoOUiwa/YRsc64vR87olQywb0NYjyAY8lUG/sT7wdXfIraDX7mX7/JShoBdx8
vzy4WGe5M68U5QguR0/8epUsZeN1EqSW+kP3A1q1Y/IySL4wBqXlFyX16Sae6O6oc9byLzoiXHGM
FjCrQsAHzhYlswzHTnSAMQ3ketjUn0zqeOdZ6AgV0s9FIqeV0xawKhbx2gkEpWWYPn5jvVmHaSBJ
DTplbe3VppLH+XBLUIUA28mSzRWGCZ0zPy98qQg0vPAcBT33LCSbe0AKyf3Q96bSWDCWhLQI/TyQ
Un8OlT9Ju849IZX9cxwnw1OjVys2VugG2l/lYajklXQsfBbSOmUi/jjcImAV8mxpu/An6INUd101
LTiTphYRYZwibUsZE6yF2e/7XDLw21LV1czIxcFpJ+/4SLII7id9EPWGKixiuZCrMaCwe2uwyjrt
boiwzAUFDR2XIsnza7hW0otHm73obzyCr/YEtHt6PUSuKjzAVTBNyHll1WyHFvLDXLc9CUFssFuk
jwHUTGBDGjbaVNpQLejdHuHrf6bx9JWAEdOtjcVdNrTfgEuTxYXEE4MbDCvR7J3a6LpH69+e+KD0
VrBnDuWWXAb6b1m+ePylak/4fNTdo+x+2vwOcA1XoJlKJOfmZPXk1ykFREn5jA1SgtXbxoLf+9ee
1dJxZrYheoDbNekdNjn1olfmbO49ueq3FAT06HmMyPxslSpoffGN6AWmI2fjk2VEwdeUON+6PdGx
xQevaYBSn7CMmPGffARHs2lWCUi0n0LpsMUAx1iamqCWZS178aUv78U1A5htxFcYpx6LxT8l+QIB
bViBHR1hLK3YopSjErj/sbNtteVIAi7LfRTlHzqne5BdODFhUUZ74nF5lr8rdQK0+iUjcJ6UJgMq
zBiBfrR/4KUy2wGzQHb5HhlxjvVjHEi4XXxSN3b6L/LrWomPDCu6OlnBpb3MFhS24UxnlgsiBt68
diLPIb/Vu77WkytQM4RjRFwrtfyNApo4P6KCwezKEeTTbPPkV1v+npNUwjDifv4+SyOWRAifJuBq
2e6pjuoqbwI18UUFT3vjLCE11eEAoEB8S96hGd+HISr9dBMQNHY4iSJ95qc5AwkP44vpSvMsghG4
h2F7JAsAn/2/RoarGGFEjcPsMwqM3cgSc8Ukpc9hQWYnOj2Sd00lUAbRl8hz4lw4cz7okP00b18K
wigLmWgA+X6MK9Gm8ciFomfQI/OnaIMORXBliY3rxRzuEFYH7DG4DeVY47iZQLJlzpOHivrkrVOY
wI8XdjqCCxiGv6ZMFsxIhd9guHESrz756QKTH2g8EEnMD3JhTIyEyfRRBxJnG7pYDMZJBWUyn1+U
VSkWtAIv/ncd2E2v/06dQeTFyWkPYTz1vN5BPI3+MrFjVR/KtYFXF84VUk3jMjTLy6Ku9EXUj177
VCwEbJru1iFhSLhKFLCeOaf/uYIIfDJh0swx5yjfEBJRDv5PF8V5/3rg3B94ijv7OxsPqDShNCEX
DPmRyqUKdeWPA25jIBtUJHo+y3ZAvVfTAFc/dZDs9S4RjKujZWNWRaXZLYV4uXJyuAdGa8lPX46C
crQjCYK3mhEoepB9qLyJPE0hhnwb2biV2re7D7UcMNRZyAszWS0nYlTtjyp7xZHf8YQluuxeAYeP
ar/OddNtHzouxdG5uNRnPGlP5Y1QVLW77sZOuo0jsNhQ5OExDN9DEGmfDAUCH9fhyMxNu6czUCK2
gBnQF4ZK9B/AFEoADw0swxKY4pjCq/EhqoIl8+zqrDn85szlgAK8MUtbeaXHdx49oD6L2WKdMw/d
xKgwh1i1GHCt4mS6yZDUgCNyIworIGHGQeiFxF5uunkw6nFGVpmmc2GEC4Z3f96LD49SNb9Xca8s
tBjZRd6ho0DtOrsIeLsynkq6cXoh7b9O//J596gb9c3PldeC3MNgQyz/1nY5BDpM248nyrJNhyiW
oZQRA/w8omTphiU3LG2xu2uXBCW+TxGI/qgGDHtT1zfmLwFMGQSQGFQLi5D8bGx00MXgsann3LK3
ubC8E9STyUUGBhoEn2OETadlmXvi1fOuIZvR4dhxfn1KE1g/EwNVfNzf5VjWaLCxGnZR3663Zrmp
wGshAi/+pGiZzJALNkEKsAL6x77MXRy5g2nfbacOgwd633wg0ALjtz2c5lizc3Vz5KuAeOlpDRF0
h5yAJqzMhOjNxzzAgt4R3hywueTRGiegbmPcKnwMPTj5BEkUUq5oP0rxqjVKn3UHfnJ9k14ogpGM
FXjn3kR6980SpVqrkGKCcfXz8T+l6/zmUQsWEpQy3c5TQZWKznVPBGPAuFeDYvaREhgz3Wl0q+xQ
HsBFDIGdg/GodjKrgbhbzRCwD62K49aql585Hw70/K8B86Du66XCWoNAmNTdyYNj9PIQEXfhUnUp
yPjf7NftVfImEvvACr+p8gvtJ8p4OwhorVxsuyFzaLjIewjYHyo6qw9dTvHcYcYwIeehUJrgvgJq
LvARWdpmrQ72gyihQ17GYe58riUzTfgAOgTYok4DzsInrwJqjZNmuEkCUIECeO2a9UnEoE5YTR+J
J5VGnahCi7bmtw+eByXY/xsLvGYzzDFtmKIumEHqX+eJPX9tcR6rVgrMHOPwazwAq8leuL8GXCmZ
zjYzJi9J9o17PpBblwOxvCyZFuilcAArULFgduIodGglcm6Hc4TS27vJvQWbXwPZn2G7RNvIuWDF
LV5X+54J6PD4aLYJF/2QdSbQKIgzvA5mbMye0dMUbL+Iod4r/sg3ydiHsbmpS8NfQ9aNfQPpUSeL
sFQxfg9a6jpN5nC3FqVF0SCU9BLSV6P3NCalaDcDyT5K06HYQuH5UmaSgf1oaPGNsLPa6PduVgD1
4d8Ice3Qc9dSCBNyUCHNpOIcls1prn+/cvFxr4+eR3DtQfe43siBLRSPtYcPKeFVyh7GMOaa0/zD
cJ2uieytUezya9jG0fSnyToeZv8rMlOmrGMaViF+tMAd3v+D/ERYvSEC6xJOUPcc/9x2ayWGu1/h
4sr32OnBI6IAloNoc4ertEe1Pk7XMCYz+/ztykRKfkEgPaHlvUo5PAhSdxMmCTR2PxarrBmclbka
WowvzORDVet8bxb/un+XUHcCgY866lSPdlvSkltAgwFFevi+9ZwxVTxlL6/hQnz231FWa4S6PIhZ
7SSs+9u3m/Lo9mbHZjKv8vywkzgA487BcgPshktATdHlemrkXNDXw4aBObLRThfQzlXSW3DehxWr
Zwqs7VG47qkyvF+k+fNW5eiS0TH/usc1fyqS7MP3dHJpEjf5LoL5P5e1Kra4gDAFL4HTqnzH6Nd5
zes/XGB5wIT2rftifwDUNt8A4BPI6bSeHoGZiW5x0RIM8fSqlfmbRDP0/Z+zi1Sqy/NVjiOnreAq
NGvAuUT++zpk4LDVvFW/ngKda2kRvHL/mWS4IOhIgt7/KwzO3SJ1DaYBcb0evW1pn/c7gA7p6ujn
XmSQdYb/NRbiz0jQGjZKqWMFD3GHcwZLvBSPNcZTidAm5C+XpXM7HTF8xKkMZD4XqcMS8u8pVVRr
w4loLTKKOisa81ppO2Ge1oc01n2o5aV3mCTf6kIpII8uWlF6IXg8ImcNBwylAgMqPmnOGsB5aSdg
nprslTcOHpKWxpzf1iC3fXWe2yAllph559vvALR8tpRGWgn2wl7CSqO+4pJYE1p21kBNWhcXVkvi
uDNUhvdNhiyMjYHPhHn1KA+LWNarMlT/fVXGvvePfh5/rUqP5+GYVIxTtZX8P+PQ9E4odtMdTH1S
E/M59QxWtUMawTPkl9PXZznwBLXbaLZzajMiMq8XYXBxDPzX3bFlfI5QNHS6tHzcD/1VGK4cjQvW
Ho0T1/ncM8zS4uuFpByNbg0NiZGCt66LpgeuXaYzLqxUYT4vAeDkyKJkXZg7EuyacC1OK7DD67p7
LHjq1KMOoUXT8omXkVLVu2KE0Az9aFV/cQghCcpeC4tYqWB0GckgpaL5M4cfeErTwuu9i2IkBFqo
GMNGwPx6S5u/fxzurJNFlhO6RquiiC0GGFhu2lDcgd24FNyAzzTGNxsd80mpCp/46D6ixbc8AgSY
GyK2c9iGOpOfYa9XZq5rYeWc9v+l4xpb4qt+4Mp35/RM3Ko/7MMZz0f2pPJqyCyshN1ukzlO+uRr
0ZTeZkehkN+TRvesk6pjw1dTu5kLEDQN/WtKF0zpX8fQtycSk5ROs5tKDEDoK8/BTVo0uF/mhbWx
U03n2I47iu9GF3oihRt5aaMy9RC1nwKS+kVfZSnaSh6sMaPP28RZ107XLaEDFyDa+dUU6Uxy8gU/
3qhGEKG82Teb4wD6banNPXLEdMwnr8buvvdZHlSMMHLXrGYnIvM7PJT4cXiJRqoAr4g06KFQQ5se
EE7LMiPyzazDe39Go7QxwtU7eAJZ1nY4NoMImGr47ec0Z+ovYJHoUZdt6DUiJeP24TqlY8UnH1zj
QLnIN2drie0531cRzEO4XdauVGNxcS+LZiMq5SzR8j3vpeQ8tcwMgKv69NLX1oOCrT/+lEYy90VX
v0Yw2SrWWasLhHJclu4GCfHhVcb2reVeXvbVWMjzERmVkL0Intp2kOpfXrCuMGiJG45l6SXBYm2m
eZ5UcGhoGkpws6iLb2w8WDqTaUrCEZPhVCdMj0O+tngAm+prwTksmVd9mLcwSN7RQkjtV58aiu64
iUWcsKPBbHWnQb78BdbSCplQTMYZ/JXVxoZcxUssyLQ3N8JWwYALwzvDYnQpnG/eo3bgkr0KSP5c
RV9GP3exqgk5SEtTVG8zRx+vCESu4pyTaaRzOEgN1DfdOLEdQFkUIrcEAVqALrGbsr+FOzDZj8f0
GgQII2UZ0aUHtGXT9hy43NggLDzWuXKTUERe1hL+mtWcmQ7HSClGk1J4W+A4lod7OC0ri7TeMUxP
iULY5WHgNo/Rzfizz+CYJa0c12XWe445veqX/KMb3Y5UxqR2dk+iYjIUluQOXBH1m++XuGDz4KjU
1KDkFfjPrd+Cwbf1gMt0HTJKPGSE3wuIZ+hndbe27ha49r80zJPOASuzrlf8F8cYYw5aBUHvZEkP
1S7HvsZTq6FuYrK/QAKKpDjqnCQCAo/oce3eBT+lGiSH/YVdmFVA8+ivEUQqdwwmNx8+DVNovfWk
o1yqLIzhIwoDewps3MGtq83QIhP73E8zpzbFkBB5Wz/CEJNFAIfHvHOrUaZlcLVHTwe1iOzHDKyi
PUBS6FgQCyOnIYCam27vEH+zFpfbwndlDKDSE829omVqWXozewo2bUJ338GGuVqRar8s1/ySfGpg
GAot87olGa55RGJpC11rscGMAGzEB8iovdWfDyKJDWedM5e5BSs0opHV9Tkyo1HqD5bH+VaQ8Pav
Jpv/QDTBax9BQ6XJBdjSpTUDzTYC4uZLUSl7O7lusGWwpPCWsSM3HbgF6ev9Sb0UQPOEEkrXrYel
NhRUNMMJ3fmty5S1qJROadTj/26cc9MwTEA9lbF+xvtXM7Qwmmc0XJgMJ/H9isLEADtfdmkhiZ54
Embh8j4EMlu27H0dLNTlbyK2TK2GbxF68MpevUtOU02L5ufB537h0jammLcqkIuWGny30pXxe/x8
iUCDQ4d0hWWdsVAwEzcn0nCj4J/OZA8XxiKw9GfZJWfgzMPwG8B0tJsfaAkYtJZku6RHQZOyW9l3
gcFEgADhA8ojvLaZlmvaoQKg9r0koPGgi9BdU9j5MynUnrlZ+INeLwGT1R5X7ENZBK66Xgs+Wk7p
SFZIG2nZvoZf8DeDkTyGzGgcpaGXv0jXm9hAFK1MlNTQc4I7Rfkih/i6Zsj5XXT05buQAW8yABut
acHgppWNU3VhlX+mR0nBWr3lF3ufPfK3F2fq4cCa6i+5WjvbN4/AkuxsOqjHZ7BDwgUhp6kGdv7U
HUbGl9B1rLPflPBmt4gyyOX/n9XnXKIgjjixbL9tP1FkN03ukJRXSdNgflODAev1dw1AT+jWUBiy
r23YYwxKHpB8C0+W63q2oCYACEmiG0mjKLFqn3MLjXPlOqeCaRwn15E+fW0peu1Q+t+Ok/Qpk2es
/wLtQB93ye3hDVDsOVlAnnp6hafNQv+EBt8aguks8anhhga99GvrJM6aYSfIcdLL6xLpsRu1aLUA
tVPjkzwlNk/8ZjGa9CdRkRy5k2MCb0/y3FgMBoGgXg1YBT5uJlIm2z9YuTDo6OJUB0kW9/hHC6Cp
GP6ynEuB36F4MgSCocOcjHLkEDbNOerlutAxWVFdBu1J4AvelD0T3eUIr+yjQZqclrSUf10YUeD9
kgmoTyCN5Wp0YZ5P6uiphhYhKG4hurrdQcVGnsFcS3A/ulLVJ2+P8YGTesM2PjRFCP+Jx2cP3EG9
Irz7crbFKvSo01h4mH+LZ4ddv/Ew3rvOVc/7Luip97S5kIwBEm+oG2uf3fXu8Vst32RDe6D5hHvK
guujzOu8GY/LqAELQkMXoLRfTY6u91QqCt7y3fGAbpOs0oc9p531gaVLGuzdoXQjq4i1dekQgFsz
B+ZyYPzQYZHm6ujYK+lzPQkUpOm9dOHIbEOx2qmAzVgnBpmBIvuldc7v07HKoqolxYoeEXhCPO5W
ZVSi6ud6I+teVKhFNIMJRINBNAi+OVfomqykAX3/xVGrSHeCQnZ5Ys/P5S0EcCj60vh8C9i2UeJk
aybPsy5bVtR7Elyhb4TB6dJymT8lscdELe/AdET8rkTq8xd+oQJs+f5liXsS6Uw4jfWQ5kVjw+QH
/IbKQxS/qG4U3mUPQt62Kl7CzZTJ1r25IRwhLpOjPEQ+hdogQVI8TVEOxsEKJPEWEkfppTvN8tKF
uOQ5UnWWNNspa9c9UjRP/09Eg1CgaoivlAZP3rBn/Goxp0POCKriivAiqHmjMRkxJsmAG5SVHxWb
lJzgufUjcfph1/i8w52bhQEfwMOXUJwZ3yOpehmVWyi+ca853HCDQa49RD9Ezgbv+wxO88FcPuzq
41d15hg8jZTb1iorNzskLSju1rhCrw9LW5uXxreQ6CFJ+JIqNLYlmjq8KkhJsBK3amok/SB695Kd
Kr4VtJV4Bl8kKQa+vKpO+Cz9SNovE1bKWr0Gfu4R3d1nHdm9qZy8Jozz2ltoKC3zycn70pHm4pQ3
WZ3q+eG93G/EAgQegWRkU/McFoOLoHnwhBRy1Lfb12nVqaewaQw8jNZDHt59cnYM3vyonaqCgP2J
vJdr+yl3+hZ3ZXDeyaT0+T4g+CXm+/Iwtk9uqW/yeK6MfwIN/HtRqWIisVDGqEFIpwWn11UWdQkQ
74i69yYlnIJ4qnhFljNb2goEJNSashKiSimonliZWSF/IANMe7/kwf6eBL3eZaZDGb/1gXkFuQHm
1Riv112zRY0vXw7njFGfrv06zKfUh6g1uLo6pX190PUL1Wdo8sgEG/QNW0HmTliIqwFnrUAmPjXr
eQy8Cyi/W923tHCxR+rXMTKzhxCo8R3YjKZfrPc4pNS8lIju1wjTKw6NTCM3sOy6cFF4/eVWMlpT
GAgUwxaiN2Qsat3NAvN30NuMXg9gD0DoW3FBVgPcXK7gQ3D7Poyu59WSJJvqgOXOtDXqDRekCjNK
CrO0r8m0Thp5ZctKS5hh5VXTS4LIbOVnig/SVd32b2onm9UxBQkb0zb0F3S8+gs8MTQZzlGPOvni
FoJNruCiqgjja6kQ8YJnq0GLfykRSvBT+/0csxULRqkIzt4bqJYlsl645VOxh7pCJDttb+mUXkpx
Ja4NxDS8FyFurpkf55AEoN7thlpl3fsBxazW/IZ88TEhK6XZDsJ7L16qoAezBbs98NtS3BMmLC7E
1KeOhnay5VeANW4YsmoozvvgZISJlBtyhABlU/HG9uqg+bBAPBSjr/hyp2akJK/utZZDkZSMC1Oi
jOY13YCaJIAsOYHA5wtd+PlPA08MYSDKSpUCFE9tfpjWK0A3UtdUfOeWP38ttsONhEEkMsT24o5T
IZ7FAQ6MRO4W2jNDHxJxd5KH1HxokvNeZWBzP+hVZZq/xUunBcGqFNBKfaG4DcU5KM4z5YvB4+D4
uJKnKL6wtZot2NVDWcYJCjrFANqHuHlLOmdPYQQfYeko+2+ILs/yMDqQ62/OGNLa4WNvUNAJYOTO
SkOIzw1Dn1scN/x8qGzI471KbRPhym+YpN15/Y5tfQZI9Kuy86z3jtyn/aT8kdcPYezGzWOaEvs1
8aQqnPrLNGsWARtKcPqNCTNRH4y9lSkJWRVUBduiH5r26U4gGaPBRg3cjPq/Riyl3nFCIvkfhsac
4+NMFLKp62aXG6ACdoavNFh/vsA0kNFrSIFAf5xZxPpWChqapgg/p5WxOocYm49d+ugqZjSH/qBt
IZjEfe0NZkutvdtKCaQUQyTFl6ztdx/716SR71Kn8XLIXNUyMNJtWABQI9LgakGnILyrrmu+KmjI
+ZDJtJtDByKebYgZ1AfIct7neZtd5kBhwTBr8A0Z7hM8eaN4+OKF1qEas20hr8bque8poMR+vPlT
mwTliizJ6qNDvm62Eq9TIW8R1KP6+6JOYuDdbY4EBN460JSIfMt99A9fi6KY/4wQTJzkZxx2PIVR
9EZm6vsaPGxVIYX9f1uiyYTbMUEoOkuXonUeHNJUHUxUnb+YKl+uX6mhm8M+HSzD8B2TOelAoxFv
wLP19p8vJCVRpNSbtJgT7fJfJJRH5He3wmiuGzh1U+ls5HV4orcF55FofynsaiSiTDbh+CVb05hP
We7AasA+J1X2qv4IxUs2Av8wtbfmzRCga2f67OS1/kUKGQk48a73U/LYO0PPQgjbI/FmkU06Lec1
rPwpzuFaRG4Id9LnMide5Ix1cMidWOGGY2ecwG1dFKGBufplUu7OR2J28NrJP/IYywSbLOQLjFLU
a2uYmu0xRWBboaw6yHBeZfP8xP6IvWGBoEXIQYBt4nPHVbq21jZRf2XxCsO5NIhzriwSTTdQGQq+
f5NINJQvVNl7jzU9wZ4g4ZpLxVSKHCd0QB93t9KVJszXpyTbcXHFFs86tEDhwZRMeoDxXnjp5ZxV
KwZhARNaJMcsi8H7sVqHdwR+w/DE1Jcp6HP+DymXPjL5O1FvmljTLKkLhWDIGyls2AuEGnv49qg4
PMCYkDTdeQ4wOcOE1Fqkqw8JaF/fUjgW1jDV4utw9uAG/tgKsqYKQFJb6MzTWARYvUAvIZw03oHG
5e9cv4kUzbKsbsiAmxLAi149MSgt0K3r0FqewcMmKU5p3ff/KCfXWz2ZOU1p3JMdRcDioA7PtoW0
aNXR40NC81KWmfelYStyBRoLxGs/aI4QTaFYvbZVfKy1Y/EOcI8YIASfIznIfRvd2TdFkkPRoAEW
LrSlYheO9P6a34wXzAZDaFt9WMCJ6AtfDJFPMeTTTvsbidkZEl9oa2/3XV52h9nC/tEbv0RovR0a
G1JqyenOYOqvnxKevMgmbdQNYo2/ZxmgRzTImOidkf742ta3+EIs/G/WS1BOPww/VbZGu0C3CZS/
NuNoERMTgsWQlGrEdXu5NK50vXmCiP62JLT+VA4KX/qyVzHn6fIj7HOlRqjCn5gRAFEIl4JBoze3
WhQwxR5Hszw7Sbr6UxCwQfSnojvXpa8XG0blOsxMZ6Q779mDTiuoFxfWs/bfgfbhKjh7xx6f/8t4
UNyEvakGaS70CQg//9BMKxjiv8KbjNV74cftyVSdwYHXn91wQGwurU2XYGrdTuD8UrlAVEAM1Y13
HDfXFNh4feCWuSemo5dtunyN1EDTAwAmRuicXBas6dsBqPZt8njDClZ/vOryUDIQqF+zh0hiQaOG
kT4MYioJzyYGDtg2I/zZIS1vj8N5kRCzxNLNEIGbEvExsqnbsGWzD5oSVzo+1+yntpeKjPdoHyfb
OK7O2BvkMQbI/TAtgY5b+lL5pEh7G7sKexBFExYl7src8wZ2wssOoiwq9bh4xR6APdoLh6rniACi
y0E/gQP268VHNSuTfnQzgBTQZEVVOHMZGWBQmcgqhx87pHqVNtQDQYN6npJJxvty0WOniF7yTQat
zUOYzUkLoupNTH/ZcxwkmhEyhLw1YVu+wqTdvhCZ9dBmmdzbgr5iXT31iyg405aJCwatqGXaBnCl
twiC/qzn5G6BblG18qRUi1rr0/y2HLCzGITlXTFDm9pDhJQTYvid32ovHHijtnSjKxQ+OkhtHX8C
XLqsRQGvA+j0Utck+jjskQvTUiHl7DMxvoWqJAdX+KvYdNXiaipG4zVLf60B6BRcToZOmcGQt+ls
aca8eU42GkIxBo1bTw0173Ang6f+prWAz2pPHfr+WWLTfvropp/5yqfLC7q7mTffEdfP6m8Qi5tU
88OZXJIuegjHpKuHp6jXzgSquVbvZuzKHt5jyWFkH7IVrkHEkEKXjgryFFNTj/DEucp+oNQYdqeT
Yu2Cx5cMF0Afbvjdb1FrCom5JqlvwBXDk0Y1efYAufiavbmXstYrjpkWfFxEWQQqzA5EeANzvLO9
gQtAjaix9i1QSCP2kntjCnaybDEMZ99NX6u6cOaWYIkSwnH5IWyXaOjeMHc0oB/9yz2TV7WAYp2d
Ll5iFADcxK6TFM7XhmOewpWEw1p4qL77RjhMP+5ukElvfOrKdDm3YGrH7h87Gu0zm5ATckVC3T5C
Rhx+ZKDMIZDF1aP3cO9WxefGC2TOeT6Nt8MXE1IB9vKxYWlFpVeATeMgS9tb9hPFPLYmyDUtDxkV
FjCwQ6OOiLC6nGnOFw9DEYWhpshJLTtT+NI8sZNP0QvtHyjffViPJLgsNnoHoXA1wpQEuPA7JQvy
sUMgI1iNMz6LvHd2GnOHOXrbu4ewgrfFI+aSGY02Yz2i2Opv8q/ELutbH8Y6dUXHIlIlMK8EP9Rr
PoRzRyFbX75+IdZtmAVEOThJwyVaXbBjun3tdVzCZjWD/uqdUEgS2wXJip+KSmnQbvRm2vFZD4TP
rqOT20EVPhMOj4zcCL6QkKxQm8w2vUt22SdEFuuZd3amUcj5kV30xe96+JB2Acv34kPASjNXdBvh
WDsuaK4vx/wE1uHYPoTTULyO2oJOZNhda+MfienO3vE/kqUSqJlWKYMrkfEbhAOwkQfrd3/ruWCO
87nBd3/ip8VhgjO4XjvqRdxdNCiDGGZ1H+Ldsd6ok5N8aMpuVbmAJO84xLGC9bk6ixMUGShOwHpv
KORYaCzlyGnF2lG0RySCuaDGx2nUR3S/uqZGSAeIcjgHRWgrn+g+YmxAl9aGJ/XJM0ZXjC7DJ0GF
8CT1IZHcGWm8Q/GAp/HK75NPiyVsMTqpxcYrwDNYbUKkTLMHMPMc8pEnv7VYRULhfMI00y3QeNAN
cKEyGB79soTe3Ez1X1mTmh3doW/Q4EfUCos9vms5ze94tsVW9xswehg3HicmyjzIkQ+8+XWvHdxt
KWl9c/Ti1vcOLFcstocssa+oOy3vDXf7aEHsaFcOVu123CS2YIvjzvuHSiHAWEr6mS6s5M4HHFqL
q104S1gdsfU95NZdhJYj3XVJYcTHkQZBKLf1OtqjTxialXfaE9uFI3wVO3tunpKGCb6eeVfCmM6L
4S60XNj7GeNM1JTWTF5ZU1x4EX2PW+ZdYJOvn9XEsgfPlzL8zd/mjPfFwWJ8wFml++80egcFXgu5
XX1VCfJBLZmG9Mz2429c4UUdLEuX/Ncr9MLaXNSUCGVtI6XO8ucAl7fOfy0Ao3Oht3nKEfONnems
5/bbACAR/PeG4eqKtsg8C8ouQkv2BiUx+k6ao4HsQjOLK4u/gIE/wu8MSPZEibUJHl68tlTnD931
1HJe1Yvdy0PMiFUfhj8i7EehYH9ofwpCoC/9qqehR6zgIP1mrAk4cUQim2/PL8I+sgopGanwmb1k
lQCcUFRKMhG1jDOF9k6THw8e9pQ+ZSYcnspQ4eKAFFyPbYm/yg98F9yVEwTRUNgnJ2i/cRazTL/G
H9xXA+g9zcuplexQgW1bcbS3HvSRVaSeJ8fXfzqSsKGyXG9m+F/1S5DF3B5Y2pSOOExKzMcE/ZdI
d9f7gswwsyD8SV8r+oJh+mAw3eQdRBQkifLb+n4VhuMjbbdt8JyMawvNxWHvI6tFywZV4lDB9ZS5
a61biV9L4x5hF6Q9LFHiqxO2xiT2RdPflq2YA/pcQe23xNQgv9auKqtP5YOrMnG9dq6a/QhDJ70d
TVU3O6dB/n80AW0TSbK9G62KpoO7432bmL830vJuf45BypWA+Avo8/oddAb60TSruUMeSeqHiCMN
BphpgRqj0DY3QzKv7XNAGRskxK7MvtaUrJPPuLq36f/frYFKr89ElUDkA7/yVqi2i5eicnnd6LRj
GlNObdQloLn3IKj+hhEeWkExhJsoaKgp2G6CjQrnYvXEnp+9p5oswn294DrviRZSOI14KGKvTG3o
HTMsOyvh/PgSrjX0mRPTcUB8193zBjpxxyfFn5RSjvgYIyTrp6dNPIDDuFPsjfdF8LpexwoC7/el
bEqC/SynqBrhWxzdB83I0AMC36RzOQyO6FfFRktOSZLMhwSnBoqh/f1JmZfrTB1rDJYxiA19GAR4
7ehwUmUcXrKP+l9jzUK61WcnhmJ8E2WvydsCla9OVPoOkKg/Bojhq2ERKgkuZFuE/S5bxHAeseUH
KK64X/lRI2969XeuH6jVWvFGCAX1a8SrxMSS4bQvlOc/ue5LwJmHamYAh6RRutE6qWLv0Fie8Qzx
uartxgWvuYJaACd9Qc8mU1b9XLnlpibRPdXHu+D+gLltp2LVFKgHOLT1Hd6YUGfl6m167Gci5lNN
ybPhWqsM7WdH4tTDGbXE8309O0W0RpdJQzNqxS7wz3OPAx2byu339+xeav0UtI08eKuaHqIDO21z
n6eDqk1dpdbB0K5v4AU5SLk8dHQWY8FTk8YOvhuw/KZMlHfHleAZbYIs+Lu1FDFwetuuVj1R+Fi9
iVsyS5Z02wNrHiXAMnr4/7TeMGpNnyn6twE5LD0JHh94HrFJER5rbroIP25cDA+HHo4QtF3cZMAz
9vIHuoOek9Nc1yLJUUhnypptkkVeI0hU954E6Jzp/tRmAfFpVuJWqCHwHyodVq39GD15aMMrKwnx
b3txmGeye7LBPEDjdU2LznlLcwN7H/KNFX6uoOl+J+Da29zi7wiWDZdmv73cxB0dSJo5C0x9utw+
e5AKv1wlyb5tcA5ovPAu/0TEwxT2ieAS29K+TLrNbjC4JoFpLP31JnDnKXhRrjAJ5NU0/3oHH65O
LwWqVK218pGkMAse0OV6VO3eEw1Q1FVChuBKkXySD5Vsu0vl38Twim8bOktrNFvRNa6VC+y1jX6O
jDfLsVGyzy9Wvcti0IAEdhzI2JYMMWFSI/Rb3R7caMquja5AGqnh8otonVtBnHzrwE+KgBBykRAA
QHuyULWRdj4Vm2ENFvC1K3eVuuDKURDr9X9PHus6kgdgViTGu0LTM86E2bGpKPNutSnBF7Gv+Io+
TAPSSnfd3KSsRcmTWn/KqNgzwChnSTjdsD0onMiLta34ye4ks+u57nr5aD58ZRgJZE9t10/RjwSd
bAH4J23SGi5U16nbZswRagBCZEKJzwQgxmKxLGtQg54SFDm0/RVgXIHLI0Y2BBp7qJbeBAQkbOB/
fyyP9F8cWMpjiU5FodoMaxyaMaQFXBKQ/ViSy0DdNOGYsRm1x1C9gcP1JEPXWqcG0Xh4voHGvWP6
96tN8oWFFz2zV90cykAs14t6plmACrh08AlnffQvEcRRJiTWN2qGNSav1lPK+vSNvUqxGwRquHgz
DhFImDhl8tfOOf1m8CNby0UwVYRP/mUZAQUi3fGSx0gpNNywlHUa1a6rNIe5x0CoubgXSBlQvgFz
P4O8Q6TWuf1iBz+QNp1Rdp0f8Y/JCcGBvCCDYPv+8mRB1kndeZp/v9rJJOQWqtEYObmnBzW1XvZP
jbzmtCvHQafaFeLCzBJ2hVSkJE92a4EpPjmMeZBF6b5PRlEvI+ZqxtGvqUCODn2+r4mVYh3cLkdF
JImWAIqLr8jGO3hH4iu6pRZlkW1NZULptPRIHEyWDysAw3RmucabZ7U5iotrOLQzqImvMG0J6lXT
yPOUKi/Xiecp9uWX3by5b9nVt8No9/BKdMwvnUZEwqjQRlr4uaX65sYYi8DdTQ4lOjyb0PXG7GIb
89RCEMazxb5KHRRYWEfHbCb/O+cAuHM3N1w5WCwHRfv4JfcbZUmsXv8VhTv0LabPL+sl+8JJiawo
aDOmvi1auzW3gooTmFuZbWKTOsP48qLlHa74pVhZFkwg1r5GzpmVk+e7Vo/6KlvccmWtnJptf0R0
8huX7VM2GmZ6DF84d4pgz3nZ8CafeLbU9N8M+JTBUpISobyGnEHEU2cawDtFlwvTLTXWDOUY3Qeb
T08cRnlS3vssE0G4sV4WpdT5hAQlDO7wx/em1hlXZT8/3Usq7GIKOLxV2rEXDuRE6aMpHL9MzAeX
MttBcacAJJCtIsqK1gbdLJ/N7MCfhFZ0N1JhLIA+8ar7VPwRB4xwudoti99zRh3kDMBRVak57byU
nsqO9/GVpWjUs3BVYeYHjbhTThU0R4qHNxTE1cxhiKVj1mxu9MSCxFSB3lSGgOvhu9LV+f39ykMU
uKN9h5joFAPp+L4biWTXxQLUXk9mGfHBKen63HZ0BbBbdFNlPkFRE0N/rAtVWKiZbYMrDKgCgz+W
vQqD33eLBAjDRNuQM2x8nFczlgXs8xteaT01zJKjs0ktKBh1KKey/q5hzt7/U8zdKUiFiPMGd4bd
a5iO+UW/PVgZqIVZxhH2cF0nkJ9c6Px4+RLCazFPCSuu89+sEj03Ii2azZq/8dOVTiTY5zJLyKab
jY7/hkcBT4aEvYZnTrvadX1MIYM9EoRWjdJcPMHQLKUc9Zbek0+SUyI6s/rSX6tKiPKPGSY4gXKo
rzXOfIIxUhCNAanmG2yYcSs2Zq6IJGmzZZEsCxCyn6aGZO0RUv9UsKarRnL1ruzudVb0EgnXfIIE
ktP+8ouok4DGCkGvcKS2sXkKCMTzECrjFtARy7oRraw7mdPpOm8PazOQTY3f2FXN6HcFCvEGjrVN
iKjYTFXPeYvHO66LrNVx6GJFZjb1ngsEcF4Ld/4bltgQKsSlSB8CD8bmFUVnVbtIhFbjKqVz8JmD
iGY8BFA1H5b0xAWNcwCldXwyPQTK5S/nxdWyKXi0SrZm4MdiYIVPvbA8L1QvLNe7IuSLZr3bmi2u
XLX9VKZDyYGOJ20YYCspCZTvEyWcRJXi4oCDw68y74b2cFeVvyhDHcXm2MzPctcPWX9VnZiw6pVF
QAKenKiOQVj9qY10nhXvaY1HgMQXFSyeAiy9loHp/zpECTc+DVdveJoCdDLHoSeyF7NfrZ/9jak0
FVNinDBp2aVR+LA/j2D2oEngoZsMtZ9TnIjRra/9gGhz8MPJ3PP0xDd6ykVus3Qqays8tQMIx7as
cdJTwZ77qndmDRzbxnlz7cHkzgF1AMripplnokY3GFral0RESp3NdrccDxQIocWKrlQQV2NrVl7j
BtUIpBSJn0tWbmvDwtVXzXLadgk0zajvPx2Vm+Z+ozTtISyusBxkWxO8u5+BuixSXUOsqHkOkiix
4Xhq1mSjIyINt+fLEIHy+6t5EaMSKqEDr88loXhvylagwJj6odyPFIiaS+EAoVBklgWNbtwYbSjh
X1oAclEct3tuN34mJxCC4eXoHotaezNGRKfecDoW1ITLYR1zlggbnh3rRIcgIJpNk2RDipo5EBAv
ST2qNmGRB2jOdray/fr64cvwYDQHyBB542mA0bpFlXwB26uUOvpZuPnJl5Oew9mv+1GYt3EEHTZt
JrjHrw/5qt3IsVXzPyl3Qc5emU3f/btjofl5OGN4c7Bus9bFEj2W539gkxtspvRxRaEAnmZOs/Hk
mUKJiSjwZLoiWz/Cntr56rdaeqaRW3FIXYH+EN/gKWzzUPWRKjUuIGKXueOd1Jpq9SG99YxWse/6
2E2CrdvuZEiH8XCAcEE1ClcXx36D/H7FctNHTVTBSBAi/9/QmFNB3e6SNqy4EWsIwQ93SdIDiJ2M
gkyebzvKuszh9vinRJryoEIygNZAJgZKknarffaVzF9pS8V+bKJ6/t2CG08GeoAbBiAX1TRhXIwa
WREXyZxkbp+WqvqlYY0v6aFuEpU5MTn3FhSXh1qiKf67NyqionXhtxP5HafmMKkdQ7Se5cWa0Ume
Cz8w4vgW3kc5hlF6eK+P0AuxDjSzrTAItzLhO3st6E3hEfEcrYdNH1MsqbX4BXImughLWzSb5l7n
9A4lCu8KsfRyr443BXpvccCdQl04LVcJ617zBVfIz2m3hgV3w0XQs9I4lYidUBYYsm0oCHuRhS19
r5s61maNaKb/srrIxiBY66qmxwjueGVv+ceojIAHAzL8qAeO4rbyq992Oz1JcFuL0+fsoAr5oDzF
QMsGyPiLGg2DuT8xrmbiFQjkxWqDCeyMEqDR1wxQim9qXzbrRDRP6J0xakSnRwFP/guEVsocl8Sg
HPD7yf7pR3gyogRclyPlwdlVtIIVUAW02CJ6DUzT9OwxdaLIpbyXGSnxKa6N0lC8qRM8km0sYNAi
2v+rujPBxuFhyXv6WLxfGLnpPC8+OCJclxmd8PPwMaJriO/74sdoSRd9TktQ79lJK7yER2/pROgm
GK6WGs7tvW6P7sdXkPXT5D+2sPw8jV01akNSxfoKOXJF3uu7AGzR4eh2lSsASVbbeeYwhWczqmc9
mDQISrw0MIcereqJCY7hWBFMtZ5ndRadappwYiARcFOtLrgrMo6Ep+QG3ubnJRw8QSnP75b7PRsy
f45bkxvTH6T8r7Kowd3x4t0DrY98mXRwLEoAeh/cgj777Mt9JwEjGEqzbtEhyly8zLZiAkBEA08S
Yvk40DhOOL302xnL056waCkJgedi8cahdKFZ8bHzE1xh7y82BHVtxusVZ5YccWAb4xfozc4BMKnq
kf1xHfTe28mprEhdlLdAFmPrfx2t4yf2TE9xwVpgYKBHoxUaXrPS3Qj92ACQDs/EOKDwxXLxpP5+
PECvz9O8+Qfx6MXD4Oi/GZkD3RLTiuMwY2ZvgggTBrMG+W+M1gqadcpqvAL/b0Tb3BZj5zK2JLGw
GReqk3IhRr+GhrmwX+MV59KQaKgeYjXLJIUcO0CoNuJSLrYLcvNmr1iyfsH51NkGZfqNhwpqsplw
Sx3HcGjY811FGYlYKvGWh4ueifKcv5tbJ6uWCaDJpyfo7IEXw10yVz+4cCWGXyrKI5foz+abIOfl
qVyrKwuJgiNju5ohHo8OotfzCkxxX2knY9npzW4Au2UvTURWjJvkyj/U8gbL/AcxnmwsP5DKe5tI
eQVoMtbzTUO5IYU1akBnIzHK2ZjGeVVNJH8DjciImkGSaY6XpPuu9nckIx3EylKVufoj2PD1tJX0
yQlGn8DLQFYx/mseIpR8Jo7WLkOlrVgQ72S2DAY86IP2h1epk+OMbMaJCWogG7JkP+0WpJPNDoUm
MS73SN7aXA2wy1wyqQoq/R1JeukFAjjN/Wtq5t7iJsRvQUvRiiSwEqt0lxMAJIsDpKZ2OJ8cfuvg
xRUbzJLaSpQDpoDKfsPLUgKe1m9vkL8WWeKU5COFL9T2KiqiAoiSdj47QfMlu4F2nRmmsCF22ZJN
X0rPzCHfd6n7xQKdGvugu4P3ytXB3+ysscFGOT/6Lac00S3hDZWcEDzkLu0E8kXUNsZNX6+IqKZ2
uaIFpbWq13z9E+yE1FNcYFUT0jiWdwqFfU1LZ4a9iG2906wuQwGjwd7eGkM+jGC0eCM8SG+02wSu
iFal0ZErqnrzGSW7XKLfcrp2MnJN11BtXSTgafHb9ZnIgxU96A5HACmT9MrYGdBP9zFHwm0ONkb6
9poQWi+G9sZWumxLXA8bnNrn2d5Qu8I0u1sIsmhHPy6hL3o+ryXggTl2RSWyhamRNQpDPMBBYOwD
n6W6jxPzgQVR/cc1Y3LtWaTl64t+rCrtzy4bBOdGTbrXwSWRU6iwJq6YQUfPh+7GyWD9NzkLgx4h
YewjKQLwTpMPWx/0WVcZSfpkizS2WI7x1rW7GcxEtI7XKo34QgxW87xin977baQPyB3AhCkYKxhn
H3QHWNq4wkM9C6PjDhBJ64ZczpLeSEHdmCmQYG1v0tA2sRAnN5PVLa4PWdUPylSb+Qk4nnp9JX6y
q0noFucSge1bTQwLnvVzcIU3EHWZUduNUeLHHAZ1pdmdh1+JtZlAuW2SRXiGs86CnMcTOrkAhu1v
mYfi8bNAN5PN2QsTq3EJWdNKeYhqWPL/41bbM2Wr7KHW0u9/04Zqnf5WMX22GC2DSZfyyaPwmq/Y
ziB6bpnai4pGiRGQgcDfAjJldnveMA5VjeHsvvh2e5bwk/IvtIL2RfvXbse6vxVZPD2TA66EhHkj
+8vAcHxJlumdct/g6W1wUXa+1VFJCrFAVyKDJFb5MGIF1C05bNTx+awJb978KyppY9YRWFgETu4a
+MAeS6ExHTmP6cNuWFl37UWBbyvvo3tOY9vixOZOvvMse8/TewMta2Gf4qAiZow3FVWSzqD3PxzA
QElIpHpQBuQBc7BTy7ER6SX8Wm+ang3ETxNQAwtwUQ8SOyakn/32OnuVknBfaaHGMGHthBIut91L
WUFL9llljHkCzkQ4GUPPcFpj2jbhIqmenFqYGNVIxEfwGh9kFyWeUi/dmdqskh2r8bUzBHERGPue
gqvDS+0HAwnY74CfJd2t/utp4ICjwEcLfAeqNU7OSwXJu/Fj38940/5ivFQqTcq9+pUSe90+gBQn
X5L6F//p+aVyGEHLOfQn24MdhyqzZoHPb98DPVZSWC+8b2i4L5lFzsamzz8tm5I8KCUg4qRpOslm
u5h2nkeCdXuPXutrgDAgH6RGfL6JqDiv8Iedx1/ToieSrSOtsLPD70iJpKUI126SeG010KIVy+E9
KNPjXNP5GHTcf02NDOzQaBbWxkDvohlw41YuCpJaxh2zL/5G9Roo0jSrT+CwlvjDo7E5bLMcPxor
UxtT1GK/9V3z4o5xTfeSbUff6u0ElNL/Q5c+CB7hYC2H+HTZMNm/i4vZO8g0ywkG0dXYjlZcGgXG
V7jP0tJya106hiz4/oUL++bGuAi3j3HRPqmPG9L0r88bsoedXxN1B/O2m++HTii5ATLfCgDFxuFj
KtF7XMMLNJzpoH+uQlSStjazJm6XZIsOa9ZTcswzXs2y3+BLRz3EXPSPfKGPfGgW7iya2NpDMpJQ
RlZJsmzjOy9N7jKyAR+VQM5BFaGug3LXNvWkOMcnSUzFduDg0aK1j5SgVULuOuwzw97/xrk3xsHJ
/5J72QXeeiksgdZMCxVTDGoT808j6IlGeysuzEudcYbWXUPEntG+t7K8q1iAZYbFb6B3FAemJdI8
4WUWUK0ojLPfzenWqZxnB1DgJiHu5vsW1psIfNPAn1t4/g1NBCrEHnt6NrYQva0T2xiAtAnvtIwl
Xswi626IDAXNi7p6sSBb8coAlQZzd9a7W20Vi9BXU+5/nf3vaPw6H/a0ge2zsIbL3vklIkrCnw3b
55AGglhy6YSOLFP1CDwtUGaS70QArCv4fO8iQi7dVBiyfOyWhbvbJ9QZAP0vDEWvmU+3WPB2yX3s
2GtJbY4F/7EPTjPsTIuceaDppLkty+7R4teOCbSnmpyfJ7ToclcyRYuQ1caqyxUK/rqhGAPgcCb7
651DMCqMhcDqT7AqX8GiHeb0b7XZFds0qy4GQveXyi+j5xlaNJgiNGQhE5laxXmYTh/vzue4IbqF
0buvASpz4lXVfeApYoX6a5GLZzNTY9WIKqGsCSyiKbc2NEIpwjJ7B41nh6+3LhZEKzIBqMSamSX0
kJqWW7d6VO06q8joBHRG7O5hTQSzoaHP/Amlm9f/Pr/G97ALU52N2551W4Z0Qer0zI+p+105Q5Ic
68TWw6J3dtYStoi2Ni8phPY+tTpFRy7isMxOMu4W7RGm4u5HUOrr8l2la4f9/EN7HqvHR8npn2ND
yq4NpK63PChny01RXf9kcwOzaZbICOo+BGkAweArHmsSarkG8B/RCntqLChp+ltGus8/47rbXwri
9hZ+eHVlTvOQWKMVuCOc8NGXMCfl4z7fWB3pBzF2SNPWySCyyf3ngKVJNvifFj5ztemE+pGXRxpE
JQjW3YBx1RsCzWP30tjRQGlWWKOA1WM/gbGHNTPW5TQdeBA2t5NFUVaVpsa6jgHcLJXf6njUeXkm
7grSTP5kG2oZex1M3rYl0D1Xi5UrWxZXOxFnhX3JJqVY1nlscJjVSm03QiuUlaEnVrO7O5L8UNjG
QzT5xno4HwReaVQRMFmSmwJK/C1hkDKQSXHoVunoyq6Gtf3Uy2nho1T7cMdqJy5qVmo+qnz/rsVL
PX4XrkXphJn99FJK++K9hFXRV0qJ2qOtBnuxVCI24LYsrj2IMZOyTPRVXmiD1kGF2ovjHGEEy89n
dnjlVM8ewrorPyatW5MlYOAkDptLq4w8VXvuTMGvpaGVC4LyyvRMUlgGmVLJSEOEUEXnPz+Kyc3W
vWbJrdH+n0D3qx2nkMFIBg1k9IlgeJ7hb+Ul4LfPopsb43r57J/0acUIPQweoLQw2o0zXdWHNRF+
NV9wbU53IUy5V1YzHWwqgo8zcmDnTqTfbYMk8JR6ZoAKsELQBZFtok5Y4ijFvo0CIWmZMUuTEYeH
JHWb27hIfkFNi7eBE+0oT6WuE21ejfXh2nmIRDN0uhWxh0peYQErnVXqvJPH8rnIo9fS8m1bSyA6
kIgnzFVCAIP811gYPMSgTCMknkLXD3v5VYx92G2kJPGuVMXdx0ED93oLQcexFoVeKZXiuslYOMZ3
qL1XOvLNXK8dry437I7dvogUKUrEBCvohdGnUUZbdStGWo/Kkt9YsYk2NCk5hpoMQQbQVtbDyF65
qNIMb/vaCkWWJa524zrHvAT8aGr3gMgA5dq4jsuK6p3J+WCKHagr2S8awKS9h6Fl2z3cFH77nY1o
fsJtaS/t/dzdTPTFi+t8bbsDgy3bz/miVn32tPBjrP+WLzGSlJaQ1JyEggTiKt4a4WTEFmYU8Rrt
Qnx7Bj6MfTdX8FftYUf67eR8RgFzq+HgDIQP762ATmQ93pozlPcDDwqGyc9Xys4FRud96YZRbhLL
v3mMLFwQQLsJtTDQ9iguehTE4T1kXR/xA8+inPZvuxU7Uj3SWceMILbzVk9qEjjJdAdDEZba6oDG
hzQzBE90etAeAqiJK2G6a37L8fEM/K1lDxtLGyRZoxDba8XtZGRGDiVhZSFgkcfxsm47+rQ9Xg61
dsCXpr1Ijr7LVxaIfGPBrWrWCm+gRyJngCpQKCzUapJrpMOf/4kOMJ6q9a0JE3CI3my2x5M1MDNb
pdc6xMM0knjbRkcm54xEflSmDL2uYRhXO6lSwfl9ZYKStkEHDmLkPYhYusY0vbsF+SI7ZsEcIOgZ
owgq3Wr0nOZurTxECpHsy/2OkDSpKNddhLZjxLjJo5Xnp9r1fuQgTBkcgvSgP6pVoRVw/QodGyKG
PNMMO7HJedQSiazxbKjN8Abk6c/YqvO3MIt1MrVfWTMEcCPDTgxAK/N9oZ/zlkpDGTwVdh7lZx9J
T60gdy7pVIyw1Q0o9p/mFZEmWYDVA5M1/slsYrU5NsnL1CtfJXXpzIwTzYNFSH3n0oE/kBkAid11
flCF1NeEWafAAMW4gmGmH9/VT96o1KZmr3/Q+TpnrvsK3f++5ApnphMHBNSlIqbXrnh3m4JpqBzd
RDmgfd9CbFbCtnsCGz9Mmu0mf9MUYjPwpXnEJqjYHk9LMKMh488SuSv0zFnBwshW+npZsEXHlbQO
ruVjCwJ+kTXUVFEJajFE33dcW15+0R49fwJHLMo0Eo0tsxa/kSPwzE6MzXymXNbHxQUYNFd/Y7C5
vYp3wOQAa1ybhvLNq1aQz/6P8r9UUVzF/3JPAp0P0LZuWmJ/1+dPoYFMYuo/DdUL2LTx6eBuNsHn
LZ/3kKj2uf3tkwj0qzN9ouSScm6cBT5w6x/wN8SKIpiNg49PTp8lryPv2Gr933yHKwwAJjNVyRyu
DexnkY3xHuKtNnqJiDAPkZEVtsy4Ad9sgqW6tlIubp8AMYaGr584ZDtTefSxk6QjENs3e5b85xxh
ebk2DFgEvI697v3P38hzGO19IfD3vojmwZcrmPLrE3s7bU+qjJoDtc9XjyR8TkagHttw/NbbS5z7
HuLMzWdMUPZPu5wvWyGzSj+XYkypHKjhc2gBbdL6lTfP8F7oSkS+Ag2xwrCy4UQOXNirzYVBkMyw
CsEMuvUmApVlAofN80rKjvpGSWpclEYbX2EC72nOqSujx3ioHkIZ/u8oJYoyd9ADHpgyqvLESXVe
GXYKFJjTFn9Jzg/CYkyD8o3wm3jE/18jDuEbrRIia/mzf+6vMinQ6w/Epk1tWylFq22/xfdkF/y2
DBmBIt3Iy8TMdLOuvASY32On3YpKlx95J4qM1knkhnb+gfrGFSBk4YmWXy0NpTKiO4PvKXtDh9kr
22ruC6XwfjUeXSSJL6xXEFKe6cSERBsahUXdb9mCcWdtFhwJIs0dOGoxSxd5d8qwSGx/YJjJBBlJ
NJUsisadQA1ufzbpxgoNsbanEFow2nL0nMOyU6ATsa+YyVGeJ5oFZniXAtelKlLZ8YAI3jn/+Yil
PbJPpXKV1F0CaUBTVQXpZYFf9+6yoCOWMDFmYky7z42hEkJ0468fUDiZLMx3GbF4eb8WPPKZwpos
e5S/JaQKgqclyMnz18b2biRtzbgKXRgp6R5Kh4eu/ogMxF5Ummf8mzwbLhC86QTNO5W+Vudc5XpL
vLqjNE8BPxFa5WgOlcPiOKMigdKlGiFTa25iRli8tZIX9xEwjd0FHBx6IrgORx6qaBJyP+1QpfuO
Mdm0Ee3KS7NkCkZtkqIDxGZUZtScqR2FNgRb5jbKW8OAtwEioNVzxc+5nTgxIhY9MGev/kU0eyZd
U2PcZHLhNOvPoZBgbsS/fF2bjG9OP7uugQyORait2beI+IMzpN2aezgaf+pGNs69x/+W4a/dowLB
28W5HxozoiAvUVkwaYnmbSdxbBOSQIyxxGNeXZ6dKwM+yBUa2166QDfMNSGBi42DBrUfMJymXQuv
ZwmGkNjps4fyZH3zTKUbUEMDK5tYEUh2iWgoYPDRzuE55USzESCAfOLf1cfa/YxkfHSG1uY/0FZd
ERu7gyqwFgsZO+WDcG87oGIrje8+yXuyfErRbnMHwIvrTwcu8N0LtPM56mq6EF9cDlqbhSKwyyKe
C5+rkAgiDf7y0t8xToXf/poYkF3s09Iue8jjvY6x5iot9DJsjln3nMd2JrpOATCt6b9LSxha03/X
WwaRXK73a6Kpp/O+pSMRYBhULRasBcLmyBV2bW/1aDLMigeYEQNHJ1YW1JdrrfCzDoD1qlTCR3+8
2Tj7agcLA7E3P4g7EQRaUxwUTdCm/axNnqTAVL1iX5MydWmmiJBDYGoSWnd3nQ/OeH65Du/WC2HX
XyWvsIoGTbEqnUI3MAIqRVLUHY/NepbksJjZAzsIPnxSvmbVzKJ2UCHLb/IXwz77xAKZUi0PRmuN
iaEE6KpMFTdK5SgYueIxwi3PwL9BTfQg7f57+msVxb3J7LM5t/H12AIvHUmSugZ+CYHcysvIVKkt
AkMUFZS4s8+G4m3xl9D0nTzMoU6/8+rwgiCugk6nqsb0iQWsc3Bevwh6MIiR1y8R6wF9SInU2RWT
ZbxVtPv9htJqUDSZLb66EVR52pvSk83L84Y7LbW6UTNJZFb/8ftweyx9Jssdrg3DRZhpcvVAkM5/
x9ceHhvkafiG8o10Ay/JjazaTyjjdbr86v0ypFbNpaH2SjatCwVdKZvajpXSYz56rKFWq0a+CJES
IhaNAqPJg1ah4iwbdtz3S2nb8Sh2sQsaBHcBNe1O0M+ANKx/qpGaACqwPAHDQKsavukSVp7D0tOu
1Xzk5vFQiMPOXGjegzvdOqk6WPNZiRLprQQxmst/jtvuNhMvkmgKB01H6loYhDW9tUMrqDqdcB8r
YhvXkUHZxlqKpYvn/hDBfWhxlx6Lpn6wmYnjAZWlwibNi4Ceq8ppo48DNIZ17hCksbjezHrRumOT
L6EJR6lQZNqBMrSz4+z8JhVxD3a1wx1cttY1ZfMYBSeyOvJhitulFSSS4qVfrKw2zD4d6XUtGfrD
T8nBsjZ51sy4qWXLBFpwfFPMgOmhax15Tapp/5c59WIchsJmQR7VOVSmrFQx7D7LTOSeUzqB7ePr
L65/kLbZ7UKQNt0r5cla7BFd3yKY38OBO/8IjvKGfXrhBoGoPT41Cm5j/6MQ/vAAuJ+QkXGj/cHY
0DdsqyNbJf2jjJkkTkPg07xggGjCdSkkTJG90V1dlesE500i9j/ZhqcfQ70FISZxSxqT+1N1Gg/1
CVIaAbiufeWhiC3yaAEd8mRcd0nuCS86lvW582eR0fcccQOs7jEdklFl38DSuL38CTtJCbZnwsZi
iMUOcP/Up9Jt3f50h0Lor2zpr3VszWXV7i8DvVQZN/LQxm+oG3BQ4ge8Rd7cJApQbYprGAe7LOCs
b6kgtBSx5C+/wjhXismIgeV2dFEr+diPcOJToGgF3IzUUW4WOCapfPNH36DDRH3J1hnLFfmiI1uf
oT7yEMVP5+Td8YPX1IPugTZSkPjucz6ZQdPQuDTFjPZXsY2q/iZv1mq4hhczLecGmJMCa+/goirS
OqcbOrNodU+HTMXsOpy53HpSv02bAD+kxE2YogzFvp2vVDRw19nLGz5VRQwC7C0FIx5NLK1QEloq
y7wL4eMAiyAqFRn6E2sj9bZbLauKKEyzfL7ZrD0GlHB3m3VXHkXk3zjMRXLADDsSFRUj0uQqSJiw
NJXextq4r0X8XU6T7lhDNUfnrx+mYNnNk8ieKAqPGeh9k+nG62To6emVMrn2fTriVts6bKlmQ7US
jRbEWVQmZ3S78cAbw5SBJtsjH4yg0NjFDWg08y4wSYgFQBHxLBjqakBaLl/fz4bcfzTGBOAzcvBn
+tryVMgKRAIl5T/NjLbi74G1/8JR4lGQAJJFpVqK0zgBSRubAC6QANksWysRt57O8GfXrLkZjnyQ
UQWbxWAoXqpDvP5Mb9KcC2VH85HppRiOSmruOWcnomJIBLrsAjf+MOlDLoNoW1IEFzXNQzCYw/zK
RNwxUGL8dRnfzZXZU+De10YfWBT+Iorp+oZsTJCsFpqr2Rm7EbgC3EijDycCeFI97NSm3z/1rpPQ
e+UTarKNLN3coepij8tooxBHZs+r0itwtRnlT5ZeTbt5TPzVg2euaE/8ST20hf6Sn8YFSvtS8ym7
tpSB/mw5ND7MftezT8b5vRiBN5OT8AinpSoZmzYxlgHCixSinQR7bcA3CYhTFmyDDaQdfaZg8zTh
4FRmLRB7vAtDVZYRMAfffxFfRBI5zKCZhZ32m3Z1C8LmqJUrC49Zuk+UAvhufg0axCa5bGBvemBJ
1Q13+8ucUc9PADs+CH/dcRLTey2XrW8POBHtE5Leapq+PtzFJtEsMY19K9uUos5A7RfJETpPtvtb
3A5TNUPQvfohQmzPUqeOFKOU7QJkquwHjPy8gmZaGZlXGSxPlV4xhqBf3pyTizy6quhKV/Eu5K/m
TNKA7Cqv8KUqXFAjgSF8Ha83Q4T4O5NvFtVkq9JV5atXWKB8hUCLuVTd4bDzMuTwrpctJoZzDC+n
QyTcLtFA4z8BpGxemBOgefENHjR6ECeB3jnOLLT7WZ/7AfZXaiZ8IwHzYLgP1ud1TSnOiFLajrY9
AVmUsFIAls2qDxZGTSuSflsza+bEdlBbbLAtM1guqD2wPo/2eEyuMfo0UVwoi3SEIWJsZ9wQCTJT
NR/4WXslImzj1WO762M85IUzhjyPD9AZO93PT3Ub/Ui0RdOMJvleBaPVelp4I8M0djH8+rUCerma
VeO7LBFxVUa7ttohA4RK1Y/pvDvO0CT5atf5dla2dK/Da7hgTKkBbJ1v9hcdMsnsiJyErUDCQhAb
/20Fw9GM8OqPIEQ+HWn2OWPDqN12lfAEuoMljn3o6nXk8TsSiE6SpBUtli6mhVHPOW7jmStgfAPQ
zWKZgE0KTta/1VtiBki03lAkoRn/m0q02ycHTMHLJ1AzbdCJQhq+5dH8UbOcx89Jux2/xgEy9X3K
Y2yPgI6Aam5kf0s7rq21NEzTJbxX13sIx7ARlxen8I0J3I6u6fY1GiaInrp0jEtZ4+OFvItmCqWa
SkNVVsnNLhLtgVbzr0mkPw7qas+EZFm4V/hC5qIa45VeKWP+9DawDqemW8JLDtwPWNuviY5jvzal
tl0O0f3O8r6TF1HZsk53ODXx7IqfcVt6xbRHJqlldjmJhUvvq9Y4ZAGOox7oDQXaiZRQ801x+xcq
QtnKSeIgYskZvAVi8TBZnRGppSvomyP6CPfJ3xd9W2tUTgCH3WGzlKsmBnLhptm33aY6cXMB6jso
ov+T3+acv2tiRI8jmyHvX5ywR+7oZ+Fb+jT4mVJ1rXKsXy3tFTwNNtS14VAdhLO8tfp+AOqAlGO/
9fJtti4bcp8iG9MEvRIqzju7Iylic2vtivxDxyUxpebfYJeGKm6hKCy4++vdvnbDEnuyRSTOG5WB
M1F2QPENSEhrCly0POx3ga1bOcNClRJs9IVGIG8klg2vC3Asyjpq0ZW6rIL+efFbkChiIb2qRzPN
jRw7QqDkV+j8Nz+pZBZMXvQLDjd4P8D6c5p2xionjaV5SVJ2HDz1/id/UVSJ4ERAufrFDWxRwt5j
vDEeSxObfRyBdHACOvQaWYGQ2LvuJv02ek3NaSW7GARNE3k5ajfD9Bj2aYc2dh/oEIHh3G3Vo6zG
wdTNU6cqRMIcb659QDcYJo4t3d5PFXxFf3MlLWjHifRw/K5bJKTZ5sJVoubLIkz/HGsTahY/AeiS
jJ3DvIvfnMXA8DQmu2yfSUzuzIow1OQ+Mz0BHxXhEUGkW3TIvcFw4ibiGiWrS1iAOYumclD2uBGL
t97Vz6YCqlPkEs6UUnVHL8EMbX3ycKcTLvND6hdy7m842+/TlxBGs0VNL5RTRx6QeYq/r6YTQjFe
56biNWq15dOlf0eO0HjCfU/sNKf7I2f95xtUiuZUIz3CLF0A5PuEsDg+FvP/eSZM4+YN7hpm0702
EGM/OAs86sMw/e4l4+w0AQcAsIwtl3Nl6KBoc/71FjQK4EHSQPapJbIxGJUDqIsS5PFVQDMnLNHw
odQghytcxYpWEsacwnISCP8jx2yOkMy2PbYrNAGh3zvxfaFrnTvJlQoIBy2pcN+d1E0EvHlUe116
k7jYqR8T22irdnPRyXTsrnuelCY0Y+0vfoGiTqM+8OPa2rxHvHF8ilpyy5eGJa9ePHarOSK+cTnm
ZOD9TxoM2pnL2k4jOMXM5TcVU4QhOyi13fsjVUZsC3e3YpVNoOvjVtOjiQfevxOMGTXPd0Mp0eFR
DyJkd3Or8eRiE1+GINXqs7/UvPNHAMkA+DADyLGTmDH5iFf9hbt97G3HcCHVMp2tskml97A2DTe9
3uHqL+D+3yvkripaChFnRs/ZRBeBBiV/2sp35WrgrkbQ2O7dVp8vivO+Lbdp+5Q4RmfGHpw6JGxf
wWEQxCB8N0e++PcJeaJxRfqqpM2tY+9MJMXghVPP6e5wZhtUj4ZdV+mgweTq4TmgnviEKb19h6kN
cuL3cYFb08vNcATvsaMH7ZFcMxUBKGqRmrOTeQGfaMzjogaG597cnZL7BHf3ET6S5m+xcSe3wSdw
BY4zIVZL7Quva1oBcENW6exBOv5GyFc07ZzRTaG9OmOpkRczhn4KBBnReLGkfOB4tNSxGl2BmtPa
C2TUROzegrS0Gq1i2pmut93KBPh4eC3hThrwFaaGcp7yo6dHcGR5m6Vt0GsYGhmshPrTywRq2r78
znTs6EyoLU51A4ErBMJl/KGnzfTeRWSA6QhAdeWukn/na4j5tcumqKaHoaKSzNkYiW49P6zuYjU5
D1LdMIioNqN/+c/pD6DDpdORHUEHihVzOlXC9ZDwT27eIjWnFgwdqrEwVKfTC3Pu8CphLVWPOe1n
45O+C2oLEpO4ldtIMPh/GY+FUW/e8FNKrQxkYP34xdNalgyOJ0IFIxSkPzfl8TDnv4kH710pMsiZ
oslN6sTdNNR1AILGWLv9gdPrn5HSg1D2Wn1qWcdDO7teuBZCmGwmrasXrqQezN5ikOFYQ7rj4+X7
qmd9jgo5ShjVLSb1Zz91fY+LCXNdqsOew/tA9qDPxj0D6iE8JkgTHu3GPw7peytdCrLq7fshybWN
LlOlt6eMUVgTplJpr0zzxbfSJDZIAtZbnSrV/Tr2YZHY5vuN3M7NpaGl0usHLiy7fs352pemEQi2
eTbL4l/7w6EcScifOMYyqSeNg36sAq2RnQKoBuGPGhXnCmiNEYErD/Ym/61LCzgnAIn8ZQDzDqJW
y2j8PHPBr5ivixRz/TfNBAdQdA8BjehOsuHNciyDPXR2mfxeTtvu1kWZCxMJ3XBCe8PQcQ/Rn23k
JL0UlB8UkWulDE7SCUXQagkd2XkkzJR9777Z9CjQo+ntWxA8/G4alYv3tJBp6x8ituKEsYaRJCr3
xe+z8FDuLbn3kK4Z8kRvhnI0zqhPZe+wDOCo6im2k55jk4/+wuu5Dg/6yXw1XDuesL+53JZil3JM
NcPLnqbUDpw30mflemseJH8TYyOD+Us7RgwGR844RD9Sj7WGkaFBWCtmSzjT/KGLewahfcBubBKF
9/4EnYcQ9Ov8P/OEwh3Boa7MfunBTnqEqsTd6bSNpuOPP9B36sI3jEvXATH8wMSNPVN/rBbtQXXv
dcZsmmKH9+97y6ddzPK0g1fytkbrbXDNYrw1pY213xhjMyU4wHZDOQ8zR/2A4zc0m8J2gL2oZU6E
Vp4p8Q9d9r/DC2HP/1cmaeFe5Wk12TIyFZ3/dwMzrCqMR81OIcAe+q6Fo3hjt77UC/xUhXZ7Yr20
NiC3FI1COdTdBJUGPFKsgC2lxfklVLdelT7RjEPl0drtpOeYf3/VeYHR3HxtK7jXzrqgdklmsLQU
xfjpSzvzeBDM5O8c0JP2hGRV2X8r880oVwlzi/moaW2Drlyk6JRuvjjmzPA+Y58nlv4h8Qxl5jKV
VwiUWaDKKIFR/I0t5Zz7owQ50mmfbap+X9mP7UclzohnWYsyCIVT4+P2QnNLjujpNBkwd8C63R1l
ox31XhdohMYdlqSYxGaIANsQIGk6vWstpyuIs/JZUiHhgLXcvoSRCd3UajLmssPN6t5/tVmaUpYN
+G0I4ABztQLIE2On2WH1IN9CRqL0ZiZiYemWXGBKh3WYj8FaWDVjgK2hX/093A7gKd5vGsdoDa1d
ZnOzsm5uYHdFxp80jC+Kdx+oTSoJoTMZMwbZ4cr9nTWdssgCgKNyjsNe+Y7YWp1TLGn7dKsxqtTw
B5NHNaJsyBxmnihDmVRwIUzDTV/9RLbuE8JXfJ1Och71a66OxrQHRmN17Z8FPqlG+aSfv5Wjnb9i
blmyIPLcsVvGOc3qNX09z9WCjS9GYY1nemGPuBTaLG/+ZuUeKwjIjlaoqN/BRP3l3FYs3PJi82ss
Xxc/kmELk5zy03u5H3mCpMiZtZjOjs4yKXgpXCr/GknNQbLLEWJeTQ9Gl0wrLROEhRtHOfsB3P/B
XPJbpEiKAqZKCakezOmYMqfb5rxn3Q4pSqXUL3jb14zoQIA/k6KsPvrcndS6FTKGHeiaA5jD3Qwb
jfvi0wZLeRNCqKbv2dq6bwrO/5COcbTyIZUlEJxFGWgm6T0zY666bbt1/uJPFbaenYFOeSSPQcKO
7foHgn2S5oEDXVY9yI0ltZtuqnMyOVyrBNYSbjaFn8V8xR+/DHbdLU2Q9XrU3UxhINWWKDRd+gVB
p6IYOYX4FxduJHB6eIOIOGKOcHTAZlEaKwiXT3/U9sBz2yaAqT78iP29BmXnNVxHmKJ9RoFY8P5/
iU6GdKBLd3iyOFnMG1btuwL+z7VVfc6vT/L4xJsQde42qCcVI4iwcadU89FOjeknrMRe2fHT8Ugw
slzpk8ZmGzx53w1ct7XIr48JJ+UW1UVvX1c33ZFxgvnzWw3yTzm890lb5PNQVKpujk7emRIt67+A
PJtRvTGPpNgg7Qf4ZGgrKXDhjWe9y3Dm9y+uRMmlmQ6VjVtlDmAZYL0ENRZvKFGAJfw8zODNkf6N
wnDLCo3Za6nscO9NzMiKsxupHfjlGDOHXUo+ejDlmmfg3vjBG5GmVGkLOhHKVh5rzyBN9XJs4aF+
lN0dq91zwoCex7Cbrj2SL9FvEaTvB90BJUiYfib/OJEOQb7wL4/AMtri/bpIAj+OCwYDlDkbkE9P
XenKoVnrt7aDuZBwRU764eYTZkAlwftszu14LZw7pyQHIL/nBswdUmC9ztn0RXuzw3zoc1EdCTGx
O4zizDFwTNNrfkHJduP1E0Q+SklK5W19MkO+fK3RLV/vFmrOnlHOFJLrssrzUpEL8NcYJaVz53/4
2HsLe5wVHRjE9PMfNcA9EHF/4kefVHxhVJ72sHC2a+lKMOw+TOQSiPPpfQgd/X8kaAfTE85H9eW0
9R3TgXIJQaaGZonYgOT/mhACy2YisE+pvZjKAJrXi5EqqJtkz57R14c3cAR9nrUWjECy5ey0kcMa
R+5JjN3eTLX5sfnRI4oIXGGntoh8vi/+LmBGkXDFKJFjAxC+ykCEyu/ntMfG7BJlWEz3T3CNz5nr
FFlZTWuiYIhwYVaEGaAQwoWr/br3IL/3X/owWG/VlX5qMFMhbFH0nqR1NEf1NWtoeWJfPMWfe5r3
EGv01v0G47C1BIeOs0CUHPddrlmt6c7dUWvJ6kPvCoIbR5i9ucYepoU8Nn+pfJmhY2ep6HEm/QJL
mt4S0V35My2IDwkPdSk5XOKMX+Vhj0dJYDTMrMPXJ1rlfmGDZgFmZ1BB59uvaVtskSX3J+GZpnRe
Wk30gG835BIpv0pgY5jqD2j2kco5ZMTlQ/ODfh+BZz3VKoadesTt9v6freFCgRc+qv0Iy3o0YbNh
35snPC0g4sLZzH0KL6OVaTRwGM4z5QTPysf+UOQh5ebBTmQZJDxuKpBWhinZb755j3cN+xTzsp6E
JkzuNi6xrGcEJYvrj1a8jFob6+UM4vEBGtvxz8jzc3KtjG5TO9Qw/rrn1/bsv8W+PDFl45bKgO7S
SRkbC2Xr4FVn3lHQc6KovmlIUK3wx3duxr7ebMlWOeGpWWEYkofcKwEBowkC6w7blD6tYCJCV4WB
P9woTk4z/uTVS+dabRpibxdGZMGWtUt8a/sOnEBIxZT45RCESd5O3Vz6TEBy67J1MIGjpbl4Zsvu
8IocPcotfrehyXiz4ce3nPeGnVm2iDV6GdbHntFrNkIqsTUb+dHPjA9nQYwZvP5MisbT5/QysAtA
z+03C8PVV4zuL242vLXXBp3bzT+OaIqyABy4bBjm6Edh20BPI4F2yZJoeXwQmYL3U5+syTDRLVHN
rFZxRlnXWTG6SyZR+S8z+RQLvq37i1vwwFIvwo0A6HTgLQnbz9A2UFlo0Y9KmeSxNhlLTeEo97EE
O5zMIiNmLZjg29nRBpe3DfzPTjMyxA5JcqDY2fjFglzv11MJzavAT+CpNp56RbsCOQ5gDytIkbk5
0wAiRwDOreDCaJRiYPDuUjxz+fncdRq5qcij36fuvjANvpMVN3kxRumRUyFwnpo4h1tUyEAom2Tw
2ZEQiKBo4BczwZoF80ZYamgHPHROuz79ClenzaNYksG2NKO4d1H+HPOtwuSqd2u+mrwBYN+hus56
AsL6k3Rah6YB3vXd04ynxnc5L5hOcm4a7iNVaMWaeFN1hny0F0EKDwsd09pJEiWFZUfjCPcd2R8I
4qTK5II6X9GX6I1Smo3f4xceBJ4G0AbtMpuf7JXKYlaL6f7Zz99rfhUOh6oE/KHdGqKdPiICsz3m
jn0Mw1352FHI9UpRhKUROdMYjd5GOUrlPBpiB9bW9USN5p2ROamCgKjMrhdFZycOHzxG05Hasbzh
sg1O2KX7XfzADQMaUmwromRymmyfHjg3ozuD32VW6Qx+DoCHyf47f+m8KhvIeGB0JTdUEHQdSShh
PIYdPM8N5ucn2AbxSTmLqX5TUG5tN6etd3B1qZi3S3wuTkynWH1Fj+ynRKOuwuI+yN9Ul++NlrvL
aAZ1UM2Flnql1C88EhxFBQCPh38uRjqth93QvJXKj3Ba5bzxwXwzClvsB3zCI1v41xnxEUSNxXyf
2WTlSkfak+kuAec4V5QljldBwUt2wGGJN3IBp5IyYcT5XAnSqnRJT6sSiR4O7FwsZGT1P9uNLfj4
6wU0aw186IEVou4n6IaNnlpzMdxHRuiNmvQqvz3i7OuxhXnBVF8oAQuVdDyv7NlFZ99i8+Ii7GDh
ozWK8cGfY1CENXLUjN+l1z1yHkc93uj/e+rRNfpez0fNEm9yt0iF1PYUCGmDNuS2dQEfj16tO2xc
aLXdf5gafbmnS6DfFc3MUB0+AiPNNpTCfKxjYVHixo/55WeLhhk4D6lM4iDpaFfWE4bCxn3A1/UH
ogPTbfRO5KVlGUE9/RfYm2XtTJwJaKY1T6owIFdvzCDLEl4H73vg7vrU/sslxxOBf65ZLp8SxpF2
vBk0dQmIgVl7Xq575VkNcgMZL27dHmLPiXrFmp5R9DM4IpVJOqXIn3m7cApYgowIVBcWZ9dw9jgq
+uk2DzYc29VHgjbrVmg4Hg12ZNuORAXb6kCQomXlBxs6HAMhpJGHk3MyRlGtyhbbTJH2PGv/lNRa
hxT0oBLwsUAXb+MHweCVi/F1w2V+eBrbqVqpzd0PePkBY7x+hImY3aiMonSi0v3ufgIqM20EJYdr
LQAs0xFgTFZvarnOPXW3BY1imyn7YqgavpWSEI3IctyMwpci+bqMKxvxj80HS3ZgTUukgqiI8Lpo
6hUVEDp71CUg9JVjBtxoVE8mTedQ/beL6nDINoDEsR/5abq5Pi7czf8bF3/SqmGjIKQiFodUlg0L
A2hB4qZl7PcVdhXBwd9gsm9GTAeF0aH7DNq90vz6wekD9LDzzCR5agdCDabD0eHWuL6GErhe84P6
klR+u4awv+C+rvaIu1MZnwhF2RRpqO4nDhBvOhFOe7igCgllRvWVDP4RHUvqAIZ0zP24Ar8NRGJp
qE9Wt1nEqCqyicgspDOSjBX8k8V+HyfqYWnvSq6Q157sKMnBDXQxaj3Rsk5JhXq7SjpShjnlAMYM
ZLihhKxu82lsubUpq+JcPkcKpstY/zvVacklptjlolZmgm45GUlOOFiGsBVOdKntmUr/u/5Z3MRZ
y4oN+oB49OOEgF9wSYHq0j7lQBJEZVDoSV2egUqejmh+E5c3kV33BF7rU/iiT1XTRqgMHS2dnYCw
JXKxzm/Wx+Y364jOmLUw1QcKy1oRHY/6eGJFSugsdciAqTwMgLUYmFcbOkr461SOOfOCfEvcEowZ
vEJNkdoJcdnhj6XsF6oF8oLnJUesQOeoejoRhi8RJG93QxXMLX4slHo9TpBG7yYFHlchTVu6QEen
POS6F+8hB5Ak5UoGr5y9DWJB60OBX3RV7r1rr2UYU5BvXsGNCwNmQRC+TwH3A/0ONS3n0f4v4r6p
qrMSF3NHBORyp9GlVJj6iwEeF2rQ5INC5jnpCHRcZeB4QE/j7sONRaeBqPPf6u184B4t1r7Hs8X8
7uiN0iPKFoLijGPw/Ib8Wi/HY6QwooLOCEOKg8wAy4OYkCrj8PmFgi6h1nrQ9EpKtld5viDbnGcX
HCVB458yavdreUuSjlOpd6FAUSECvQoRzZpSH+bQsAGdO0G/H2rBnCtarOfGx7KpEItAyZcG06Ze
ZNALr9aROKnk6S+YsYoAPqF9NpOBrDxvYAGRNwEXedNAuEBN2DdmOYmJNuDDT+I+ly/MmucwivBo
7uCtTs1CzOEmDABYvb3feMFwHdpo0NUu6DjQh33gTYYP6WkcNIQ44SV8ZVxoo3rFzDcRXhCVt5XP
2blf3KXVmoYOnlHNpJoB4NRggoPNwTrGX6iNbAO+l9GcP0xet8Zn7OWY1xZ5t7c7ww2o97xo4iEq
BBKMLAUv7bd/6aYlnDeqs0kb3Sk5g3H4emyh2nWB70GbOMsTlwRuSNxI41E7QPFlgcwpUe+Lb1yM
kGCXXW5qpoA1BHQCZx/PCtFt5LOJ5Q0YGeHROdwXtA4NGkgsu1kZwyqW4Mt1RIyJ53pL8L8k1TXn
iKgv9f4QY9Qq0n1zkKl8/2sWIOmJijO0rVlQyw25bxt20mCuOR41v2LeOZlRcu3mdP18rfX691vG
azD+zaxIU76HHE/KRTAR7K+29JEbcPYeRYjaYCmwxiG04a+dM8+Qj9F5U184BKoe6rBqAP/g6i1i
kQfslFGGISJhT0XoanUM4UPoVHM7mVPeCzP8qlY1TfJfo1E+rFh9JPFzbldkG6bp0MqSYwxQcW7b
2QhmKKZWweSjlNtrdanBtMNAkf7rrNITvxfeDx8NPrDyWhdaI2mkcQk5wYl6k42KwCtt7jYNQ9m0
z/P8rPMtL1BEw8PUAxxiuhO6POvtREWTJ2ZJKr/D5AH5WPsTPTdLvWTv4cupu5B7sefYEnHwqiAa
ibDirpXdTMXlcbflf5aTM8em4OY+/Sz7hw3ClvGkQHmMF/2nCcsZdA3n/cOFwJFESCmtiq1VDdTf
EnR1Df9+a11nN4usq1bCsKpMqVcSzgltJ5HOjHRncrNVxh/x6X+46SoAOBYtOS3/taWJAPx35XnL
9Zc5umO0B6eDDPX4r4l5GHgdx5+o9JWHcUCmL4ZLM25q+zu/dbx3ZlAkWK04U56BlJvlDs98rLsK
8X+n59riXml55/27uYQPaHfvDeQHDkYVFRzYqjvZi1RiCLjsq/GJsNUrPHUNoV2e5J1q/hdd/fzG
e4beNjYgRp244b3xRTwiuov003zsxb7U2BUlBKY75I+94C3MizuDCBLqEQfXd24lDhC8xyuOT7cA
GfWqHxZ/Uvb1bZ5+p151H3La9JvqsYSq2K6AbgId5Zed92OTSnBkZvoNqjfBRzfpNiIUPnGP1Xth
nw/mUUN7JXXrYUFe4lcvw7eYDM06nWx3jEjJbT3swRM1fkAhUSL6naY94Vu5Cbg7mSQ/rHE95w1y
fSrYKoHRykBEo04FKKxurRmVI1E8xIosRee+zyzeJozTjg+Gv5wQ86pRKfvy8GTbsLzxfXYMaNrl
RmaUqNr+fbO4sL+5MmnJX/qXwUCad3G+9XbZA45g/RkeJ9Zw2RMz1SwGbxga0ZcdLak1b6uCSJIj
+HTBGU7Z07i+HwBSPc+qhK+kaY+G/oX/n4rUmRrZ3UYMgwK3Lz6no02YknSaptNxH8M9cBwibsY6
lDMMAgsuPjXiB9sCja5Sn9HdU/i2lzWw0tFz/V9xABMJcvjcAYZu0eyHoUkj5dJ7CepI4G4dFWig
Ol3Ez8N5z3wFCzhJg7XkfrqsJcUpVMQbGA8g0OKrulQ8Loyx50PIQr/pwPeCqfyoMOustqbJpGe+
IHtivIeRh9vN5GC4A1NVHokAsWFbS1nIYxLcDkeQGJg8e+OdZF/uY3JhKWLiuWqyex7rXBO657XZ
d1m0zM0QIdp/JiwejvU6PU0jJZATBf9ZfaxauGHDJ/eWgYKdB7W2UWx2GV7pMFnRPjbMZgl11DEG
PQLw2aFvyvsAB9LdbfwhHd5kHOSfYa6AKvmy10dI/PVpQ6M3TjTVKU3HsRsHIrTUrqoJVBqGKuV/
CyN0p2W69q8F62asj0PO5YuvjS1wqKQ6GxCISlFYLqv4SsI0kcRF7KZrUKhPb55eNFhUIWvryi4D
EmpxGOhRmf8mXj++8faRJhXj+R1UORa6V7gePGFx3EAQZnqw15zkVY41c+vFiD3J8bJSF8+TWenS
WKPMh17t/zgfXIA5ITiW2GyFgE+E0QPA5boolyn9c0rpjofjC4JwTq9A17iDokqOE4UtX/a2ZD2J
Yvl9bdBLhAUggL9206J/l6bokyCfQUg2lanNgAlRfh+uL3ETlGjTXCc2dL8R6JtHsVikTuYDJfKV
wNdzcAivb8h+jzK/aGiEPkJCf4YbHye+UGzVkhMjUjEaCyWGBBmrdJ4SR3MjmIOyYC2x1VozVotm
2i6jtkUE8YeYeORjo0K/TfsbGgDNHAdgBISAdae6unjx1ZyU3VQVMEm5xvIOWuPd3/4KsNeTP+4v
eQX6bLZBt5YMJGInAtYxCNxyADvF2XIVn+lAIVbmv2Jc6TTHqNHkFd1j6SIUAknCaoT2bM5g7AiN
fGaoOIJq/X6e5amJeL8EENbZGjnSQtoQLHF/o+voFhh2h72LydpuOMXP9jrScpECYpFyOGXUmEL9
4qGNA+waUbpTtzGoiPV/bcXqm3jsZCOKL+1XrIjZ3M/hcmGK7ZOgGn3oOGGCcZwsNRvH0IDVFzNS
pjR6gibjyASEgCzcoyNVaTlus1zYN6oKmdU1a2pwrnIZcJ4+zmKA3zhNZSwynrEtJcWVKqbdmK9K
+J70xI3b1zhUEBksz1hpX/kyKxcsnYQYoI3EPbwGi24HiHnThy5281qC6yjoPfJ0ATF1GG/Z90QZ
j9HdO/LKEum0HvEoQCrY1o60wN18V/F3xMHwODDhopA49gA8FCzvfk9j6OcXa8DRI/vlsSatK1uy
O6EWbnwpStpiFe3ieB+6cg7vtuMmGeMaT0xRiatiJgtxhWg94MJ2F4adSxZG68hu9i3aEkttQPVL
LxyAckhhMenX1EDev8uIzxLlKWl7V7AW3Zwjnb8dmbMJmRXgdaQu/VRwasIClaAPOZtff4qt53M+
X91+Kz46IMDDFswYKmuGavxnvfLnl1LoGbQDAKy3VeXv3yB8j504Um00CTbOHvYNqgZBsMfYMa5J
5D/YOBCxs9e57v1FDfINuxIHmkDja0EkCw7d3Kir9qDJdtdXxCq7QS+MSi/C8hXpFMF0jJTgbU8P
nqH7NjB9cSEUEbUM1I7NmvlCRIk7vicoCrmWZGP/S3f4dwhivdWxIFYFUKtN45jwOjeU9okuXR1K
5lwhTlu9JFNHOPi6EDlYvQvNd76IeA95LQ5/zAHRXq5TKEPe5K0JO/L5dn0NrETgmw5v9Y5hX+on
OEv0CKo6v0V9jWE5EUgDagvmDH7mV1MzXe1ro07bjYVrERZCF0Tz8a3DaX2RR/LQBCPPDmv8KuJL
aFmwStr9g8gMCrJg8Y51Z4BQlm7OSNTfsC/YSCcuoYEbIhyx1VeJDWOs+HzHsJCQdL8T0j1lLCzO
UbqHO28n43rQ0tvEG7pKq947uHYKM8zsNdosLBFEsAgyrDJqJTKUiItl4MfDvAqpkUfyo4kJKp7A
IyzAj8ejz/tOoxKy9VXL4ayUWOUdQHmZMkBhnRVvpjhqn6Yfsl/4KUBCmw+25uQMy6LdPvYJTwpW
Tj2T0Aq+jRALpRRKIJ3HIWzgFn9P5lmm5cCTrGiEnX5cRvNc9HhXOzouxAV2Ute9uhTZEEgOczsn
FLOETHY8WGOGDHTNVnwohDhNtG8hpsb+Du3ANho6HG/U0CLhuqeoTcMCa9SO9zJneihPjF7SCm5Q
AbhfQRUsMrPx80xRU6tUa2gHvZueSH4bpRQ6E6iCFS84rUAvQWc5CwMtsQgiKizFRI1Udo1EyAD0
UDqPp3bSnR3zwFjyTU64s6a5Y8Kc0mTDk/I6d1NsT16P8qHWx6ZiMF7X/oNOIbESza19ACnMV02g
/+wf3IeCm1M28MHskxIXlvnt7WGyiz9P/sdXN1qc4Kp4rkCEnC2OMS7viF5OJrvhDqfAgBx/s0zT
HLzSraCK4enH3hQVORi8w7vRJhtyt0wKyJxT/5n4iKFYgv58Vav15Ks4kKKCO9zl/dJJvzF/WQmM
4WOEQktAcFbYDfqVl2irDA+yujGi17hN+M2ZrP4wV1DdEWA5K8V2BlWQNQnFihqSXRsx261TNyv1
N2de3/bhDWZUSmYC5jqhZwwJZn4BYDQd9P2gv82uVRy3GRCOhuHHvA3x+e7qBwJEgKveZAvp+KNQ
5MhBNW8p/KHT/cG8Hqiz97yFtoZahZ4YFQupnOVHBs9zIeXrZiyhjGAzLnpqnWr4AgO4NRTXZvRH
Ad3QhkQ/nNxp5dU/w3Usye2cSbMtUjKgoTAxLgQyP+csWD8lhoEFoZM7IO7Dxo46SI8AmT79Hu+I
9may3twceFxB+jADlsz84DQETbxm05RHQC9kahU269ozBR8utapznl/3J4T63JQUgzY+6GjSSYnQ
OZze1GRQoNSVhZjNIo3CdY/DgepVl3Ci3d/Pcm2z4iz4xsxxO3sHQ73BE8MOaAFiLOjBLissLXaF
KEy56vDypU/YtkQsd8pZaOM/b2yYoAb2O8yhCqyFKENrplMQbHo7o64i5jnbzhWiSvOhfoydviui
glGtTASQpyTCidPP6Rcsz7aaT8GLk82tbYDXa01nOk6CId9l1WTjzg3efqqimeugbvi+TelIe6nZ
FckmG5gIizPhEdtI6modBS15icio0Y/bORlNfmWJ04DPjaKPHMcC1Rpf+xYeOmkTbuvzkrB0X9cL
yN7WvPeuc2GHA8Prdpv7CXdgGopFxBeDMgKsOlF2akbYk1wMwQFjilK8oMq8q3b6UIzm2EmbWixi
iWAbeUUHkE1aCHd21KdoTjnB+3IPg9RAHRCh3sX5bUEg4NWzOeRdYXkmoVnFKK9ZGYgBnWbEZlGN
+urNoVuF2qSw08VKwWX3lYXpfCn3y70sdJH/5XG9bfpLqaKko7/m/EVYpQRZfoegCNaUTRdFoPKk
MWyN9mrALsMvBRHqHdAnzZZcIPNKpadLffLGJrtCEU+Po08NIMs0S8s3OuGtyfix8ELiGX75fHMo
c3r7FDH71FWYXVALZye/rQTwEjV8JEa/utb4VmfD1vCKvmdKh45eVSI7OAjIZ5NSs75rg9dpdWCZ
FiV6/kiUDBw7/Q10Ig5jqX7jMC/b0zsyTUxbuxgVxZ2O0oZVYRRc8BkmQHlk77wuSIm37991pN8P
OGGN1S+/x7bindiOmVyPiBXCzSU4w0XUc7Ibfv5iLKkrQRJWtqp5kCtZipbC5U4Ay3jwRAk3lvRH
yBa1am0A2a4H5IBwel9OLTC4oASvTxbl5bZ7uax9E15OzBivStg5OReonNwlL8z/RzHOzJVJH217
SWZXP56WzkKYB9RarIXEJmL4MmMV3IU50UyOjpHPMRHf4beHUl4Ho7LwebIMOsKjMibR2ADfkfxh
Ax+xHVz5yFUHx29ji+IJ4wpYRdx3sYxpA4MAHJ9krrFcMSQWJbCcbZqPJJleQVfGkOTDlBpC1P/H
GbgGytNAVi/pEfNnk6LwjAe0C/VKzhcrYj+aocc73iO4jN5/L/zA95No17RQrpn8SS00CJlMBOMT
uSKA7+i5SjwrnBgoWZcmGNqELg0Ft+97pnDcXV7U/yLYNs3WzNeY+mNEbOLzjOicnuAHrKP0W1Bh
UkPlc0G0I9nEOkmvoTzU2mY4h/d500gx7uayfY8/H9yaLLXw5c8wlvylzhbl9f+XQ6Q3YfxhvyNX
vllP9bfx0WNNMGkeL9mojDI2nLUIRHLKHZfm8P8HWniNJqWms9kYPWX2X/S5JCDumSt4l5fIW+Ue
zTw7va1FyBO08lzjWBKEUERQlTCNbcnyI5C8i+36YGhHK95qn7FTq8LOYFhBCRGMQ9dw3jTWAPhg
o/TMl3hKslIbdjDmSlloEzHheK4EzUcszalz9RRDGpYyRchk6m+dnAZYLEeRS7Wc+sedkHGDZnXD
9VPd1IUGm0WlMUFCsPsYpJs6GpAJrOrSoGjqWhOCqLv/NWc3bl6Ul9jYWOTnZPsg6A6/d/ZcXFn+
Nst69i76f5lRQDeNd6/JeJwCkxuTHlBMVc9Icno/UPyDAsNIi1HjnvEY0AewWS2SZFt/d+UAbqgA
q7GIsg9swE81VMpZsX2JASRcNCADhBImDnJVc6LoEkSOzeu16lhKsZ6tqzl+oBxX9fNfe4DtjS9o
NBYB911X/AnvOHyOOVTcWPM2gg5tM43GvySSJG4omu1Sfd0vmHAPshrpuV58lNgAKD/5fOogB9sO
OAWzjdR3WLuy/1X0HmdEbWM938o4IhnrCa7XL4bkaXWuo0vP9DntT9Y0bGw3KXh2EQEjgD18xgtf
6QnUCb/+8/0xqvm6TGsyRqh7VvyVxo6i8HFtjIqjBRi2auZAuYquTcC4fFxHupkiOyFPrxQ+TY+j
hRwP+dOYLb1p8gUSzneqS467UU7LRY8lR/OCYQTvVTJxSd1VVkyqbZPcre8CKQvO5krPkmLdNYlN
qBfCopXIyhMua+HmL4LwWctv/Ah6DEM+ri64jfLFvfvU0pe92xFLkcUv5/ZnuV0dMg+rl6/INp62
3ThYPjOU/brBp5YhxPsKLqe7w5E84UyCtILkmmd0R04RssEmtTHalkBN9appD2/Hb1YH3RpH8Z44
56iry7sWN0d5rzM2wCcIkDRErQMdByPRER7z6TdU9UDOXWztS2u/hnWn0zzM7jaDuaMAaLXBo0nx
F9TQqjwD4wULG/ovbgjVH/oyhxwshjOe5Ccajy0GDiav9qrHgZnrDxmauGyypi2cmqfZfOiNEuwZ
ZvBnSgigpeQIHZT17Zf/ew+iZM9sGIQ0CKWS0db8lJcR0u6NlAUobmp+FBZmWLxAknT6X8bTmLx/
y+7Kue2b1Kk7azy8rp2pUW8wCa1xnns/xI1aK2n2V+qCWXoP/W/3vYcXiG+P6HjkqzX13njydUcP
7MKNoO4yxomvFZd1Sq7zre95DTWu00McBTGRme4QXvh7PdqYnobnCOOB8Bvj2hUFR1XCyGkDqpam
PNOx3E8MjMLbYfZfEzmfv575uTr4Iqtd9GhD5FGwShhRzdvK3+MuIuMC2xd9/YlqobccsJ3b0VRA
oY5mUZWwj49JusPCmQ7/uvG25n01TrLjll4jozrw+1aqxs/NuiWoCQzjfouhkS170FDy+0UIxvEN
T9a0TCGQ6ffwJ05kBmTDEcCM66gVREA69LrXlVq+LHDAYMBw5Si2NXg1g3rycdz8yrMG8oy+MmD4
RZ6l3ai/LwQKjs+ecQ56SYyuFq9fGcbIj+slVBW/SUDUeaOZApssvPbEctFmzH51IdKeRl/OPJvK
l1HwujoyZNCCeFS6BtPL1GL6ZKQ1WbYT4eKINWP3kyy+XpDirN3GaA5Geu2UEw3jgIw2Xa/o400l
J+xOETWNaDfAPDjIuVMsb5l/yCtsDPBF9YxczXocEsQZHev3GwEGKvPrtkNQTCrO88+13DzmOEtW
aYeZxOB9fC0GJ0/JbjkDM6mMu7M4fsZTm4fEP72qRFIAGXL2/vRXhhmCoIlYufd3/ilT+1NoEutR
a08daUO32qwcbv8KgIm1Mtk4Lw/xEzej0iD4bTc4ksEZKvnYfzzYCbFtgFciMwtcC7DtU4U/4FqN
iC5P9f8cpPU4ittH7apd8XaoF6PCRmh2ubccXVVNLMmXw212V/J1SNqSs8Squs5umFhrd3wCGZpv
Hz/x6xWmonAaeHcao3/CrNR1+6PBLtt9VKmyYZpzFTeReErK01KxgbF0GJhyBzDGEe7yP14x8cpi
jkU+4wnInlvbT5xReCdCStc9M1IY5u9F0HgYouw7j0ySZ0CSc0BU1O/tkvnfRLxfwIU7IAHAwGsb
pHETXFfAdu5sgMwmFqd2hqaf3osidR1lrkDv0jd/rKTlwbxbXGzzrAialSqUZBlJk8/TLjjHvmi1
2TcjVUNrWrMxPacFJBvVly8vR3pnLeDIkgVclp+ytKFnUfwwER16XSi2W1gfDGIBnMU25GL1wV8J
2BcO8YplmR+sc8dqxdzV+2T3k3st4LFu/6pujyGVk+zMqTophwkHRbg6u+83BhVnnL3byX9f7qzG
updEZiyla4mflxYSq+kPZzkrPRfm/G5bFGkXV5zeyl5pw8ptvcBeZeifGeY7JARizMCuTt0rQfl5
ThKl53g/dBEX8+EInZqrRlshXC95lgs5FBinDYXbGDUSfqzteldP1u1WeVd0NJAOvnBTGLvGqP1F
iYNrSVtgZ8d+97ylCOyVgVHSnxQ7egVQTvpSSoa265FEIdQh1ckqeM13Gifv8d8ykIMWMUONHWFZ
ShkYagqOChdNS0tQ/djdBiTrCRy7v5WrLB0V3TpZHsMZ8RkPslMEvmfQtcR98Jbx5QWSQGLnCeCw
+WJocXU4QSTpcmWW5aIrcvaS4npprKzz6c/u2WA6g9TINV195BvNu4sHaEw8Rt3PfMf6e3dyuF9V
Td8cxPbVZb2RJ9TKdVAJCm8lSXIEX0ybeHiugjrtp/jEc1OV00uaX1zAEh1/xjUOGVuz/NHlZMbM
0azW8bwjdsCGL+t++ThWoHToej3y9ta9uQAJoHJ9YXjfrGx2OvsX2AoGSqC3f8/Bww1StPE74rIC
HjmIMhxloOtWAyfPFCnQfLvtygWCLqJ3W+Dck6nE3GJYYFWXrOsqf6sr5wpTf1+xlwQTay36Na0Y
KvOoNZO5oT1Kipz/6rXjhxop3lAmA1xrdOwvhR0xUddsf39KoPB86WZltox32g1Q9gTmPAS0veHN
9GKirtNNy79MisjtUOj7vBn7jntDeEYCRIJ5aAe9Kd5RFBqE/j+oaZgKVsZi8Mp/xwUikBbC1nIB
EK2Mu1hXQyxDkxDRt+eflQ438uU+Tsp7Ofg8+IjEA5L6TymykGaXAk0uhPzgPFWCMZD84ux7tra8
WsBV4UajbzSL59jGcR39l5kk6/9xUwGGRZe3j7PD+WriFlZmsIsl2eRNvYelGHkug8ffmK9Bp+co
SY6OigyDJOqqNccMsHWNNu/QUdsd7XTh55nnowTkK3VQzxAPQcgXV/hxsytYuh2xCGYT3Cfdn/X3
w4tK2lnTMOEGFjwM6kniirwx4+cUW+QKP0nMDO8rFw/+zuvBdmxoqp+0E6qOjGmnChwr6EHJWXm4
vWTkrO5bqvKAAN9W5ujD9umFIKHrSUqoOk8bqbC0GmvtPOEm9PskGWQncerkCu6SyHwtoGjbwmpP
U4Cmx2ShLrtPXu6zCt7DJE3KxVSqfXJeX/Xu8yqzPIjN5CcbLpIGaSncr9ZNNbDcIL+UGZGWxjk3
DDQznqHLk3oZN+TewaSGeLSDpIYqPIoWRee1OnJOxIjz+eJhSnryoH4zj2LrUAPLzuP2x1HlCU1L
5HNq6EscWDRzQHz2Z41EfniDiux/iE3906OTfP/ZJBjKTnubjyXQ0uamO/0VhSbEjjTQkv24g/f/
Q6Ii/Qr0H+mG0DOHcEtJC40fatsqqupy3aFkGHbwOs1oiDAm46gnegwxCs7OoQLtpL3RdppSG3/z
fdkLPaxcvghzGbCgE4PNAXR5qjChqBNIeJ/RUOvH7UVQLn9P/wQNaoVnDJHFJUEA2t3XZg55pPMG
if2OiEWxxs9zCmI7HKLGkovTvAZAHdm23s89hjyXZG2rBMO1mnM2zIaDSRVu9lg3SvH7L3pcjOIR
1InjK+JHsm2+IeJ0Qyvang4Ahvr23UG7oJ/kNdY09knLtsLoTlaIbXwa+NE23OrtU4VGbAfieh2U
aEBDSkC3HdXwVrJQNfIdpuY8eCTWkMEQcjlAi8P1fjd/EHjHZtUVhmmrxw/4O9+2nWsLpMym7hBG
Ln9cT28xqZ6cAIpMnuus0UgdSu8ISE8P07HKEAmTBcGCqiLPIrNeR7xv5L4WxvfrYcYi/ove66F2
kNIoFYM56c9OimLh9yT52hjbyLujYxiwRGLYy06ctG9w3dAy5qtQuuIBsAejxb5qIsGMvCG3oLXC
KSCHOOxF0caW7LvbUhhOoGOYRMEYUkrVWVjzyGiqlSzUECburFOYCcKbEvR3UUBbJ7D33GdR4kFy
opqL74e3ra5jaqHh+CJyX8EeHF/i7S6SjPFdih2Ir90rT7sKCnkvKUmeYWDwQXqNnV1T0GL70Xw5
aEa+/KGS/FF/5iyygTaX73u17L8ePB5ca2jTEeofptbRuRzRRcFxif8Z9hFar/rRrC2IUHn0M0Hi
t14uu4ET8hCnuJSMRa4PlAc3dRGce9VrfZkMHsfk34i4Bt0ClzQ0ai9+xhcru5xEXYOFdmr9LhGc
/GFinXt+kR8ITbIFVDAsB9EZk+vNLC06UMhuZjDFMbcMNfD6SbhK6MPmIDsBc9vPVZok2WRRWuoY
2J16CX/PwcXsXo1mGIufAZzQogbrPTdAvlHlHQO2Gix2wJlrsIS5evWadzF7JLHv2OUGc5b2VT3S
CDHTegoPhtM/Xvax/YHtNZOgAIEg5w+8/K8jYIgOGV3rxYuQYtzCZI3ULZI2GTGYsFNuFvlPwZiP
mp/j/kykgK0L/5JKIf2Tu6ZMDvMpgj/27TAQlq105GAp9XjSZ9YcTILW1udl50rQ2E8NTrZ+8Mfp
v7DNM9WUjAEQiXTE0UHxMfu9+EKBpu3qGmnidFJL7khIPiJBlu2An5YQW6vAfImsi2Eu+YsNALiB
iKw4wo2GtV/MSKebsMJlWF4Xp8Mh+oIrBcIDlhJBNproBAMpR0ZUvN473368qwp15D8OBXAXWcvw
XEeyWW9ocMeVnhUjrf8u61f3Vttk0kTx7XUQ5OLlQ5TnE/FKz6A0UfwZiFI9JygxO1EQen8vU5rh
MJQeXhEK+lEmspMow3Mz5voPwYeexLd17u6IYvh9Zqm9Wd3dX4CyEVglMSHJZSJT8gEdn6X4hKqw
Qot93v3fQGevvNZnbUwMn09d2Hn3UHuqtAX74ahVhCNr2aUR+RFTPxQcLoKYP+loOQvqMt4rmZEw
116cyhbWEDuRWqq3cI0nh/yqXArn84N0ou4qovA+lYGIaQ1lvpCTTQ6ZiHs6m6qALR2o0+2/1IAr
iGKOwak5enctuOggPiMGL59iowxhpVyM5/ywTH1CeM3EfdXVE3Y1tIjsULZY6OHImurFFddh4Zc5
FEMsduUNK5lFYrs0oaoM3twlabvqOy5O6PeUN+P783qnNJ7lNxnSr/ZNc2hbQZZsHlnjFNW0CsHf
CRlBkSl+irbH+Ed/EqVs4ypgVya2EzPN0LZn80FAwuUUMLRceaWhm36fMBJRlj2KOzpdMHjY1Mab
WHLGPkm7ruaHIVjp40qDSe7ZExCZH/gzhEccMEsUdLu5+dklnVuqYkdE/oF62z2zdwB45Cx2hQDE
LMd6wHmDjFvm4Om8FTPiE+ePYUynSN/1AjQxP4pVPyo2X4HNOW9QKpVB9hKMphxtVscyfDWLE68d
u9qHEJ/9CkckJZL/mAM5pcWq9PG5ztxLPQypcT09V/c1FG5bfP/LjTm8VEsX6gaqJ25m1rnbCUXa
TSCvIGv/LjH6CTzoZbJUPfUvI7gKRjYkrj5pg7tR4y7VSXc4DiF4J43F42bau94ilKhWK8bA+ErH
V9ZrXShFYyOQMilXArkqmKj41IxNDX+It1liPBqE0DhGZQ02L2wZ3yX1aafcXYuYQijCs+mgY3V9
HZtKvpWphwPswD/E4EDnmrhKyqEMffNYFmY8j8tnbhcGUVVNPpJ8SROmjt6g8xyd3MY3O3GRQ62d
jyV1dn7jHNUgmchAkOWqeYWE5uZvr/VzVtY56AMjCq02sck/OFQyAnVkGJCC+2hsoAx9JdQnO53B
p0PsbfAwDnya25PnvVQoCC53XpRqqOpoQJsoFPkhtFuyE9yjPary5pmif+1xIfUhOfqCBS80nb5U
95aCMC2ID8G1QhiXoC7q+D2kJ95E9hPWIVCtjGT1ZizRBIs++NT6b6xjBAF1n3lUkHLFMTLN/Wvf
sHJIOYzeSbTi9x/xVijs/thMI3hLYWL+L2jA/gRVwjYmhPHOCUj6kpdTn7v0oF9nVqtAbzm1nGC6
wnUAckJUB15IhPPYr9qefnrpaVMVEireNeh3uFwfj5VyDu4I1TYtoaX2FiYGx3SqUDpubMImNR3F
psAPkcL52kQhpmqMqxw76vWCzCv0cc86LGB/GORVCzEDxkLSwF+a+g5GXnkYbaKbPwhGlKFMZuIZ
D9X/VNi77Eyvp5L95qnJfEw7CK+aho3gO4ut3a7t8v8ufTDu5HIiXe/EYEpQ5bJ81tdtcCb2Yc9Y
GcG8dDFQ8ycGhlf077z6loFJpa9985kB7/FZOx3oVSZrJChOyrrVDizBXHhXpwSn14WX5+ip6y0R
POGr+z4dKSNYemuxEllvy0GdHlxDfhUqgL7HOTvPRPyE6sO8Dp82lSnZLpevRi/bYJfb6E6niduG
0Nkf5aMRLFe4sXw0P+IQa+WGl+bEJlSwEZDv+FROFQ6jlvIJCJ2uwu7GU4jh4zmaHVCNdXXvem8L
tlDgfE1ANBg1GeQgOjmF4du+Jr1h6McfWFBq4/mkzsCB4oi7n1/LC0j2E9/OQ7CVpVykMsE1oqiM
1jU+nTVCBkMesHQC0Uvyqo1R09R4w56bk03DgxDKpb9OuyiW+x87ynwDF4HgPso4IMSNlXwHmlLx
/kSPOtiLhcbrThIO7eIaQ4wQC2+ooYd4WH1Zw2Bt6ScEOZwRkj5mw9gX9CvqX3pkpEsyJyWYhkmW
GVmb1/1ntdDtReBATWy4S7gL58Vjrx7yuESKNtlgOPjf+u4BI1kFb/waDaSE2e+VNa3pjYlQZl+Y
dPAWBu3QCqTHhBvdiW4/eph2Y5SuqjxL15VT4T079dk2DNvByYPPVVLy/2as6nSsi7pDaKd9jT9K
SKrKCRsiMcX5zzN70YpsSsa+67kMENjjec6ziz8nIE+cbI/khD+b68tHYMhcxRpwFP0evxm3DzOq
FDu0zwFC1mCBXvBpOrKbKbVFYWSNs4Q8m6ZzARrQdmJnCG0fSP/GaU6I/JLy0pXJXNO/jLnc0nBO
CshAWIxZOVhNUvRGBofBNEC9InQqeNEy6m0BSGcP98wgnvL0I3s2EIEN6pjGF13iHldgg9x9CvYT
vyWicn+y91EtQSkBBBBQXepxpVphEqumzRphr18X51CrEe+mumb5YogbdZE8YCXsouDC6VeZPtze
lPX/o0UncmUVutjERfdWFdZwbC3aebxSPg2jchcXffDu4cOHYn1e8W9K1AoKt9pefaQkljONDOEC
21qGWY89QDHVhwN88RYTjXmeGgaOlJQ6qF55xk5xaSjDA/O51VvSUXmNNZ/Q788OmOP4hv2TH825
dE092BDjLBXA/pMPKzhJ44bzTKXt1slSRuR0ewuBCT7wLHL8b2c4sGwnbWRKOYb2OtLv6y5iwOTn
foLsYYFke1l2vl6iHSbuzzjvZa4TUz9MkIfpjiM83QDRGdg40BrTnwM1/mYx8L4NWqw7FbR51lr1
s40UNh14zx1PIF9eYMac8EFYnPqXvPMl9pEqBY9YNCL2pQ/gxSLRBgFNbsSvotbg3o7pXK416mqb
SJBRyyLnjF4WwdSMFP4kGvNzpaQi1OMg1wm/m8akuIxMWrMU+y2ghAPTLdhodY8epswjleulbZcS
1t5xE4mMV/gykqRaG0fY1tBBtOYZ/NVR3CXPbEvsAxERYLkZI7BamObkAjTtVjRYklcp9kJQt5UR
amw8U2Xk1AySx1qI+Yx+2bIQcjHG6+tNtgHPGuYWTQbhLXofQGqSj/RhuQ/SFAlxjk9fwPEXmF14
1HfMxiHni4WaIK0wzNwqLFAfSPAIy7suCki6i9pqshgWxCa+cByrulNDkipDuLervXJSq9sQHXyi
x/xbA8fAEgaVIPvrPLGV4UEBcxy83oy4WOH6e4zT0iGKAhQ9KPjH0AphXJW8zt/ae5TrfwmttaNX
P0xF851fgZk8jn+6nG2Kd7+qZstjW/YDsg40tR/ZHRjV1PrUW/EP1IVA2rpmh3ISBpDth0nLzYws
naD6tXMTLS8UiK5a4+e/ZuOc5mxzhWV6624/sPWfbI0b4qNaOQ06UqFzLODg6Y5OKd2Wa1YJT6jI
+DMLzkR02oPjpL2tODK4HeFnukcUfeO3/p2IFOcPHXiv7wzSf99awehm1vvqj/IvOWTH4iL8024g
d4hLbZ1xekXCphlNnUkHJCLYzfCnZ9x5WiS7QO7knqEQ1wVSBmKLZpgHwOTzMQ0JrABaRTlSHwZz
Y9kvq1b1oJRE1ZsgDjxED19cLOUIvrSolYfz70jnvR2JupvP7SgRrj5kGUPyEloBjD1RS9nQx4L5
qFnRC7R3D+nl3t0hfYbXyLK6569oscVEShiPAIQ1npvcZIUC/fginJD9f4ssgceC3wrsMV7mkgJR
Q2q4vfv3vxPbnvMivfAfvkANyHJHehnAg5g2N8ZOrlv/Cu5GlW3iYkMWnxR23AaxNczeE0kdrmh0
VdEkhexo+F2T52DgM1pqTOSKLjjIJHqY4QAvppoAkT7Doa7Bv2aKQNEjbZEYT2y5CGVxZSyCOMQH
AM/uRcwI3WKAvmnMxhc3PRCj2lCFPR+DUqDWx5TCWbFcaT8YvEy7pG5EEelW6v0baaT8LFWz27z0
adDpDLO/muYa7d2eTaxV0P51L64AK8tn3YWVIXHQ7cpRBD6Ztx5Giq/6tZiMbfL6x09EeIDKcIHm
HM0ADNuTylIDMkMQiRaQQ+Zj6lEaMQjPjR095sRbw7q79pC7v/1aTtYP8RkwWTiInoSlZZupVohH
GmR8qW5DnT5+RiwICb+oNZGcv+Ru2EQ5hW7ZVqwQd1Y29WsfVNZFB395Dh/73eSiC317Rur2+HRO
a3R4v4a2uFxU/k/Gp6Aax+ZbKs5BXGgCzXyBRGwEXxc5NmJn7K1Z4vHd6BQnmXbtg7qg1Ib/Hjuq
6XPb2wY2KhnjzNGj0iuLslPu8QcYBZuMq+9nXOStFAPERIncgKdUOvPHSReuAZR9ldTmEiTRGoMf
AT/OwDzkDk9rZIzZqQEqeSw+tZfeIJLLR7+pNKipW+32ondhJse0NQsAfy1VLaV56U0xhszzepkt
ic3+mS3zX9fIToL3piYSrTBkO3KGIdpRk3nVnocXgq/btdJdMff3GsSxR9ISV30whTUh/ZugBRtM
B5tXpxtBoeA/RQCF1c2gPVaBULRIfxBcIxXTLhl2Zaz+NjuzrtprVHNjMiTYBh6m5UJgf7zE+m6c
nr72zZJs2YWYGw1/af1inalxL2mDJb7vO2pSjzyn7Z5sfH3EUPM/RVoSQUHOqZPjWEubvTJMEMwy
0GPa0DJGneSXYAZeMscY8wLJhClZFBet2ZRaBPgjkUg1KSlgMjEFvfW5zirnbRpaFdWapRFaKjjo
3D9+5VnYkX0YeZ8U/F+7rUl8B/E6mi6EdZl4Dp1XT5V8Tpfjsgf3OFq121Rrs49s2cit570zSUPj
CAzFdViVvR4f/0av3vH+gESoLYVvlipuwZ7k1J4w1kTJw+2E0IggwNDG0NQMXBIZuAR8xyd6WGG5
eWQG0e2NdcnK7WfXbs79tZEOXmtltcNU+EzHO09v+OMNXORBrtYM6m0xUbKxbnPGEZ8OAL+EUQf9
Z1kS/x8wdPqW35rtqu9IAE2Q9E2FHNg9ECRnyZ/W2WUXEvuJWInr6vnHeKV2dMoihREu4ErJ+M3Z
ksW1WjZOHCq5HLNhOdv9sDH7OPx9+iMjueCcumjeK+qqwQAOS+JPxRO1Eewu0dVOv+/b+A5n74Ay
szea5BZ98P0Pj5pEVgFIl8HVjahDmbQ5T5FmjhlyhnYnBb+yfhb+I7groMVGuTZ2gNoZjA62gjmE
vTJ/E2h0j7pgTt4GRUjs8K0AAVKOBRWjbEUcGRKG4JxkaaZgDm60+5CCzimnpXpmMF7K6FEbpGCk
4S/aNZSGv536WRWcfGcHbAx3ACVb7mFBlKb4bjRoQfxBjrrZ7nIH34nSMqKPx15fbNOY8wZuw7Dr
PPNxOCvVTQp1qKmohjQ7Fv0saxsk0k41pLqzQeYNkRssl99Jj/s9/7TxBFQ81WCz+UI2gklORoxy
uqG62rtfpbH/cz1ntwjoX7AyhD2c93zgQOHllyCEvRN/5P50MJ729Z5GyqOr6K1LKLq+GZCTIZ4S
3TFf3H3/t6R1itLXs1dV09alAN3790urNM4zuRxu7S6xEXhz0QZgMyNluantkbRgY5pkB+5CXvck
SrOTx+aazipgBUpUvEEEsTsHQVN06Fcc0zdIl9QIn/pSoez7z+/Z1S04KC+kSCJkU2AVMVHWU1iO
AE/+dUMbDJZXT7VM3TLgBvnS4bNAa3osWp05O4TG1cDyjwFU/1I0Cq3EfJAkIojsa0whim/aQtcR
agMBfWogIDiinMR0AlPpmlPEXaIqg6yvnCnPGAYjDAtPgOiMtGwVIJyKGdceYXt8R0QbjRPlRNm7
TBWSkgfHD0cB0XUI2Yn7kvML03pLPka3dSnGEraLB4JeFQzutV0P5m1FQGCyPx1f4RNwyM2z+ply
Sn7Q4Ro2/ShC2m+vQi+9AiFpr2f7Ftl7s06SRp+xDkRiOfKCzpiXqhQi9l1aN/VMJmXPRA1Y9aE8
kpQfNSDwW76nBaOufEwoK1LlnO5olOTuTaApzitIUlcRXIqqXt8kqV5cWwPeA1F127+wM37iii2V
K824Po8rktHOm1cMUfUqVL3GnwEGxZdMhPzz1qRK+3W1mDiJzqv5NeytaloME7HvzviL4cZwSUmY
BHxy6QJKJtLt2R2QsqOV0ODcrzq5TFr+YxqvqTUa3JpbpkfKAxTOo2c6ljxVfi9GXKV44iiaIida
aTcb8pkdmAxn02qxCTPS9YlZechG2y6UPGd85wVTIWqqbxDui/KfB9Pn3uCXr5ry1eg1XZor3HV8
9L7qnJAuzV2f8Wg3j/bJjt0BmOTqfXc+Att+QzcSK9zraOb0uL9FnXgexOXpqqevDRHBRmUswuWc
edX4nRn8AIEGc6zW1xQBOIyFBx9AtkcTBBDV9bzE+hvI//7bdTEfcQ9Rc8D2wUhTvv3xG+lwx1sI
gmtDB/AnZEk0oWZsilP8q7SbGI8RTA4zzOanMsd7lqsbCkk79tgtr67nONAdF9vDzcmyDr/tOjZO
vRG+z03ZHh+J+35HKKRet252gFuW34K8aKvJqohISVURtTfG3KRVleM/kLaEUZseel2ay6rEU8Iq
Di1qaPet41zh2gyu3hRFI8uYXIw5JQbqqWhisOK60sY+ycZsvz9/RlIGvZ+ptrnrSWYIYZ6JdNyG
mTazxiMayYLN1pa+oIQOkJTSUp+puoz8gou41aWXipwXkhqMdAz4CyaA6JXWU7NTzEayVOmcmLQB
+4MuFHLxLg5ShALMJ4sQGDodtD/cBjyqTZ1xlxSPV08se0XPejEHVIBLnb0Tpt1e+a2p3vTlIQbw
AM2HXN97g9VA4JNhitzCkku/zgkCur5b4CYvDKW85rLYZEdMvjvy0GrsMvuRfIDpHqcLR+zxWzuF
V77VWbsdLEODKE6+WOUz838W3mdq4yyf1LGNFEcSz06gmyD7slUWVKktSXDpieOrI1Zcmi3LbXax
dPjEIsaXmDjdePQa7erwtHq2OGqKO4pT8NF/YmX9hhwqcWbHIZnCmtnFzXnVgM16jljnAHQslOxK
eJieyLBuqvJJ3XF6b8J3rJia7MOK24Kba3V7/hBEznXGf37KM2kxq3V2qbufV7LESCe1qsABB1d5
9jj0i+RCdiUXMGdcptJiolUF98S06C4Ms64e2go2uxs6V5kdMRBAxcJDmTFWtXWK4gAwxrU6pIwO
5r/bOd0o4xaQecXiF+QIrmpsmu+8VRYSYdDKDxqUeSuyJD7TQ6qAdLa+xk5WwagnuzHooKKtKNeb
n2Xrte72IqSJM+bdX63TSFs8zFSZl4jC7+PRvWkANgU1AaElEkeypob18uXte8FgK6tsOhwzS5K1
83p30rYkS3dn7571zuSmLOmYPsYnwUVD+Ztkw83dIdsz/WW9ka90hCH4Y8wW9i9XwfQlnaexag7p
CHvf0snl7+2v9JU5bLLiL2a45mb0zdhtDe8Ks1pr1E49JaexkJTK/wLrUEqT4pWgHa9eDXLGY15u
V1G1W4q+AH21tApcDiNRPf4ewZuF5jGBV9dGvofLpXRKEwEetNgTsAccTi4VXxYQS6IVI8oo1+I2
K5zeJ+pRKmDcDv/z8SW52h3kD4YYcezm17bRlPKteeF2F9rPhHkhKYNSL80soCrD4cmb8P5pBLWh
c7DSdnPblgDtWCD5KQsoHB+Ny1OxLcVfU1xa83DiV4QFDoB1PsOom5BlLJEgxobe+TajKaYlpVn7
J1bNuoueeN4o3Mf3nywYoY5IYsi1Zok2BC9Rys3Hyj9Poi5Pf6sYhvQgapKVNtU0m9SL34pbz9Cm
a54BFc/MfEmDDi2j33yiayIHRXzmwBG08imIh0aiPocWXR/PiuFRlV33ts0LDHeVn8y0A3BT0+G9
echbnGVCiAV/b/4OCLEjtk2rRdkyKNvMRUbX8/JIsikztZd3RgBhI5BFSt+OheFuSh6XUiZvJXXa
quPuDoXRZVEjrGoP1dbI1rbEDIVx41yaki9HC62JQ0eWFKu+ZBX3s7csxZYadyKE8L5k1y1RfI8N
r2yQ74IlzgzN1AEVmVzoTn01bzkBcbChTrwWrsjGNO9GEQ/vaWM3Dr+ttmlaxfUf59VrNV817yr0
mFMtv3YW9CEFbehOFVUeMcUOMVFJV6q5KJ7ldhHeQXwDqMnDFF57H/28QPOJ3FenZIlizXHFjOJl
vA5rXktQUXH1zIfh+MerLJZNvhLqPMS0nG02w4WRKHwr00/HvFAK9isuD/TqCg3K6MWpiBUMHsNy
7JAT4ppZ7DvAXUjcgYxi16aiAxo1F+hjEz4MDeG5xgPvsfIDzsuSCo9EqoEtNiO0If26Xho3gUaD
JpIVwqDwyZ0CVGXomIdCCt3N9yaLAsVSdMjad2vHzJZhj8fcLGaA7shxIJEll1PCgFsISsOLQtLD
0jnMBunuQNXI13k2lWQnBOo7L9toGbgMJJp/+OzX3x1cdkppeA2RSiuMZCzTxzm2ygETM+ZO72CV
bTHpTXpiEmW9LIz+OOvGBhgiADuKOar15Ud0X0k7h5qTkSSu8CFOCoDJ3B/1koAd3nzLcoBQ5kCg
dU2kZNMoaQ+St3B4snFJkXhgVEuhkoTRnfIpWy3ydKi/I9GxufdmWb76rJyl/0pzDxZisu/sKmyu
FdP5WeKBgZhacYf6GEFTPf2sW/L17ylPz9dmsscCeNi5D2IK25/VTe8J3lQ5j+R6nuacfPjvTbt8
/HaLZ4HAKikbQwwCE/LhjpG2qy1ZYQipSm7LVS6Gb1yJH87rRq3Fty9Bu/gxQmOEe2M6IoNlH85L
usn+TasrXG0y8JpiH5Uobl489NiSnY4TjE7kzAJAuy+ZRZiNhsTJxu+Jqstid4OAO921MEucSpWQ
wYxM4uiSdTd4gHhpzY9qASTkkw+hbY3fID/9zdKSHOfIHFY/EZIf1UH47FiKojESXO94ODMCc3Y+
8Ztpc8oMHW2/OPRPL+YDzd0Mf8aseFfgZbS4I5AcwlfpRPLY+yY6NZzyy1Jl7EVNQFjXUJkhYZdO
O6im3eOkFomymf/iokdbASMqItNdbMVtkQl3dzzb/CvtrEcBhHRe3qMVndog3xaEVN9PFgr3/yhG
cdiqrk4sp6+/xFCUqm3s+loSvTH80EdXrbETFqO0xugm0c6h1r+RJRcVjaKrKT8BdjvYHfUcin+i
Qg/y5ajuZX/EVMDV4qVpGVslv4a9tqm1/14mmT7WTaJ7+RRr9v9ccuTV/zkT9u8WYsS6p3c7yR/q
ilZuI4txQA1PDbW4P3qKMVCTbxRGdRXQcoqEgmrAllt9Uq/wngKodHYDc7v1IU6/FgxPkx9Spcp/
wwoV4PBzCDPkm3ilfrej5YuibGEx+BVl4XeCR9NvAkr5mQBt6CUn5lwtATojt5TzTAnLCWz0TSDD
3lKJWyHzINwisNW2zD9Nrvuzbhsm7EiydcDGpII4O6Ss6obuFradTzx6QJsqQ1hoR0Fuh1gpLNYc
SpPVn+rxsi3yMxoJdelIpVRLAC9olpGat9R76onqiyQVLwImlmfIbcwpojE08w+PKOUWFKWcOi1P
nV6/Fz+ZZAtKCbcm6txr+r+iI7XVwUBes5A+Tm3ADz5iEHzRnwvkOa0HHocx18GP2ASs8ZKm5pq1
PYAX2FdXbCTCGQVWBxDKhYxoVt7PnwIQLq5S+kI11znYED8EI+l/fQmvZQo8FTICpd8pksmVl2TB
Biv8s/Rk5fAJUPfOqCI38T8y7v4Bk0egf5xQHcoB+VuZmhmYawS+MttM3RXoK38Qgmnw9f/fu8aA
LP9kMKkSDJWVJ5FyzakWxcXciTs58X+NNxAvrs6dJdk6ve6zupk3Cm0k5C/lJWHEo5VPqYBSU6Qh
oJz7zRONjBx+BC+ISSg2nveZr54RhgB56wuOpcGZdh0XFnMWZxg5twHUUcpRCRU50zwdM7s4Zcpq
Y69PpVk/pCmqOIuikQvrsysC4kFfYMbr9Xwnb2OH37lOjFnjEs1S9qcybEUEH04p3qdKm/u0BYRx
gZ+GcBAeOlOwqxpzilpb3k6G3sLX9vHyRHbmdqpy8/XkojfsspuwvS56GVoITSN549ifa99yiSmK
sEVahzDkf6O3htfhz7Qn2Pc3QPdvT+zfGwWBnlAHx9o0D+BOLp96S7f+pdZbNGOjtneRp31UKEFh
JIoDnEVQePeGKPsKVJPM4isJH++Ph6MeECtzKlK8YEr5nFZU7EzHHIbEx/bwpm83aUr8Zvbjkx0u
qltbFsQreC2bvVWFA659DXTyjM3XK6WS9ojRaXA4iSsFwpGZzwv+xw452CCmsiYK39a1h47idcWE
fWd3qrD4qvDwdai7x/TZPRgNggyamvdRZTaP1cR3l9D7lVb+LYE/prfApZ/WW8VZKOT85zOwa76I
g8hTLcOO/kLz8AjQNGOQ0qVgTzDQj0V/2gztZ2eL5UP38pMsC0iqJH+VWK0YPG8lMaxx3HRZJYQ1
Eayj9ZbXERAATHK8x86zSxVLL0KToPjt0ZxycNy1GHXt2Ccr/FyLrCshn3IAN8MKkPz8iQyq9Li5
NSIJgg0XFloR4autbM6MrKYwcmVOZaE8/t4+Mz0W1hXvyGKglUGTpRE9Q66IhFgQ8BC0BhcWYlG5
Z3Yyy7zppdFmFScX7aYwXif8mZ11qIk/WBdZrOVx94PdfYYfTLg3iHLIFxP7eJ2lniKNcVHqX5W2
mycpI3/lw173iCwvqnNEMuxibeQ5QIcOo0rEhsDVSiliyF0+vd1KRggxrfiRcjgTOZmFFlFv+4+h
Vh4c/qpgN1NddMXlylI4z5uRKUR011eZMBZ3jCamknfD9tqa/MFz6EXFsG8tU1vbpaMFbzOOjJW2
l/QFTswSbAEbN3pu+3otJTMTNvvNwwW4DsxF8Nyh81EAJ9xTg82ECWYJHn9aGfC2bjqfiQzYJ1cJ
n3T/GBGAATv14YcVlI7JrxbboJ3xmYQ03ot7TVwwFVqmm6Oi1/QhxXvMEngqngDo/kiBzL8gwBhC
IY9RsSFWyGxdbwtAlLq9qnDWc3oC2MHBnGc1xqlj5SO4fffb1awOS97O/aRxq+1IMjXsg2F5IZgm
sCHiwOiXNDlEIP6pNcf64s/ZUPR1riAlm9UGKImnP8dgpm9ZBhlcjew/k5cgYbx/sSKJ8w+VPGbz
70yZPUnTu0guGc1CcLpKaH5Yn6tAZBpCO/2xIY57x7xuERtO1Dclap/T6H5e9CYpuRKpAXs+s9jL
ecOYDzDrjSkt681M/BL9OLlidMqGfvNPj+dlOPv8zE/bUlJBSHlZDWlqZrNK4iv1Q2cJhsvDh6Qv
9juzccGTKEZT2rorNzFuZHsSVzmr7daWUdpTb0du6dgj/i6/AAzGq0yVWjls8K5Cj9G+2dywPW/8
Ez4srKKTtl/8dBg+7I8MaR+5pMhezLi06aYQNdXsBc/SswlkmndDJNYVVjHulnrliN7PBivMpc4h
x8olyBEr2YHOyz9kavGd906jlCmmREOMcE3TxXYKlgGEn4SrIx7Wio4VfJtnKezlrTMCZqAeBj+9
KXBqP5RLUl2if4SShI8FGSm90iiHE7Old/BZ7l3bTUyYGJTqPI8B7Tk1ZhO9EewcMQbZkzz288V3
5T6Vyi8s3UcPMswHYh8ovESg2typFmwa0DU1x2OL8KPb66bmaeiG+KUaqdUQGUVACtoHxUDuJVjj
4LDaOZWt8KFuk2zhR2ET6IbURZYqLlZsfayqeOPLqyfKiarS3cv7hrpAGqfTDs8JLVG6xLTUMWps
3guz0IIZBzpB35UUKXeysPcMPMImzG9+Kvcb601WgVy5u7zy5Pe5e0aM+kUMtRZ+wGm7xtDxyNxO
9HKvT1j7eSZCkBYGQGHfgEP4DHw3XRidjTqXy3M4orYe1oFcu4Fd4wVwKBRZLY+niJeBjZcWYqH9
G9eF67lJ4HIQYfg94P/xPEf3aYcbi+z3BtXRnedIMdC0mcFP16Pu8RTpb5a1TiD643/EbpzGn9NQ
WjP/qAS3E6h6sDjnQ5FKc1lmcHWZu6hXk+N852ZGkGP4eQlNgCm8UYwfnGuTRhfPuVreVZL8lOQn
GeI7h+BNYY956k+r23wHVrfOU3ssDji6sgIzf2UCOfr8ZT2LCx7gQ4jjnY9hqVaBgYYtY5iDj9LU
0J1gTJOBtCRfB6xwFCQwNY0khJwVA3dqDKd8f0zlWE0M5xS5mxeyQ+tPWc+hgfVpisy29p00sncU
cp19ECyhSiW/tWyaD5GYnd704bx61LY9Meq6ztcxW2cCsJOUZ7hsTZ3L0YQVC6+E2vYfYLKlga3R
YOHGeVeE73gmJShXg4oJu1o6QUZtvyKe40SXpfTsZj/2/nb25pUqpcjLXvfFuuqJgYdWEeY3PjiC
cD72TjRxlGm3YX06HcLp0DewqNgn8Ayf7vu2UU2lpQFANovRiv5uPryUts2De+qs47dsV+25aWYE
yGK33P8PZB/4ok5zOfeED6wi+ztQPlMt1sa1UcnAAk9vlnVzpmycvueYE7mvms0mtG+o8DkdIwIJ
9SmQO82Fj85zFZT6wxTmhls/W9JZyAegBOGQfYXspZBQuTV04muSDYSBoHT4Tr67YwlLd1Vs0A+R
L/A8kaKU9BN9qszS9lUnBUVRibcuYUKHgiVGgoqBcN7FRxPbNkMp62RuOYvVLcvTk6fkhGce6jdZ
y5l+46tcN/txzBtA5Lho/PhSt+srKKjgqOploejIpIXo7CLgNmHqQDFU2X7QYYgCHML5To80WEMC
re2LfTJ/CGlTyGr8dIY13eJVofhLXgoQc9AAEUCPVIXmIsOAlBeqnz7QhpwF2hXLQTrj2kiywI8q
muIH+0xGoFXQEMImZc44NcyxnuE3jXHnhWul/v9X7xPYqL8kxlnqT6ifpddC2du2OBIHzwByzmOZ
jEjtseb/RyProib9/yIkzSKebBvDopvGrtYdqjlawIGyYdUXOUKd7YeCCBKXuLveJiWD3k9xTH3M
BodQZ7S157icsmqgwSyo2SgMbQBnSNAMG/XlYa9ok8SxwellQxwg1NrcpB0PKLjkpx3LspjfWGVc
gvOIlpqd8rQEAZGisRXnMjfYFuYGtnzX/1/+4jY7R1Wkd3sOiZJP/hCpKjbq+UjrYd77UR25Tvaf
YHN1ajuCcK7wuKELuMOug9I/JS/O8s38WM6TRfD3zvjtdodeTPT1yvP/AK+bSpAiw2aMK9os0feb
j/jqmuWpyb8TkEVjK2tDDxB7ugIH0SofeqL1XcA5MbPtRZiX4nfpeUTw3U0UMqSw2KaJNloAJYMF
6B9tbX18w0tc4U/QNY/oSzMEc86g9FWvAgW5P4R0MqUswqB/YxvYbOs1V8Y7LOE2zgZCf1+N5q2K
z9O+Qz3snc/ZiYIpXKB+KMqcYduP8eMVLUE9N5PN4Jel10vLRA59pHAr6p/eWlIjDXKAdQ4fYClZ
zr78cT45MsIHv2PNfU7pC7E/9i+mvCqOULvUZL5y3KPCZsH8s8OIktSYYlJb2zNzkjZMYyegWHV0
t+cP/sgK35sDENph1smpUQXvXsNV7ltWL60TLcgauv4u73Ku927LWL3Ab7nAKdEysau5aWs0r0Gc
fH6MKR24nMoqfQ2ITk7PuWiwJ8bWWmHMIroQgl6TxJjcS8fbzNOYAdmTKFpiU1U8lYCptF+CzdAl
tIdZ7LxMlKqYt/W2BNUEmtkepv5MryZSWJi1JGBV1W6O4X9x8iHCTVdzktI9lRgpEwpF3Hmjysw2
P5ApItbs7wA97pDBFq2+FvyW821rqG6pR2kxQInuGuV3Hh26D0ucqCmgoO0NxCJHbnLl1+QvLS6g
ivaMcZlbq5YcBFpxuOl13wG1FGY/N05mXBwJRRrrFN6nEwoFtI7cmuck3BUKKtdQg7mtkBO43liX
BgJnq12ExTkBwOJRexVDNyU9gDJo/KKikpXNSsp+Jhp+qr4BdbZyPO16BT7behzfGA3wwSJYvhL6
yFt1yHdLAUBnFc4EbAZ2pH7BI6V5f9HyiA4GooI+JLsUAdBt/8oZrdcFX3P0YYIANGG23nfZOQT8
OkgtmWmpPganeVD4Ht7TJ5i0ZfwDMFse1y0335hBBLRgA/lT1xHNcy/zF95SFWXdS7bTTiA/etH0
xV/O5YiNmnGAes+VEj7W5ewMAekHMqtgkpgtvP53nbhO/iuRaZO7adOVEorkLHHZV9yicCYEwfRC
uBfIx8zadVl7iHwUPJU67wM8Y0ityiFeb47MAToLnqmJX0wo1yG6sguk6yCBpB5M2bKNnX8ll+Ow
2ATDOqxkY4GOpJbZShJ2NYwtOmT+MYysZaSkOT1ZfPBLPeK46fIZUBjXZ8sgRubTn5QKo+UPeG7M
lfh3hbQ3FnKFn0x+S9xFANZ37K+uqunCUJp1NuAabVS31syjAG7BV9XM97MfpznLKoSZ6ualXolb
8zwwZ48N+FuAzQ2rOynImvmxutRy9hMKTxC5QNUdezLkx9oi3D67Dq6wFbvv5li0fjVInhFdYMKY
Ace163HqdEg/35bWGaGyrLw9CSH78A0WRaQ2SnecaqiBwQv3HRxu0QBDNCywkRJUM6m8V5oWOpFB
jnGtMAaEwd904nkQFCoWXhxGs69O3w1pbRwM74qOZ9AL388k5cCCoLiFiovvLgTgeiWEH6zEaavt
l77VkGH9l3YIIiCTzmwXNwWtRXRKsnwSyZ/H8YLXim8erZ45sRuL9ApTrhdQ+S/gRldRu7mt6sZx
knbKtItKDoiz8Lfy1qaB8d3Nqy1d3V3hpkQAwpsz/nsH9is/tJ5d1mrJt+ku2XBMzIXwgjMYfMA3
WB7QHCSdEUuYZfvTBuNcNgizbqp8DrqqtGKVthdNivxauhQuxe6d17JlD+PcsZIF510sZLyCD9eG
rOzVrvhqX9+a4mCsdeMQlu7mr/jNG3BCWiT4nOdx7x7NEbbqVDbDWuznXR7ef8zsAGPl8m27y28Q
Ss3kF+bjWfK+y85lMOC4sYmXoshHTG5XFoDF/1/vJerpyRQYZijflGlAM6fLd5IhtKArzPPUahfV
FpBEBqN9GdQ2Dma0gnvTHUzGYg3lYb6i8eNQKwqLl0/2BcDtUls4OAH8ivjoru4WhXUqJikD+AbU
Q9zvosrcBIy9Vv1ZWUajrgDVL/2lnTYN0vejaLTWuDPC5RQauiFqx1PVt4Dcv/pNocNgMo+j8SG4
T0GonULWeuIESrcckg+lTFTXnNuDRV82D3hvEc4MeTGIXJUBiUI9J0GMUcOjY0z2p6t9eeAE21XF
xok7SCx1md7vtXJaTn4EZJhzg4X94m6Vra0DgCOX5IRyIEwOx9GFfRUg+PjaASDoPTacpx9JloHv
h3CD8xRWYH+xofSqfCo47cowrfOhVT/my2ZkMatC7ngeF92svT3DH1X440BncqJfC8yDby0AeL0h
u2cQUrjWqW31X+IjYvk9J2Tsw9+C3YGLAyft7iWbSiRlQWmb43gMU6X0zaxDW+b+EV6HrS76Cejk
o6hbc72ovzmGg66Aj5KMkk5tMEo8IvwruGph0GLbfcsB0jEMNiubSC31We9mb4kKDd5FDRhW4rfq
ELqvpyby+eid1JyZ8826ZVQfHFN9wn9wM6uUHTuclYTdhaDle4jmmKfwHEn9Bdm7mekp8nEGrnZq
9KF3gpVhCbgq+kZDQ2zS6Sb2zjml+oNHZT+CCqYHBWiA0EHYauPqfEzZ/sCJgdBE0/Q8y5xt0tBY
7wvhhMf6Lv6YoWwmdWMQJYK4Bq2ei0MdQa252Xijya/UPd4UxQbl0bVVEu6lpz/c95fh66LhZ0sl
4Wq6+ZIWyG8zu2inPI67WPUgT+gvhuMP3X7EgzQzGPdpjZLcr7S9LcKxdBkrIeghE3izUitAn2Jm
A2SAnBcxC4f/Nv+HG0VaXlykGrIxAvm6Sb6NT8aEGFLa9kW8NK1UKSlA2LRrUfExiQzFWHXpSdTp
v5E2CeK1glJligndVklnSDeiUsmTHaeWTAIObC3J/35ZkB6kQUBPXEuNc7A6CYEqd2EVsBoXbFyV
KWLunvQeKQQQojZF0TmRh6JJ3aR+2ccwsnZaan+M9fxvvhHYOyeD2M6sHFb4Qy5lzf/ACenh7MQ9
3SOPU3SAFFWvI+mBDxb2qugNo8PKA3grqXREJg/YyQ/c9dAlEUl1/hSaibTnvVzIiw2XtibDfLDz
FgRSDKJtaCp8ifHUgiKPJOgLVbLQFzX68onoH7YkJNTgzZKKnGTH4gO/frKJ8M5AcYfxNNRHdrEO
5YaC4v5L2rJofMXWRQH59YfpVfDO56VuqxeNc8GfK2AUSl6IjPz3u8WprDus5cUeVDIvSvGH4AJs
RZBd915usV7rsnTyHS6HYUdirWhRFTWOZRPW1QBY7R6vnPllwuFaPH8QkxYhqpo9c0E/b8UBzWrV
qZLwzzQpcAi8PbTI8t8HXLfiRpew9fw3hQ7L2DG3/iFDFMLGv+XAxi0OIVfpvMXX32iCd9HRcLlS
sZYd8ip5A8FYMqDeAMbLqzBto4/FN52r5LD83NABqo/T7VlaCYAF+gMx9XT0hwRr/BrsJfvcR0QN
LlEn00mr/r9msHxJj/PI5zsJN8dkfnVd6Hw4uGcRCNema8I8B/ll4EYrYZPuMPsF09vfqRsSgWRo
DRGf5oCiJ+cieQ0BFivHex7AWrHKnHvzDyFk50N+pG0DjcK5PWX9ll+DmGesWpTIMpVJ3jiWOho2
7KOnSeK++4Ejj4PA/5gliSswTnJDWgSD2kJ046byUudLXbQ+RqMenqkeIWTSveiNgyRnGADY4s8J
ImH24OifiAZ3VBhJkxBg3LQolkLH1sJpFLQ/vtro2HZMLhls8U28Gt4Wxms7nsqOtxtb8JmC0OSx
GxHTU5eXuMV/grpcZo4g3jCO6KD0Q1WRBEJricLWXFyVVpfPq9thjylf8jC/NxBjJfKJK9ndfzxU
wCQPzPct14q2LBkF9RLnXTZr/RdaFnoh/EOl3edJi37AeJw14EAvHMg8GuNb77NqfpTN8jm5jtyq
/sHkrtu5CbVd3cn4+yqTGnKmS5iOhxBq6OEFe+mFhI4awBQMfr3pmZ6Q2A8hxzms1+xoBqZ9AjIK
+Luw6nHMAUAV8Kzx+N84TPf2TOthLEGwTKdOALd5ng+IhSeWgSGmbqfY1y/MldynpZO4REGqZVfc
cfdm+qR/rErJQGoWTqmk0I7mWGR4xhsIu19kJVhPfJfN9qXFlsAW5exOShDs8FQvx1N6znhYRqiu
HTclgL4XOEWyyosMKiBitTMy+halnES4BXYqZ1k966sN48iGPSsS8VKmMNqob9+Ld0tLHfihjhOU
BlZEXtnhooREYjvWvQ43KIbdMjHEnI2z8Xs2a9xGHHZUVmycY95uzWTna55K3Au34bovU1Ep73YM
1zEef3NWWMB+Pg34QJWkaQ7bSuwsXK3pkuQN+/bCiNaeClywelg4BBjopxz3Hm6AaNAeEo54+iXn
OcvGyc/1MhV6FyvPG7ioeM0zBq679gBE3JnkspUruomyZl6pdXAdLM4F+OgPXTujbFTW6KxcnxIw
JIz32CGo7tSPSOM3uIJytyasgQCclhkIxMNE58rD8j4Sg55E77+opTTPysdfhaJJDcvc2Pi0KbpY
uPalNbvUoOZ1AV75p7Sj55uobbOF4cjCKYgoLhzTqyNbYp4NWzSzBAT8KfnpoYDF3QkNwgHiSbbS
pWF6Cn2Y/2UKyYMeXtWVADqTXvJZYwC208iJeV5x/YUJlhHSXI1NIm/YzJQOSk0gcz8+87K9TA+6
1xpAV+LyI0+S78ZGPOXtFpLskAc5QUmzTqTHD6Tx+i26LBDwF8M88OuN3ElEV5L7mIPpopxEowUJ
dLzhp8+hZrrrtrTNq9t4UL2WlnBCJDANcHIeh3ShR5xNMabqMAegkLP4zB4Z4/2UetkKpVFzZIUk
WUSypm3nQ6sJZfmdgSIavZRLvWdHsGzkyg2XyV9/U0uc1vBIu7eSFQU5sOqr0ElhAwml33pstlxz
uI3QQHtKJcGowAZEDKEM8lJ8eydX/fwsoumZw3GjjpYxH8ltK7c9sTYR8LO6IrOg1KqDIpLPik5z
LofC6pyzA/8n1yg+Ws50KOeNiY5oQX/bmWv+OVsnxH5sN7lF8dE4TCY2ceLpm8mFwJkerg52+yG+
t9SYa0AwGKe/6K5teugZMjxM/io7lqLAiHSfYAwZKX0oNZoiB8dvquuhSp5BMrVfAfci4ZfZ5IZv
csszQ4C/th+h8X47XT3x3ghgWbYyff8LOt1z8iElXh0NT4S6DDFxg4CMzYXCXeIhTWwF6oe+DjHM
mvkFquEn5rUFQf17lStiv65PSvZe/EngmuUYqtOuiZT7yfDTbBZj2yOqCbRBHWIepn21Kajh2LIJ
JKjCENscqJvDKiMk+R5V+MB1LE6FRksCF1DTGZ6C4/YzagmeOmfUE0WsYNGHQnswZt9laIP7fAjZ
8b3W/kuOpYLx1nwbnxuttWN5hc8GZieVZoBvMiV7e6hu3IuT3cqwzTbXHbK7iDHsFNZBhxic+ds4
JWfWHo/To+jJjkm4RlkM+ikM80U26c5jIFEP9AjPG94MgqFp3LXyqoeqf566SZoR5bbrzAOjcRAK
dTPpJFdCmxP2PLQ1yKenvH0IMn3lJ9527xHUwpI8TksoY8ys7SipQxBXbhYJQyddqfvgx9mqXbEs
mo3jO26TxilMpPe0Xg3srR9JewGuI12G8LdoNiZayREdQD5Fqqo2JuVDIU8pzYrj7a/xD1PqB/pA
5T6XONAojP6Okyuan4Tu8Ot6/nLdGfUQfCw4Oqzv2wVMgxYEi+dmzATVCXInbLO8hc6ZNT708+zN
FTh0lBUrE8xnNePvpwGhtbAbkRD3xzy3GdUoVb4cM/QqipWyE2IydW7ZLSIMrmGNw/v8vnI4tag7
zQk4+On4C8P18uMIm68fHK6Mf+BEE0V5kRg9KTKvbkbC3BhpeagRORJaG7tgF4olGImcgYIO4Dis
hSeyU/knss1LrXMlr4A9Nc4Wc+EbgcCntdN2eRYp3+brEA4qq9+h5Y+wbq7VugDjkKNhpGuV8bAl
xJ5Qdk5CpvthRAAINgIeYeH+qcJkzbuce4EEk0KORmyceGvwvI51uzg/i6uDMM0Dw1avICzXjmK3
WuOeb2iF+Y+w+NgSRe+5WPTVHJUj2ILyOha4KfpXQFXRCoJ6rPGkgbSvpJ8+JD+/4EzplITa1wCe
C1OtMqz7tHgpkRsUihrWQMpM77vWWzenRr7tkHOPrhW0KGCqTSIRdE0Sr3DH9MRjgEs1Aptj3Q0X
GnPDKqlBb+KZFExI86ey0GdUtSrPk22JU2n7/LB5MV/mSQId1YL2UB3plvucwMLK0YIA5xvdzi4D
lvjO/vyIc5fCgr6geCbPsnTDylCilkXbAzIV5O8JLbzf+rW3IM9jnFje1PKvS0URYF8FX6rDClHw
Yp2MQfA8MTcpQfRMl80MifLXdu+0Oz9dXw9eGT8i8/9u13fydpu0vzc1PuCQFp/s4GrRJe/wdiOb
xGsDcO4KiS43eLCpbngca120pEAJ8vFsl0ij6U801F2rrhHY5u602V6Tv/KH3N10jw+iC+9Di/8F
3AzfQrWJoszaUEsClRWRswKdcptnjiPnAdcjcKAqLTTIBp6BEMReTeMzANaAy885l35IdgaZ3pQn
kLvYu4mnmroIe1NRNF8JP1rvuWmFuG8Gh23KhJBFjtLdK6NTjEpltblonn687Cgc4CTRee1897vy
B8l0ChcNiaDZ1Tx0c9rXtZLuUxVK9QnZvUElicmUBrUBZmnycTZ16DLGTsMMpDjR+/NgD0apuvsO
ipMd1WeEEo8TG+z3Zfx1IbWeVVddnk5IURqvuIQ/6jxnqD63xtnjPu8GyuIjCf6qxdGa8r002Cuz
SlyonWbaIL56iC4f2ezeEVnDTXz6NQ8ze9oArrRWwIeOfCiHXphAyDsqwpPpJt1kmdXeDx6EGCqN
Dkd88Z6nRL4UeERHfu/e1yanA5faSBbRn8ucH744I4T0CdRZIPY62mDY+2knfpZqfvEMdk5LDIlj
Fv6u6raV1rR+8sG0FZXB0ZQCbv7PycUguYysqvLCXvuXqvZnjOxwlP0XELy+73i/9yh3GPvLaquU
9kIJoTeQpmQh/ygYH+larzfwIdzQRY5538qZIuPiQJFkM+4t2b7MJ0o84W32XD+2a+jdrV4ABXIU
6Z+rB7yXG6lsSP678p9Nb86tolnB0N9yaMGs9MQvgHSFiLJw6yl/HpO/UJ/O9IpInQvfA2haHj+H
olnA9EtoJ0XGUss2iylSVibTrJ3/5WIJQkhUzNHNPXeS7S0xTIwtjmhl6TibBa1c3w4Shzl7Edx7
U2zaEEoShcuZ0Nb+hd2Pvr1W6ixzSM2Idu9Wc/ZLS3V76TcnqZWg3kxczzFws3r6MvCoiKWO0lJM
zyQfCiLzqQ9GJMfowg/F1Nv0iP+RvFDqCoC7jpqyenn2kbmnP1oJ9UgtPG0R+rL91D+InXDWkCjV
v0sXf1u/5uZfzIdXDnLo+q6QrCks3Mcd/NUr0NPYff9wdVDTjCqMUZVRA2D3p5Ipq6D/tYU9OFEE
qadz1XC3nAL6Qy73j203UVBmW5R6V2fDGA/c84PQVERyaegr4UjgTGZLgjAwKR8R9XfpQnGgs9HD
0vWBHAxgQg9K5qoyB3BGiXBsEeg6DdwEriFLoSaUuKolDWhN2xMtQETOABe/XtvRuVwcraJAlobU
8f2Tp5qdpqT5xViKMG+lRjmIMd9KFKdfSogDM5uhu5FLf6uvRUrRKU9wO1AEjEnjYjjW0K7+kOUz
Vo9PfR2mViLeizXowhDMOcU3LqDnxFlQsTx148c38y0ob1/h3rW9F1kw4R6qa8CK31YRyHWPxCdu
dR+7FwVzOXGi1HZrWV6CGJUMYkCxlk8gGnZDOnRfJlhkEZ+AzJ83o60fYsbiEhAcn1cfciOtnhF1
ETTSku5w4GwvgswNnBBfKQP5LlF5cm8Un/188qaagvz+UL5JHPUI9bjhc0G6NoYn3L6hQ1zYomME
EttAliXXNaerXfGeH0k52fdgurfnAT9TsNZRmzniPm43L6cN//clWmZMJtc+qKWpCX4iuWMjkU3T
Ea8c1PHG8fE+CTTiRI5+l00zlLnIm8CgYgA5P4Fy28ubf2tafa6qg0fSLKiVjoSWQwlxIMkPfO1u
RcudBGPKct4RP3RyBeDnnGHR2TT9oIgqfTEV47oCqS1/tzH/VULg4ZWUct3soMw1VK8ENnm6gRJ1
kJd0+ZF3WrT+NzjHVssZxufa03LWnYrBS4e0lQJEe4qP5VVAiXhbbAfz4e/04M3UkTMuCFG0UVh+
AD7U1bn7gIFsPhLm1gB6AdAB/NgClQQs8Cf3mMfn65UIvh6/V2fiJGX9Fu1SakaKIMsVZNTSjNYo
BgXlwN2MEyVxDZ/EdiRTpFSpS90J+8y81AHJXfAtXnZm7r7WQkuDM+sGgeI1AwbLRnxHDusntsAO
W95DKtyzzcp4QrPAINWlHD44AXku7y87OiIwK5rswkjeo2JCx/Bu/kS2BBsiyfDzsVlazY/zWI6o
/ayUFC9+RK1H8Ja+q6wBaDfsOLplBEevwowAVgVm5i5tMqib4IefF2TgIvMwwh/Syilux8Q+4Bbd
IBWlDMiFOUZ9GSVNd+qfYzWeqlRRDda4KfGR+y0i4ZbXvd96QkBuOUMwEW3Qqiim7yZmMk6RO9aI
PXxfAh2O1BfOGMhZJ0E2X4jvF97vNz8s5wGJCZHPtEQ87ZiVYOXQJfi7GyrgoqN1bMgw3DvpfWtT
7cFfKhu6ng1UMcx7rU0WWBUEnenGDbNYX3IcwEnDCXSXzrGERw7w+7PWyIcqTdXT7u4PZaF3KuqJ
gFSm+qbzI5sbNZYSFsHuWbmKRmew7vuN8mFFVmnHRfKS4hNfU9jv9MyIXmp3X55UJNUtlrCJV/MX
1tFZ8NiDKNKqYzu0/OQJeeFc+Y1LpG+FLOSc2sIOAKpHcGim0b2jHP4u2xINTQ/Rxy8XKVyn/skU
n0ePah4sQM03tQxlBt9nENIXLa4guV0ICxmzYQQLRSkncHN2l18P8tvNQu19dunknmVfY8jbG2xT
OsYV3rg7NGikE0ZGv6CeyRDxOHMa34Fgv96GZzvgtPcg7Q4IjECxuoAaU1FHRiowrk5OMAZ1M/wm
RxFuwEpAm9NDai8XjMqk6TTcHuFEL9WDrcoRjtSpJr0BkledHBDXsumillA4wRy0XJDvClyGOnzh
qfZ8TvLlMUuCS9Or62cCyWsZVkRxAh0nyppsJwIS8PWMYfYaPx9PzMBMi1vm/cQw17mWXk5O2HWj
zJpE7hQi4V2f6DLHhaz+n7a+8hIOxSChJpbg93YXxTisbrlc8OEO8fWZWzj+bwaAaYOP1eINZz7/
A3b5PbACbJk3gsghd7OKd4OnlsoEcRfJE47cUpDeWmXehp2JE9lYpti3FDFSqT1D75NllAdMFwR8
+peDxJlak2Wf8YGPdtPaqMO8FOREdlLpkvnXgJ49OFM29K/FQ+QqPqLImxmrEHYxTd+tHHiMK22s
lJ2L5ESaI7Fx4/YVUiaTn4rxQuRwpgYXX037GwEDeIDlFtNauFlymmoXvk0WnEkQcCZkXSwXyTQe
v3Uopl5bMtXcxgIcmyBbmQggI7/a2AV0MW6RjbXAuWD7eAl/s6G+bb76jDxYbY6wZWYvaLN9s/xG
plh+dGG7YaEvgnK+rd3tZx4u241ezEwcZK1nfrrJ9KkfJgO0tEv/k9jIVFzIhWWg265e0/4Rs4u3
ZP7ZaSSOThJ33BIsRy0FGuGM8V0V53IdRyEjlCMIFGTeE9U59TuPTdCaCm0l/TUt7+7yrL9hocO3
RWBx/7uMORwwU4kqIZE8ql3d/i9sFBFnJFlEvKtNU/7lFjFCqXR0wH86A9bHMQNXn8ud2mB4w/un
V/YHRs8bpgzyuAyujfiz4jSbx1QEyHSiRUSoqZh3+91T5F2LR7kWZGEry7Kooqw/elYCPbrVNMZu
ahVDDQrNhHAIC2p4gSb4tuEYii3+Ev/wfOlivIq7Ms9IQS6PUtFL6+yqbDqKk9Lz9HtJJHxz1SVo
mlALQBHzhFBS3sfHniK4Azqx+DzUFB50Zy6JOqPhe+ylfhBFXqgO/FFjN7ktDlfpCr001niJeiMw
HjyQk/FGS8QalB6EHZrrTv+IGt4qe62Ya8vG8erF3Au/bzwk5erkHGlIdLD6VVd66lhaZS6Gr147
yPtUdOuwRApledeV5HS5WWaH0JS6qOmyXyA9l7VfP7JYccXZm26boyCMy1Ri/VGHkkdjaGZpB44e
bnA13d4tTptSrxHNhuIB//6gwkFFjsx2EpZVe0DDFKtpnGVw6MFYlCObYSkzPGQVpAvPoc3QdiGz
LelSGM2y0JwVc3yVFGakVTJ3yoZrTZZc3om4kfdyD9fZN6fPsweAfcuq3Il92/a/QveT2ULQIzIu
Y+bIJzTsyUSkA0xWpG03xkBvMajBuW/7lJZgO+DTszwgW7o+n4wmLMBL6nBkgnbskQQKaf05b6T0
2Z5jnqGGI7aQ2J2cTHv4guz2LasR8hGL2GoYvHVkZa+0yFxxhFMx4pFlOMDrclIAWFvbzS3COoD+
DYCZzo+KFUKafcMPs+lYg20OL2rr9T0P6xQ8lrWXM3W1e/Aud/o4j144IhAML4gRUIqAWdR4PCIk
YuSP8bHD0GtypHm/F0bKVIPlQqMQNLGWZ0XMfJd179K/EB9CjdQajdjVkl8d22YvLghVVFfCXkb7
nz7QFAFo9MuVC6g/gmsbWsUdXgo8AIocARKTZjGSWzUNijMnsA/XqKQlrfWghWGyQAogHpMY6hpB
daNJFJFZB8ffHchBgQLTHW3PdQoUdAYy1p4B9L2Ic2tx+VHt+kHmJxDw4kpAjS07XDy0LCVqsAL6
VnBF6xXMZn+aKIAzQNfzb81uNaShGF+R7GMaRPR0sgcVmO1QtFUMCWRxBktp1JpHmfFXliTu4Pc9
l5eKTNwv/fmzOGM6h/SP8fCrP70sRaj3WanK0M3uno4r92au3R9U1V3ryVlsy0BCQdmijdLRY5m0
kcsA+5tUll7XUiaPNmBFdGfQq0oHKHwWisxwh+umutwh8NrK35bnnOTMVsKK9L+IZWLofZNNFNi9
DFUVnpCiSfNsdS/k0U0mwhtjHmAlfAVwDUmYIp1+MhwARtDl9J5I4fgKJviyfkYNK2YIl5Se+UZC
JDBccgHFFQ8hZNO+Xn0wxAz2f30hXV+iTGbgo3O1EjYmTTu6wXN2cIi+VvhF2ywbPe+UmC6ptPgS
2w2cHUoMCQjsUwWcaAIPEau6pvaSbEJN9fGc/PV116kpvHggcXN74XXZltA04MSozhbib762rtjq
3Lzu+d5hv1cFbeFeBLekOCkaadJ9XkJt0xcLc4SJwh4vjPHHpi3ZICyqpbkweYvmsQhNRuezg3U+
AAB8rco1+MCy9IJkonMOE5LWG40VZMMIutU71IybKxcYPtfl5zaRDw8cDVLaOKvozsoP3O+Ekl54
SkKuyT/bRAR7atEC1fqZNXgY9U0kbuWn2t5zgg8jfK/IVPCyoqxE4cZXQyAfDGcKi545sTb4ERp9
PfiYzL1IVZxreoi/Javn/yF/6wwdH/6yu0Bpf1xNV8sLokeD9BkeM257ZexdQkc3+05LWRtqg0dA
mEGFFXSxg49Yvc0szfYa84x42qGnSyZyWH/ce1Uc3zxbCp7M7HuYy9IpluHAPMO7uuieCx1Eg6Pf
f16FzqCotnzZB71titP0lpH0GG4DKhYT40tK03370gEBBv6fEjuHl+ptjzh5pWWttWAjZHe9SC1l
P5MB0V0yJbd0jkr5To52tXswb2VfNzi8O+nyn7P+5ymDx+PnFoebA0tPBg5X7kTf6Ye9un/ExdH3
2r485V2rIppEXPIA9hGlelv3+pSDivnYpeSz/vHezu9Ajlez/VgtAzNbp5qbBhNbAHrfiBaUzFiv
XPVLBkA0WSTk/DlbO5mthM8S8FhV/Zr9ZHxCY5ilRMV/+1d9hPtCf1zQyEbYyfY//EFF2xw/JF0b
g1VaolMwbg8+qx0yvB4Wqg2maf3gtbEcWAJ6TDT7DLhbkJwIJPPGv9UY9tto8l85apuu0+P5wOxn
a5JwrKn7E5GHSqjqOAxQuJOTYELNz1G36AC3gxfgwl8ZaAfcW++3ISHpLAHmBtLg+iB2LShdQ3bJ
kfkb0tck7b7laXlp2T6i2NxKM2Brzm46KGowuYA3Es58vL8dxAV+/LhL4z4pkmQO22stl34/cSKH
C18W5vc0JP9SaJdfhnDtCrUMYCS16XK0RVlKf7bIdpHdODocqu9blGStgsetmUg0MgHTeHCfMV8N
3ms/fvChy3sChG89t3pJlNB0N0AIuWUT6QKcKelKRbw/xxOC72YAf7yxXvyHqiUpbp+MK36FrV+/
I82fub9wi04d4TQZ116h+rZgMH+w/hCJu238pHVwQL/meWeYpEZCc7p53xrJ0p/mYP/TkMYb4p7Z
7spGx2W9Zoe04BUuYD+bKHzzL2oC4q0CadCzk2y0adpWqEzc1rfYmitGszoNYYQNkjZT8zE58c9C
Q3GfH8LXwjbipCttVxLUF/SoLERlAOBzHkjffB2oTM3tm3ufGoChQTzYra73nRiqE3GJEp8jPZYo
WkHgikqYQYoa71yOBcnBPb1hXQV1aubMmu7FRlWdL5LiGryiLEYMZ0WDkU8Xl7vclyWp402SEi9V
PuaTQnRX7PLShQI+Q5Qm3guqKyHt0oQzZEVVk+0Ti6fBzSP/D9V7AJUv+bBo/xTQrjZvgQODTqF7
9zrNDBImBzm2dU+VqdFeR/FJUglApLZmjGTWsH/FloSmpXiLLzLrtB1KuUCiPNgA/C9Xl5lQLwpA
CJJP6/KAgTNtnUrX0aHjt0IX7Ebm4jA9mJiGi7TS3uillit1l6gAVPqiVBmUMlcO9/nprzu0GcCw
QkacNS5J+5+Q1va9bNI6Ovs35jvam7pTzSJ5dAL/tDQD+HmVf4OZu8ypDOBL7Pl4bJe35thGJesU
gY8Pg+sFhEHrEesEgtAhKRZfZPZwJRHegMt5BGWMgkj6usMzUCphBF4VfRTjSwNXP+WKVOOpOUqn
bMlCY48O338Q6j4SteIynRPTyGJeX9OZH16e+oKbOZcC5myddTWunwbeMYTpuX0rGcEvQmdTZT0k
GaRN08v6wgavljCGGTc/rbgb8b76/fc+BtULvwlMY69rDvsargs+6PUO+n7Po9BHxQxUzeVEBatm
fbrVB8mE+kdtBXBKzVxMNyOW0xie9tw7Vbh8k2Rtk1SR/OTUqMvpw7ph00Pd/QedfBiPUuPiyyJp
30/sYQRVXnt6Bwdcj6xDhGsY+9D/6O0Z/+0aWJZDyR8bu+IXiHoVPfrT6QEXFnJvrXMzhl4txZ2Q
HnvPeMG0olA6oa7GtWmKfGvO/x9PbLtZLLO6YoCz//L40B5H0VpLE7NvUdSb0SUnkFVFSq2Q6A2Y
rTmKSTLJL1Yvb8rgkV9R+6s2DTVHz4UoBfOhSIPQNmTVqz3TOLSWosvTSf90XjtZCZSg2tybbbN8
dIn+PqeZe6U8xzN6oK1Y5ySqp1Q+NIw9D1K3OPgro1r2cnntD4+1c/dGvo9ehlxEX46s2mDgIyjV
i1PmdCmfiKSpnYqu0UTap7Ag3nEvlHMgFr+Hr5/+ZUSdk6M+kOsYDG54/YSCtI14UDBjb8uM8RgA
vutUJiQe5mlWnsWtp8geIr9aMwbkluYafzFVYDWj+PcoVv75rXTHnGk7liwQHVBTq2+AcbfE+7Ox
kY38UxPqi1/43z/P3JNS0TduWsnJlFR7wZ7ALKktRzD7QIPGQ7IAMDflAdQEBrucYg92LNvX/kcT
8EkFlZ/M6bS/JlleI/qElqiMQiLeberA3GoDJZ7wBm2xR6Yl8GG9rp3Lx/wOvisbpPgqcxldMW5t
iivFCCfsxIsQhZLNgWBNLKWU6EYvwWpxWVvZtLlw7l5n7Xmdc38N5mx+8NOrXxfY3029W01PUM5F
5RBNCGZkW3Rm1vuy+s51X110qFdH3cnIIE8RnDJN+0hPxR58dBGHf4/7NIh1vkirnoV+N85cpop6
IIR5hvKvy3fFSpXFD+1McPjt92V6WkVZbne0iNLgE7lhjGc0LfOJ/ddMCZd2pqFUTRWQohYvnQ3n
y11OMJv8VL0hmrtLp/8Q4A0jYcOsnD2T4RJUoFWwAn8f/yHQWAdq4m2o016jo+Exul1l4pz2ANcW
UzVsWmeryoaAp+ctOQrLw/KYpZq/kLR4ycRKm6DuELJLUGod0K6mn1T1bvXq1AN1me9F7UEGDBCq
7wDjaGyobmE8H2J7RnWkR6bbAgJ2jffmp11x82RKy4maPuvGT5/dPP5XRXZg/RbNdHRIZZPuQjhv
lV5bYLA3MEaLsKqgxK/fAAyxtBoSDZZkXaqhzar+oaTFjiLtm+zkhXBvErH0KASZ97oonxbSocfw
5cgqdfEn+aEpnKsjY3VVglP+NKkkY0gD9b2t9xq2a8IImI4oG9G84D3e8Y44A5HbacwYzfdqjTPb
S1cB5VfM7lZejrMWSxN5B2beszOLIIxBhGMoeE1YPur2aVvR2U0KKT6yXMxWGXBJA+hMEG3T+V7R
kJ9qcX6HvOdDJ0DOLwbzqEJU1jh9aP5rwwcp8317wt/Dh1oFSMuyfdU+8TvJXuo6P/okA5mRxHes
UAE27VGkJMWYgfZNRAPZ0Fz/LPCgBWUQSHgCSo/h3HxFr526pMCP1MrwiY8OSVku5iEi/Q2QRXaZ
xWIq2CBuERnIh5KFC6/rcYG/Sb0eEgAAkK82A7nWTgH7uPaTdqDXiYc4yIlvIgtH7BoLdoNvw+47
lHgvBYxyRIbktAG01zjgWo6ergWygAxb5GWXkUNXNyWf7U3LFA5kXbqhUia4l2q+v0dndnDTFqEU
Tij1YAZgq2ldhAA1bC9w4us962HgvPpJK+pmT195JQHJdIF6XXeG/IRZ8Nz/2zGhV1Jx0xzHQEAE
qsBMOD5OoAdYyv9P+PNn4bXfZQFUkxwhveBnRNUF7CTXlj0jXQLk3Ne4irKPJcKL3XYmk/CGgBfA
YafiZKXuWeTku+CQ5NMO2bxYBPpma6Q/DZty/LpWXAzkuBdV5DZLL+7dFEUEab6g2X7+F76HgGeD
zD8pLQkKULOYTxlw5pOn4NGydIMsur0ElMwPfXF7bOOsKqR2KOq8NQJtJcHTXnQOZnfzPfIQ1+vh
UOZhAt+G+MWQKXODdl4KEKAutUf4vJUS0bj9ZWdjQ3JfFRX9VLYzlTzbaK86v9IBQlrMlZJb4nt/
89d6/3FikmCq5cfqj2WjeAOzIVAU7MT957SX7Bs7Vbrwzhlh6989dLrg++ydM4wgmCbqFWyHUEhG
lshIZLI34YWmp+pEMWtAssgvzLEfvuRg31fOSPZoKbmc5R1DgewFRcaVVnrUOhkxqafefjcmrtGe
tx1/5uNm7ycJEp9tb1zXEvJBbavrVxL8EHv+/kpBv3JsnPEoGIH8eDukv4imObHiNjrKTC6R54Dz
ZF4pMwq04/vS29q6nEFq2u/BBMVCvYHlvEZG8wVVUUQTkBMiPsL9lroh9yaH8sIt4g+hqq/6FeAD
3MUEeDiPSXrf1Fa7FC060eQNO4RFAxRTiaSAESLaMr3ZUGXfOKL2CYPgvs4qdLE56bS0IoRjB3iD
Pnv3lZ2wcAzcaSc3WtHgPwdkvad0onF259VbyUuyR8+xaIz8wsx1RaSvvqdNqxlIFhO124mcQ6Lq
UlcxOfm4Qaec/x2IWMp32UgCJLhgyjCBsRflvwXzWShFyLeWAy8z/Nw+mpR87l/+p25T4U5bbOlw
O30bp++UhyUiYfvqgy4h864iFksj5GqNJFVfC2kpR9pyAxIKA5yPL68lzIIKSmTThTf4zTeYdCVy
aNS23BKqScnnrHwi+206PTiqS/1zyQgbGv69NBLXAbOyVuPhTpdfDDOQbv9NKm3FJTbwAfxY5fIq
vHGdXJk+n3z+EabjfW1Pt4TK1TrFdqzo/nJzCHgt/nbSSuqRLSga7SZwZe3/UxgK8v4t4gY8odxf
6S32SvYNem04Lo0KGvi1Bp/vOKGAtmapqN+8JAlWvgSQeB2xbSIL4b21Hk1wxezLL/xTZgOof+Ck
7pI/UACAtJUpS4JXzfXnax+QZnTlgOcV5c1gdliAZbsdvbSilFMWEZrxvmVPixyFLHH+NZYqz/6x
qvoeDUbPzelhRSvmtru788I3Uwd2XhjVE0HiPmbPf1CgFisY9MyFHnlz3lkUKdgglahWJJHr0qa2
aNOlDn7ThvHru5fDLTHzjuUUNijZGJXbz9liZJWSuvy/td8qDX8tnwQNMtyhEY3JlrvK53/5IQ9s
AjXNeE7yUI6ucA+2ZIDSILvvQt7SoC5aiAesnhY9LZ/qZ2ejjzg5hrKjKUsktTTdwdsm+e4bUzaJ
t+f1Sqomi+Jy1AUSR5cJ25WfjprPgthoeS5JhvBHD9LtmHQGEdOorau8ApwwoWbKygA9frHcnnjk
BXQcmSKchA/P3sFKLrbiLXLWAFWEWpvqJot8oVP/MWi5glBRKskcTZ4uQtN6UqqI+h5/ttezoAQ7
lpSgentvufNkUBhSyUhQbmcHEApCxDaaTw0DP8mdSEoshbJV0P73qkUI80+8Qno7Ik7MAkvYlwmZ
J1+9ToyyClKdu1WHrT6pNaTXH0jufyQWQWl9Ff3J6mh6o33+BK+Up02jocnMiJIfSZCLcfjREDJ1
nWPBN/CREvEVV7DabF74ddMHX488Zp00Pe4VXTqppMgACp1Q3SUmXscexIgpHJ/cQy60RbOEDN6w
FxeSpUeCizbXsCDL1AvmOZBK3+IVeWNQvZcFeLmRhBF3mWBXeTTKaHYCes6J8Bmh4hPPEM2E9NXf
JpJpWxntd9C47IuDijD6TADUFPKuUUHmLmnNRHIGZWwb4DkOy7Ef8aomWjuDvdeAqTpG1rA4E202
0yOgJdPhL8TK+hbBmXGsK3OqhgMRzHfKCbm7ivGAFgbCBNPIVrP1Y0jnVkZKcx9vpsBLMmMugiqe
TcieMZRsgUIvI/+B8K9viSqW6JnVMHRoY1lNZ4y4KkfGIAVpW6CyGHNHwkwD9v9QLPxoyZiXo+RE
vzdzMf54ICK3/NvRWMLTQFVFFm72TN5pjsHfYZba3yRKUtbkzHPewPJ9G1UWoqBRR1OaIPNCji5p
30qra5ACOnChveU0gergmuxOQMcNhtlL1JSAQ000MAoK48PcagrhJ/aPmdZuvynAtLZnl7cqJtj2
RNhtnrLspo4LBiPcGM68+qVzfWocYVbGgPupBYbkgjphiVtX+5ZUFUIG+iEh44YaU5LEAqG4Rseo
fmwNPLzNWkajg+YP7wBEh2YCZ51fS/KVB0MHBcuHPECQ4qtmPHX77d2i5TqGys/og3WDkR0giq3W
AaGevk6OdImKkg5RncpjYuAcQpdozPsDuibK9NexGd2AqhVv3FTbLUp5EZSgasmAoM+08vonqYyx
J4sJnAWmTojPsaUqQIylVvo8Y3Le21hSv07Gwa+/LvvN2mOZ7D00DD4VnfOFHh8mkuYx+PChAx5S
4ymh//HtUbep3q2zTzIO+hrfTBgulfcbr8r5qczzdD/0ZCnlxBmpvkdCo4lxdU84NZu07z0/MODJ
PsVL59V2KxfJMzt8Gwcqssl2pHFxuEVyYowdRBY8OiI/9GZL25MBXVkLwb+sIkwaS87RSn0Leo5f
FDwYJjzx2XDkDDXk7BPDonqb558BKyqrdCmpQ385rstclElhHGPQahNsUK51PJkEvx6i+3ertTpb
Ke5Pt5yt+2YmvdZTN3KJVCLfjjKhQcVSj7SeX/Gymi+brNBCDbKkUrTQO0MBV84m4Tx2hDchUJOF
oBeWsqi2URWLoSxOQl5UOCsgdKRBWBrahxsT57Af+7BTLVO3lSpj7Iz5vAukRagp3KCUQ2TPGb5l
L8PDLX9+gULME+qgtcCjjLRtU9QapFb8frJHFNsg7sfJjd6gPOq21qGzweBrd4pwt7qhN+092R9f
yHHeqbGSG5CiYHJxhgMWp652kGpf51NNx+3TXCqnrPF8RbEA5zJBeEez/OqGr3wkw16XzqF2Wpgt
x9wOkmwl8nUJxKRDxw7O35UOTU4Wx1bxon4DAps1Me3KpyJpaOAAPZZv8uTnP6t5pfHK+YyMvYeT
4N7/iOzrUBzul/bryCQgmABEWGnMLJuT60kD8e0kcXc1V0tv+U2cCMcSGyleSTS4LSwndB24gV4Q
tXTJKcKAq5iAHPXv9L3KZICVdNjrkYNtZoE1g9571t/F+MnlirAMGatZVSedUkK450Go7QqjdPu6
dvM+IGnRrf4amcnSoPevWWmlEq4bBm4IjY83wR08Tl4m2G/nRW61Wo4gz/8agMkiuI+IyNLxOQ/G
LArVapxcFltxaHw3Lz4a4meZYhgi2FLPCVHqg6s2LhHgkNethsZ8yqt2pX78uPVUzjRBft1Yqvcz
Kzw1IHaRaPUlUx9d1/i2eKDrqgrwwKr0aTh8gyULiTJAnbT4aph0nR3zhL8B6PMSYz8QKkz/cOcf
NclDaAO5D7XTfDHn81FHoaavKSWEQAS54StWUb/DtkR2RBZFhD8eNiUzM3ap2YyEcALXJ7LD300z
jGnNSxSSKn+jP+6CQioCdd95/W9YcRvnW1UKaTMXBhfGaG+5JAsUTngFMRTjzu/d3ouyJ6dSNDp6
Qt+/Ewa/tibBSXGbjDlcm/IQrDSyuiRIZ+eewBSKbwBo3YnrdPPhqVwJy+JDvmQGyTz+qGgaYxSK
Ki6UY7LPu4Im0cepEOxNIszP0OCE98d6WYl62IifDIrKvwpcsZmlRiO4vn/0qZ47yaL3D+ckemuk
pwSIISZPNn2c1q7AfWpQ8IPiR9xUB5HAmMtjKuuIGIukHw6uQG1JJ+7b5Y7ItqlL0uZJ/PfVCi5Q
2ira4NJPTgLld4DXpoMoRB/peTCM6VxQwCzmSirdUlGclBWXueLZ6w8W6i77P7NL0bmLnYeXhteZ
ho7Uk9OeNS9k0/fibc7yO3dtT7ZHcKTwqwzbhR4WIOAK98c/aXOwqDM5u7v1l4nkEDwuegsJjhlZ
oF+LVv9v1VCZKeLssf/XYR4Y+wTN9y+8kDf69UL4xrwe4dwM665uYM9QszIme++LKpIrlP1bVug6
qeoyiOA4El6w7Giq8Al8dtQ1K9Ghy41Dy738QZAbyYzv9R2BAiQmoQfYfLowlbecr7av+WkWMRcB
g/c/lHkgsXRdZeDplBjJb3DxmyTVAC5L9npWSR3QJt5DzPtlXBPGmqjlRsr3AvoRBAI3Z10W93RA
o6gdi2Py8/1uPSdVASqQVFY/iR4ioxWR48ajEmPA9wnvIe7NVBcgOGifV9QA2p5yUOPXcNMbhkEO
0ToOmKLMyXwbVa/Cc1kgV8DOGmgKxGNpJhxLTEjon8c549y5ZKwl5zya5tM8Uj3SzWQ95N+n+42A
KdhL97RIbF7i5BFgpyLSHJM1Ml5bFMz53pI6fpU30x4kjDlXQJkJpyhVZypHgYaGOJpOl+YFk5f2
Q6Ny0xjs9/DyfBlqONbaxDyGDB29QIV2zWZjcSXvIZ/71CGcGXJgFOdiMN+7R62OWcpVuR2CmsUH
EUtuoNJYS0Cpd1IMvNyPL4Wt+II7dLGeZMY1l7cxvCOjG+N7ndmws793aXDbQLy/xr8MOq0WKEiE
Wtxq2/QBGPEBeo8CTPLfynU+3Q2aiR9NeK3b/3jHp2yArBUUJ3J7y+lEj88GhL4vORIiyGsUf6ZT
4phkLdYJXAjNHEwg0RuTzWT9R8uQbiwFzSs9ScmFbFllW6+Y0FqcyiBC8gmiHlRtFCwHZWkf4zxT
EMm7x+jaxk8ZTxWNBPkJe4oLXtugKTp2h78CkiyjoUa1Pk42vAZ/vowc3jQzK+LAtARUKO4vVcf9
pmKjr2aj6ERxmOW1tuoVi7977QSlAm0xHf1EZHHEQ7av3+jojd4jnWd0dVDocxXoTgg84ZYyQX6w
IYhKY2CB0GuoH7Zdu8UJHeYIuvIIhwSbwBMAoEB7sf8oT9uAf82XGWXvMVKxHqHzmvxiyLC19bez
mwLYc9u31yRebhM3vPB4q0dINvfm8KaRBtx27lb8RMP2jLj4PvbU7h1XGBLsej5/BS3Hx4FexjWt
WqXjjCZPeC9NFKqnwx1rfJJO5hxzZ8fePnewlsFQCa0w0OR5+6KpH6kq+Rf1qSlcP78bj17XcfZV
yDYRKfi+YfhZF2AnI5/6KfrwD1HFyrbjYtp8zWbZQBPoI2KF6z35tS5+vtoHLK3mwvkOWretwTct
DU5t/4QhNSfboBhX/v3W93dkfDn6NiHfs0Ydd7RJcSryyrgPok/Ni11y/1VuQDLTliYI3fW2TRpW
IfBkyTvF6SZfFe+OjAYeD/gjj7VLzjWpLDkddzvjhWosgp5J+X7WfQbzhnbj19qkEpke1JAaNHo9
akT+Cm26uy3IbchfC5ahnttUxK3wNwgCwaInlcMFoX+GnSXwbRsUtFYb5BWIN5r8G+SpLXcLEXHw
U9KTcsGCxWf1UtAFNHtzrN5l07ZLguHB2Emf5YzW3xBlVf2w+PhMUl4Lab67oPs3u8PsPzq6ElEl
Jw9hXwud4yWZHcCwD5yKOgNK8gYNBISdoU+zWHXjSPDepuCXvUqJwJvomhb9iH0ag/5JaQqgwUHK
qs2DJyrDLvhS3crKKc+T0lgqm0BziuYTSienECbq5yaKnF8mbI2ZKhhCBp+lblViVJVhISJ9gi8B
pIGL6JJ8BiuMm61F3e2s0LT548/wQA2Rh9qWu2CnZVvrM6qHBNmC8UIHJeIu57M4JPoWpXlqoFXG
yAAq319yuvZNMP2Vr0o5nib4/tdBIfcXtyGmCTunTgp1e5Lt4/ruH9Fqzaa4QDaxxNJ6cYmdat0X
gzmYxLeMbki7s/qozXdhRDddYmDFilPDvQzIYT+qMq/Goo/1VZIj3P3Y0NgDgXp36bLf21fKwkVp
oaunh38fTijIc7tUH+7Da0Z/+GXfxcg3uTrTxYYqwGNu1Zc1U3nCDsVe9L9yxCO6jRPp3uva2ox6
DPdPznR3cCdmBa8ihFGYkiTSrCs08QhBv7TKMl4r8El7pnJFAi6dsRQqXhI02TIzvIE0DsIq+3+M
YSMZHctSXFzCcGNsYEiFCxjps4cd1LF85YdjAaljSjl6WvACRDRGkuPmTkWFO7aAK/ydW7Jn9lx9
G5npoO424SH1+9H2hY7rI4q4XTdkL9sIJkRWGKBOBNl1Qfn4SN6jbZJi1S6+QlL5R47dwJSz2VqX
bBWpul4aSj/l2egSSR669GVXuZpVIfI9LDZfXOXzqXR3ZcHhfG9eVac0Y5HMqKoGeOvOEPgOzqy7
UMjjyNe8OkLSlQoZPBtesvpG/AcwTcbVaGk8t41TF5pnmYnUDrDalO/zC79RimD/BYLDWcRPo2eO
ttFD279jWzWkOIl8vaIqQoOLik2cSbWqpxIixtYvU4Q7BhZ+I6Lv8lVmUBCY17MNxxZ9GWe7KEuZ
a+CGuAo11l5qamlHw64qMKzDZYY5LbSpTbRbCG68YiDiFTvJwKiauypnog9cgB0ooEnqWXppFjOn
bCp5DHNiJhtnnByadheUnYsEEEKDM64MTDCgPg2846G/+W9tDKiy7SZW/p/CuWYESb84KN4DqUpk
neRJnXPGsxx+qRbCd3pOvWkOJ6J+LuyUhnqdMaP/x3MHgVozHsYmTXGj6G9v/WInKxmT0n9pJpX4
9mM4sAp+AZbNzCiYFivmGib/Ei63NtikWId3PmnweD7bBgj6H9+EN5HtHurPFf3chnSMhj9Hkbjp
0vsREz6KaJ6OQ4Jsw0Z0Bd+ioarOOe0HvbabyNR5NEbgKGlSvXUCrZgmgBCjiPgyPkRcdj9EX6P2
TyvBryc+7imhZHK1jnVo9x7K5SV1r7nf/gf0t6Cimx9hUDS/rSBxWNeBZcEnWVRK11e/tDcQ4/Gm
4WmF+NpoTiPeT7Jem3bu4NaSAof+QSm7Cl2BUJ/iuJuivA0vnGVjdTUtKPf/eaNWXGTJ90JkV9by
3esjEaHWT51Eo82E8D+6S+Wq2/PHfOzaJXleoQZ/jw/kxQ/DrW8t3Ur1VX6AfULEr9Xnso4G2yET
zH8ZaGF0k2dBuKYjveuBaYCd9BhJksAh0uYlDADckZUA3qEYqhbs9tch/FcCmyuCqmV/zwwVV/nE
YOasVg9JEX6TEgHZWwRBttCcE+mzZyjI9lzvABTiJ0fLvio7aD0GA+3mDmKSyCPIAnKsq5nx4pY6
Ozsb6hyC6v7VONSFp3akXbsIJ5Do3OZGL3W4mUpnLUX4a5xnPM52zUMD0PmoFRfzKaQefQR3q6q/
ZFll4/ydgP99Q6ShZh32bvMgZXjp6gsikuruIpVmSiZ7OPwceDw9n5AJZdsD7B2u2J1DSwfkoI3t
zy292TUtlQ34iNQCxksDEJ0KipcBfiZ/x1t/HFTr7Vg4HsXgjGZekOWzFGl7qMtLLoum66ZVh4XL
Sr6k+HmEyop5ODZTkdwKvjXIx9ND0jDUpusXd2odBST38oc2pnbh+oM11xdXmH1mI5rlrB1sVzLp
N55aFjvSCn8Z9tzmheaRA/j1hy8waapQAO9pbsO9jkVTzeW4JrHQDzgk2pLT5Ei4UZYKKFlBoxYs
mjaCWuzfe0FGuXCCkAL0FmwvgsX8Ia3EiRVoo8aFBEHQ8g3Ey3/zinTNYdxnPeraq7j3bO+OLG7d
wMdJgJN8Y5BfpGKsJUMSNDkCAOziY28CKKr/fbsurlYZePJs8guKxaFXYo/YxA57LFShB3XLKSsg
fM4jHNQ5+0OAcakNEjuUYBVUfKPny9jhlHBiHNlEi7yRKcpXs1t9/a2/pWCKaJjWMPykkSlyoer+
IMaRbXyB8IIERm2fVI1T8RFWbkfwxSOm90Wwkgbf4OHH19MX8d/KbTRrsNXWPuKmkDUSRxwXEkKt
NGRG8Q8LsLyiz0g9Vu6+IBBm+SlIsoww+xedl7LaOd7fJk7xBfCLFY1/FgnEG1VFzeG3qquSv+mQ
DBsvg+SdmHe5/F1KCiu3cD38hdZsvYO8EXKTAk9WnRCZ1qpnp94/F3JR+ICBYk9661EC27vD78cj
x7Z3SqWPGqW+GtNlG96svVPmE2ozg/1s4ixsd6dpucansWeM/Yd2QIzJjMa9fjvk7TnMkJ2C0IlV
qjbIzdU+rmuXIAio2dSWmopf3VpnAyErmRGg13ICVoIOfUcHK9fA3AxdwzGV4KHhjgZ5W0ZwPUmx
/2bTOY5ccPRXv1HyBe6R9+j5QL0PJcOtOGKU3V1lpZ2h/feR6snLA4DnJGkasLKa2yoFrkwROLej
APNMSiJab/jfQ6Pv8HZiXulaY5w+tDJdjR9f0iedynqaJ3yYquZjPzX5j3Twlywsd63i21N77Os3
gP2BNLqOJu8q92lDk0uldGPQhXTR1//JF5HrEm78qbyYDKSkjYTPS6W6lQHl0Ha5/TgYSDITss0w
LR5ZOth08zXobcLk/KFNu46bRZcomOgaJMl473NHHucc3KamuhrcDL6jWxQ2D61KWv9yEIWu4Ql/
MlbUwDivf0fy9/HLJLvRddr99V32Y0sh9i3XD4oVusiYSvsetC0jHhUlF32/OQYswV1AZTySP32R
IHsY8Kh32oPU5SW1Bxb3lOC9zrRWxmtr2PEE4EQYDGI+s9EMy7Jq1pYiw0b9Bkc0XKBgMKtl2LMS
UPY9Xrw4JQCHC+nfMArjrQUEffmM7rOJoVvPCNNaZ1JeEh/uS+N+MD6B9H7NaNB4VaUOkSKNz/He
fTzHpozn2tT8YEZSjdKuTyqJJjbxILn5Ok5MjI7KkdrTQ14959wWeFOtbDBXq3hBxKDkHnSo1d6O
jtFSUMk7TD0Y7Xb9d6w4p8FZdAhuS3Q162kzA/xBoTn5DsrX8Pv1+bz8IpGIQg0IiPwinRsO3GWb
cX5KxmBC3qW89+hKhLuEOJcC2G0FOFFZDfnRQqtpb8i84w/D8HriJTR+C66kdJauDwhsD96tiDlY
jaL4rPf/PYkXXWBFyGXD12AZh/ib/43Csrxegd3liriZwp7Rxqab7Gsk5cRjertbWtv7A4dgn4/7
VfysUuDgNUfLErcTKsChjIDqzPnOaE/k57FtgLUIjCbv/eBbhOsFY0n9vMaAdgKgviQn0CfxyM02
0H3FJKPJttn4eBbfJqVRfdRCyTm0kb4GZcZzDtdCCJFseubAmds410fFs9yn+67g9ZefVDkR6Zwf
/H/Mas3Y2XWjKIsyd5jpisxBfjv/dMj2FABP/NME7XV41CxkM7Dfk19qVlVIqc9C9YzORA/XgKav
W/AXcY8H5v6OJPGlkEP8/78VsaTjiV60tdPbS+D9aLWtcv2oavIGJbA8EQpw7x6YevS0AjjMEGce
+52tVPjoBAJfhcMbtl+1gteMhR/4TMWVTh14wTMKN3Xnd+S4Np4f78GK9c52PQdxH2zHSrZDB/BA
d0yVajOGPU3xlndu/rOU3kzOWRBb3GdSvtU87BCzJltIZRX3sh11/BRUO6kUJ5KQb5rkmRbCNF7K
sIaymzIm8Azl51VH6Km7NgMI0ipsvdemiQpeDk9j1vlFOZ3aEVHhauszXeoSl3WCM/Af892Ao8BZ
HSx4QYLCesc45EOjZqdthIrWauxusKUe0qDTFlNRo9IGOrC4w/pPT+bFJPb1j3Gg5egEIuVSgidy
WEsZJ9fGo7jpWBA6vWFqQsknghQX74SebBZ/1tBwma9JprGlg5xGdCQNyhzxqh0ttNjUpeXpbLoy
LSSO7IESivKk1pGvYw0p5+JQZzVBVdakdP8VGJLYbSlhlsfD8gJ8ASGxYPIfT6AAXrb75byJmnxV
luMy1xhbkJlBSohZs3m16IxHgfyiWq5qUBdE/ezKyx6biREaYFdJ2j3ni+hgfJZFLzoUhVzgcBHj
0tW2j7HEU0akESISED6TUggSOwxoTieUAxI0g4O9zD+BwqO7FxZKCEVM7A9pxEorl8r+pVUHLFY6
HFw48pbKBzU/0jj1SL0QgcfncGoZcu/nyGrw/Q1dYAHZyIf3OVGV90LV9s2TgNwOn81yQGkdLHnE
w/9XpU7d0gDaa3K3YNO2G0k8rkfKGJ0IN/k6K0/htYYx1NC3UIPHi5skOgE+rfqJOPxLS+he3lIE
JsY/41jFbvbqV+TqBrxS4KPxB/l8Cpw3g1HtAj1YJpxUrCO3qxYzZEQMvCVA8jR4mMm0W2nT5GCs
VRdNf9lKIk/8+LqDolTSiHPqbwNuUv8RH54xPdNZnwRSRJVxrvkH2S08kmexgxmsMoRKWgtAsa9/
vz/j3w3F80rVrHHUjqXemdHqYr1FAUAYv7CgduzCrIIvXAAjmGKCuea4ew3qFesWSKihZmYoo5/n
xyH2i3MJJzOWrlR0tX65mHKs4IWKkGChmOkukKq6W7BYjEPm1hhq+E25OBQejFY3WiTbmzG5ccu/
702OQfTsC7t9U09Xo6XEi1l4ttGvbXMDJWupLgPx6dD5R8gfgchdsDTgZBmcH2JZGjkiCgTKrcLE
NrbtGMJ/LzAO/u7xxXjVJZtAfn/kAJ2j72MXzzwfVTuVeCRwJQZGXvdcZYoU4kvUJt5hHtoHWLxR
zFowzCrjrnc8974kyCd29ce3VydhEL42prHO7mEAT+y8AEocn8ejUoi1etCzjtKDNwFKltvxTWr5
MdcBm3hBtkd7U3kIn0XrKc2iDvTOHOYQaJBGKc/rsGMP3R92EyNJnUuatWmS215HbxYfjuYp6U9v
da6IpZWThqDhKfBr8/HNm46OLjWMt97qV+ejNxK2VLAGZ6oxnqzXDT+OPlWLTN1J3zBuH8ATCXSi
EJdMdudIux02/4E01pI7NtoayomjdbiHXVXe2w9Lsu/9g9e0NzCzbSjsrCyv/LhU+Sttf4Wnaquj
+A8u68Kr9heoVX3/fIQToBU2KTPBvB7pv7nORcqoFaHuxUEDkebLnwodYtMX7SBqNiPbyTejHdxe
/A9TysJ1VKCbUZYx+6oE9b13s6sEofGjMMpY2Q2bBNAuWqgEuIDlSdNdQ9WIbX+FhFtLtqEC4nYm
bzgtN1iurSN54Sr1rYYWqH4H1qHLSly7sa8a1xmjDsK2bRE2GtpRiqhb1vCaZyUwIPGqA/wkSTxJ
sOQ1stkWlmm4GhrkJjyXNSmNGyZ+z67O3lawij0EYKuK2fVeXPri6fejhQjaXXSsBQ2B/TLwKX98
DJANfgj+ndx8uQFv1EIQQtSSf0Q3suUOddZM19whF7fpwMW/RsGu8YEQb7xALzJYCx/Rkb1RD9JQ
jqlZC48G+zt9iK2TvtUFpRYGY6dQTlurbnpkPHALeSrGqKAPiNuh4ticOOPfkZKKJnjruEG1RjeO
cdcPebo+H+hS3ijDDg/ceMHv0vQYz+ID+p3oi46THZyl23Y9jZivAfeRKlFEQbnYMU/CXxYIKZGQ
NY/2Gcf57/uqoDB3mvpSSSGfGFsEppU7sXr9MTD04LrPek1GL0Y2caEFXU2xj8sSQrpUhS7X78gm
H9eeDQKbOge6DTtRPOnmMgEaL3EabsUeo9h6mipDpP570fUBnWmdpKyRj6K2c7jvUvdMFfkNmIdw
aJfEt7DwqopJ7Tfb26RM0tWtmXdT/t2svcJGmiJmH5SLZNoz1ZZWVVdmcL8c1jUBBbzjYwARZiBD
4c4TCZ1Kgl/ozskFgIC9lf4oibuAWgbkfI+u7fWgy72csSuIIYaQh05bOZ9mZ5SpMiiz2PdgiQXN
547oVp6U0vlcq5rS0R9rgU4QHLYhQM6jtDHJskpkTV86+t/RtjmMIRY/t5e+W58lSp5V6JbwmL87
J0fgl1jhscYu6y+9lqufuPT4zIC5zYuxIItwLJGmJKchF3FsRgPsKuU8udZdx4rdnG/LD7FWUhI0
jGvm3BK6gjkUfGMQeNllfwyJoiTSiLqhekR4ARmn9FKAzHKxnTqg+pRIM3mJoj3q3Ffx4OpyL29T
DhXRmOmCoQmE/rnUuO/iE58LfXsgrGUX41yB63n+bvN/p0JVLiYpCzAnOTWVfdIISr8j0z4QL0rI
Jf664uzf1zCD3Yk66vK3JqjEh8DvZRWXDS9HNpctvyhRVgljx9Y48e8NKRhAO9RYnkL6wU6QuRTr
BG+fYJfk3Ij9TxbS5gCCvweieFv2ovyyszi7ms76KZmzrMwcI2KY4dUIil2AvF37fzFxWXX/mgdx
VYz1+q0WEw/U7OQWSGxUI5AKj0zTnw4SFSuHAxOAqAzsQGbmiUWcyLw/xgocWCQm4b4IFnwOvkdM
tZs6Grp6HLtIwYhhP1wohoXL03rmhUgCd+jYsAhgjAbh/Kwqcq6fmqgSAKpSS8hCkl+gFYhueeLl
8BFC51LQS+QREc/WBkM3pMN257zuZCJaPnWYzoUti+KyRZigXbsJJHgLoTBvYhg6T3Y+GNooxYGt
AsAaPq4U01gDaFSwjXMgXrAdCC2C6oR8w2fEV38FjxTQKmbEK0PeAmrAC2bApFh0w22yp0VN+0k9
qqJ/ZGg7dW9eLzlWNV1tVKBqPT3wYE2dCTq53y2nVZq86FJ/QXZW7qTanZgokmaLJguBHG5swLpd
exa015bBUV90aj2u/mLF461s6p6WucFPy4f7uR7/mOYtvLj9olE5+iPagiAA34sn83gnHGXDj3aN
UJaVbXp1p1LSAq9QgNynDkzCo4+D1+DAVdrM8TcgMNDZbbB577W0fNXkvo9ciwkghVJWu+qCG8qV
gCNBCWAevu/qeL3S3g1z/r2G6ixlMQ8rW6KX9uad/s3pZdM/ovSSMFYswHz2ANY6aTMWBbfJtHA3
7bnnDjt6qoholFrQpeJnMAb1cQ8pHPvWJIFmuPlXLsmdFl/iIDdA6efLbpTu8aXW8nMVOTFZeX4o
F9HFwES8fz05ozoG62o3a2OWq3TCMKha5pG+70Cl2q0899pL+H3GS9FPnbFF9637jIyg+BUROEVb
AQrYlr9yjofvqDylbfcQlR+NLohnNpxUsMaLFH4zFiPrrWV1mu79Mkt4YamHUErARervQqSDCSYW
tPafALllhgIPtkGvUIUWrf6HTNfLGQ048IKnV5Q4RtzlHe7RHaKnSMEBxscH9SSciuGizKftPW3i
69U1Q2cZzrIq1ZMts5tnGt0tFJxmOyfPRYHbp0LUoVtr4m5+IGhdFIax/4vsqap2dC1p56PeQwS+
J0USGf5rI86IV0DrLDp0qbuz+837X0idYNo1MblckkyEJZIzavl5aygjo0FLD77lzARTDVLk/OlA
xf8+FQot5fS4lIIx3orolAiH2nlmaA1W6UDCSSFx5Nba0KLg8UXhJlLnCYSD479kF21+axcjSRvR
3cIxjZdzoH+sw2gbQd23ZILUGAUGkKeXTYhoksT/5beZZsvfV1nGJpl1+pUxmkTW1dafpaRkkKas
CgJSFF0gNqKeIT2yLgu4c7iSSad28RvWnw2NevVz8hK521pfSyM8N1r8EOwroHv151RbtjghRgk4
66q7fNnFU4HkHNTcfwdD9Qzps3nBljhJ7sBjcvLbp/KUGOlT8AllYa1CrAB9xgj3BNOckstC+hJ7
m3ALSqnn8I2ZWj7pUWExdVNQ+VTfjOPNdpnilvtbCo0FEkTUePRIHW+UwxvkzPHvtncPIMlZW3H0
ANiXJ06gDAhTOuoyeIrJDyqwLAKYsVv9g7bII5URKygMuT/tEu+WEQfpZVXa9vVPRaLbuQn5rEpN
4F1HxGKTANOIR3iMN7Gjm+EZA2yNUyhqiy/xr19a7AhORrSsk7oLkqG8aSgzi1nUbnJMb4kVtP6j
RBd05pG7xp8lqWK0VnNdzJoYr10gWC9F4m6rrJoWxK3+csjEYAO8JATY+DMpNqaiq4WdsH3lEWJb
ezg+/hr1Y0a+mamHKBg1pXju5GNSyJ6tSPoli4bc/lJW9P5Ha9TxOTzeHsCVitQXnvLXWJqmPy3r
vDZ/HaqLgV0971jbbpOGMy7sgMwZ/xT1Cl8b27gXpnod8+AAhzsPEgHT4WcCb4uh5JudONUZkm6J
x8WbD93pbj3GRIwGPEhcUUJHI5xBl+rzftHcw2aqhD2rV1FwOQo0Ycq4eV7RvIhrZ+hBifilN685
+AZ2XC9OooR2P4yHmNoyoRoqphWjJOmsXJ43VksPDLBUeAE5jDBv0TgeosB7BxzoZSzqMhZYmM09
6Wil/0p1q49WH8P8NjGnkpG75WD9rndjkEtdlsGXTAL5XDUFbMFowU9/0247TN8xKVAVaDnnAHYW
2M54Pag9tRZ+G6n9zXhEHOPFLhiAp0vXhXz1EVxzXz2TkC6rL7ytshy6hA/iUS2PC6xcd7J4RpgR
MkHCHyspEFqzVd+cYBY8fPOOptMD5vT0BeSSAZ1De+j87uvxTkvOoOq6R36m8Z74jVexJpxKrfzl
vhBexfz2ELNLWi5d/aowSPhV9fJ/dFSdRNnxbih/UvcgVkxSCVECbJ3mVHWNXUzT71ZmSHWIRBQ6
+K8kXRKIUeDdk7RW9Uj4s3ZVrvjtbAjieUdvMrm4Y/zmq1KL77y7UU9L3IDP/t7ypksQ+XmceKwy
uM/EY8/EUKtJpDSTSD8MdlY0Dik5esXlgtdF+cPvLkW7o0a4y/9Efga+a1BpC4/j0oJBWJ9IJBQq
iGiohFgXxN4OPR7OQ/RxEw2SkNArppsYRrK6WdJy/nTxcH/8/cDSZydGEeqm65jXurGIlJ03aCaH
ZFIz3Zghl/uHY6gyqySmBH/oXXDgPe0CuC0zc3vJrXb7jIJkO8i2CEBj60uStlNAA6NBANb8U8cB
bj3z61xuxeyYQftGrh0PDmjUEAN0+Es7/73O+ju1GER1bBurDDWchpolQ7tn6OOS964p/Ku/TZ91
tWee+IBDiNlJmymv1HPOnsdxQtFdvZCaxU0x5MQM354tcisEep/xbebK7SR3ekeMiQR3hg7VdRc4
0Un1bwQihUEyjQrCJ6ccZ23OLSdhKwHQ+WeSQPIga+DpXKUgFy/XiXhTrKmOCyDZtyqKjAJoPZ7l
AxvSvijhOfAP+VPZl9wNK1ub0Sxiu1wbm5Z3/EVLg5qz2LFrOswMPz5wNuinVr1COed5wiAOycR+
/qRWB/iqsH7tkF2q6Q8w0wbovIoD0Cpv3eABUL8eUtvRAcDBMZoP7xLITglLEY27NPr0iu9qiv3s
m32BimwN9mdZU2bGhphxv6RnbXBqPtBHp2vAR/E/zjDwBhh57qqU6QliDbgKUhLaN5JQ/aVm1nKf
5BK+jN4zKp+HrLAxpxqz7UrXbDOdC5+WEk+qKnDxVVpXhXE1uIMQXawXlS1j9QOAiayi72VemSv5
EVGLa6JRQo1AX4L0VsoC6xBCzfkOuUUehr5kbpEwNGsEOprqtTiPUyqV+Snw4OKoR4yNnq4NfdoE
6Me8F7RjDj4i2HuqP7IdbLGynDC/zOZbqBjj/uutjB1nF0e+vDMEe0uQO58cb+LlSeAByy6bjCtc
P7rzRjNKucSdRuGE/pRntDQEORmEBhcqVaS+2vG8+55Q1e+C+ggMnWn4irhSPZ+N6ZSId33Fv2jN
wnMlU2+BXP07AcTmnJ7P+zjR5kk6ETGd7KHK6HaHfS+JEENns9K2CE4gxVbLJ8IKD2YdLLEXVrvg
JO/NUn6vfb9v4WZrdZ902amX0o++DeSztQiizlAUvym1SckvNxwI2GrO/OboLrPvqczAd9tPl2MS
4K06lcea/uFXcAJ8yRbxXMgy3RWM+ndbOD0f3Y8sBODzv9Hf6NA/nR1A/EMdnvmyr7ifvJYZxsLz
qHjT3xKfX9Hee2hqChEnkcWPPwtX6WqXeU/hUQKuuQwOIXYZf1iIl/ahptzN4eraFSTOzaYcD585
/30oKondPERE5L6X9fohJiPyqMqvsq814uAhkfA6E8ttFj7VJMZiXk9lP7S7gAz0H4I2jfa+VRj7
Tnj/B0tnsncolpkeGLutrobRdntnqFpVF+khXhODwifneY3SeCWDHTTc+w5NClmlEWHD3tv9kNYE
iNhLm2eUZiMviAU4eSEYD81/CIwzFCOsaGUy00YCdHSom63+cNYZ4g/Vrx1c922tsGguqBhbFJz6
wlgOQ78/YoaDw5GwifIFjLOGesuLmV+9T0PY1P3sCaR/8cVp+49Ej4FVMQuA9yLN9dP4l4rOSO13
eDH7sxCMp1OqH7n9Qs+NzLNSI+pDUGxmF5rEDvgsmtal6tA5J+HdH3kl68alu/elpJGA1TnC48gQ
blJU8y7qAgiMPdcHCRoQt0NhhXY1a4iV6fxCOwW2eyR0InZnk8Un4zIvgio37uMEuQCWB0vkxH5G
nrfBm4ujOs3xhct5nE/rObXiCSN682AXszZbz/1SLQItTXxm4ZFBikhO7ti+tY4XTXwxUye0Hwkv
++9mNQv+jWT3dlWNU98fEn48cOWZlgWVZwlZlZbZOdUVO00D4tUsvXV8HKxNRYkwHK+EhFETERYe
+EKkX/2DBePCU0FzpEropBUh7glUmmSvnLcnZan1XdQ4wnl9TiUzlKA+W82K+3ht4pNr4Nf1AwKn
jxVF7gN9ZmSMZ1Wj1xRRNC4g5BgFkGnD9vB1fKJPIWfFTCyEWukSsGCJzfNoBVWnX23N8yV1wW2E
Vwr7dkYmok0RAqMstX0sIs/JTd98ZjpsJC1Kipi2pzgkbtIULQn5s6YZXSxR4EQ/VlOGIKFbpFF8
N8b0P4CFIS0EUEv8gKQhMIBpQHX4vS8+QRi3Kcr3wlzbGqeCwC7JKN/sucX2KVMa2pEMDO2wUv71
jdd2vnYlhPQ5Lt8AxIlN3oNkUSpLmA1rDFnvocVRD7ezG2umNmPrTXX4OKKscE+SoD0IYCgqKzLX
kzCDJKiNXjgU/mr0v4CtE0LkEXEjFFDivfCvz2TC1vRXLJmg6j528WAjo5O2o0vuOr2IIFM8W3jF
mWmL3O5Sc30/11eC3wbm6DOIb987j/2OPxcAacT4aKGwUTtsiljBhsndKmYSj7aQ5bry1TGmn0vC
w0IGVoak66A7ltVwj/U+8gyJXgXIds2Y3aPJAgc6qYdJEENnPwozERZD8KmVaGCn+jjxzE9C0Fee
qxI3PoQZF8D+Ea+/j06X+4Rwbx/8Oj/jqfLjkwkGt70734e+EjPdhP1FUTn66mIgeoMXWGK1Vnpl
ieIbpHzlWoPsiIqphavRkf3meMtv/h9OXkPgMtCHUBpiZrcbqkOn5KYmFhiLknyqDo+U++WYRtzW
WJAMQG8bnHqYNU7w7vTRm9uq0/GlcXE8uoyDWM1TEIM1SzQ4gXq60rXBnLINj06Gb1/jaHsJ1SyJ
LOppesknhoV22mj+IwYOHzrJrhvrB09x6N5aJl9n8KJ/Mqlysdtzlo8z9FE5qncDTVcbpQP1h7RS
5uCm0IefcwqicNQhpOe16boLRFpvtnMW19gpD73XuNVPs0a2S7iO52cTWJWFcKP2/EdeJw4a8q/N
RB2E6EiFu80Obs+TgmclXemrzFyXESYUC2JQYoAuUdE/vKHCvhqNou13JEXi4glE5nwPm4jY8HCW
cmwcQ0Qmldr3L6nBudzOH2PW5M8LP34xBaZ+hwKqHXC3vghpgcoLrdoQo1z/MG+/noWHoR8J1ui3
mrR/49Bt+F8dWkgmwHxOds/5GiTVcmk9tr6n938HyHGYzG8n0fUJ70XpkiU0I9ySRMb3lFjJEg2k
7Ew0S6moGINaEIqpzWsd2KVmZ6kYd63gg1jTRMRnVKnYS/Go9737AVq70O3iTOdb9EzLK+8TmXIV
FaCSf/U6zgbCIRGbdL24yjFgacIBgtLzDcYiVKW7W4DsE1tHLzAg+XCuvJScpjVNi0xk5+kxYCfm
+YeE9MhEVuzBKDW/Tq4I04wEoALECe5Hf3xq2Zlyg6sJ9LpMq71TN29BMZMgRFSdBuFfs20LtWIS
7Yk6OByhU4K2BLc8atlWVgRscqBARYnRahswNEP4DJEELd9rqBAgza7/q2LQZ3sxVVxK3wAM83A+
Z+3DVgo4dZcFtvLrkNIiP6m/h5jDJX1i8i0H8RWCGdhBk5ppp7DXWn966d4ZYB7sNuKti1J/yMVv
g401KDsbLz4am4dxTLgDSpTIQH3V8UZHISpsiaD1sR3iyY1Q2jhPtd91lTC7IBGOK3+hQZ7FffM9
IwwFvnfTpkvoEUw3AwCBjRD1dD90NmbaFsnWdxlpvEGXHVMnGQTEw2dkQR42mcmnBjVcg1J2jH5l
b4tjGxc+Z4F378Qp0WoOa6S0co9IhFpV7djv/rbvsHICWrMQTiuDJmqkedoe1J515Q85g2WJprhT
ERLWS7JkqtuKW1xkGXLH/UUZ1DfWdi1pUT3XobD0r4z634dkvEoXmaxqQGAzkSjA+PgBWKf7t7bC
+Qi63548MYz8f6Em80xEhZGP4o9hpPI6iy4g4KOTaSvnfMHxZxjI2dqgwDhdz6iAhB/RjSrqt9Si
I8uCYuiIEKOwQuvdDGm9Gu9RVKUuIiiQQEu2+rde9zb9pbxTJheH1LzQT+mn0pZM0WbUoZjiwHOG
0jMx4k/jAPK8PbU9G8azJwuQKWbZh8FcVr2Yp6th766cyBUM7rqJ0bQECeTXaSRknsoQpOWj1fE2
T0yZ/eeNG0W6cQ2ZTNOw+RpvfQ6LNmg0hCmK99uafXly56q4+wQTACTTHqp2diT8LRA7IRdzpyNE
evWuHyGxmTvSJzvI3Lc4PS4WkUtv+cVBCHeSIQ2Z0HYfGNHgnhdcBKtPOaDljpuisUF+FQIeClRF
W1MvS1PoSHjLxxClJr7o646xMt0qzCHmGK3Ef4UnTiRmYuiliJXKCirggsnblibUttzTAi57BLms
eIvxh0aqVfRVJW0h/+6KbSn7C2ijXUwfro5hICBxIpP4jtK8yCFKlzvwu2sq6MZJWoFk6IyCTjwi
Gi+fRNDXiy3RCLQb2cEfHa05NDAgtxwzGJsLuPovU8cJpFTZF3hqxsjEAwpK7/KMAokMkgMYXz3k
73lKOgwewKDr/uQXaHxkmmWTw2kIpiM97DfmD0Y5/PUJkgSEtWSeuHiQLaxLY+jiVPUaTN0gmENX
iYp0g4TFGcRRSe3FQKAEoh7ouP/a0bRouQjLjr2ytxCFGrznqnxTiw7AaGTWuypwIdnYTMaCP9QO
ZjZURA+eE9qMAAG/sZq0u08LF4Ti+Y7AgqNisa1gJ6rP0fYz0/icLjO9oX5+isDIL5yxWFxPTUxN
pmb5ppAiRNFQtiQ8/9G/rvPac/audQvUOs/gHikgD3DSgztMrMen4xXN7Fs6XwwdxG86MO5KRw1H
C3Ae/KsE1crRki4nlPVhd/ES/8i13az7LA1Ka2cQBHHDg6MCaGqxikLrmUEfDwgLCWkkxHod2aGP
0HmA/zQVnvUlgnsUtQU0X44BU8FmZ6Tns5p2dsYP/XxCjekXXVYZ28cGI6K4+besVCYCOad/dkHV
HdGxELA079Tj4+qYruXzQYveiDxOOANIsXALzhTGES9/Y7kr8GlHcZVKYpfEeMFURtPvPJbEERRJ
jHbufUcytl+ldXy8sY35ivzrbjHviwvfz319yLds3yYOmFmpDtZkSGm9yTbW5h4+LqQSvde7ByKm
RpPHMoxU9i21b0aRchOyUWdXy1OgJ7fskheRXTLyFgtBwAo2vvraxfwbog8Je1razwN/a2x/ohTA
nuAPelVmyoUJxuZoFn+7kCdtlnMS50PkZ03+Xv3RGysKDPjSKmvljVnrlAfIVgN8q3x8wslxYSI0
KkuaGJMAFX06ux571TiLqNlS7Y/bWmUUnYG/Bu+toTUmqkQE1jbfDr+qU8kVrmJJYA2ILnoCfIev
FVXj+63FVmbOc/9t3hocikNqc9dn+y2Mq3aVgza0xgDtac4o8+GIhoukxPB3RhLQbhhXu+0yj7bE
/0Yv0f4DILEAEJBEahHW9zeAcnKh3CmawVkjwSXVP0/O8qrHOx08RjFxIpybrxv1tf8g5JG7wdc6
kMqnMfXdDPS0BxxnKmwx0saQwoqMGsFJQNTfF8H/HGudQtEffqnelAuM8dNX7wVE4DesrkCqCrP2
eEcYIixx3JHR5wa3qOUCN3Uj2IaJzG24xAzJ3cIAIqw96Y10FOTcWKICW90R3kzHKpXmIsMJXdEv
z4Mph+JsUhIJ8VR7RUkvV+DcLAkhA67SlTmXpPOsnkvGNV5TtzEFwZn1WvIfeNWEp4MC3M2sDN7D
VsfWMdKguH+9FONiQ2NDKxXiQ5fseNSJ/Wjaj+MmGgEzDz0Gg4qPD5ARtXYB/UgO1wdb/GThzan4
PbRPRS+XmnTR3r2/Ccgq8SPr6KYXtGbe+1IRqKlDPP2+BzO1y5EHnU4jEFPubo2vZexViV927I6x
UeRQJO6E/Q5B5Y6I+8jJg43b6RqcD3Cg+5ChBmjDdJHDf+j+qmpV0D6nNBt/r67bC0AExYo8hfAu
fZsqz2K6YUMSk8RJvWb7bZcBMMt452vy3uI2/MYbXIZu0D7UX4Fd1lxrhiKa+jionvYXUIhFeWJG
Uk+lQAAMqbDppPcK0CsppaN9Q0b3+PjtRvd6xk5YI2o1VX/YKlaibxvPJc7C/NB39eDlsurmbDPN
+hzglDqfTM4jZKqt5bgMhF4oI9xzoAtGqzebkXBF5JCiuqmmV8vfksfLH5Dnghc47h/10p6XtqXG
Ml2tBWiuomu300FT3eLRd+w4vOR9CnChYfkPrfgUiwZ3KKmxKGeN/Fhvk5hig14INZOwGdWZlV71
kaWrSipHcBzX6DmnL2YqyRotXoXfIeDFlebTSiCbQs1Cwt7a1YAMKcnIEYhR3Bn8ujbiB9aid9eE
y4frCSdr/6iwgGDtEdOpE5Xge8VmJnRL+nw5ee30jRwBLg9Cj4UYu7YIB+EOLnFn64155QiYpmnH
Z8CAXWT0KZhinAFcEvCmZUiFWbuN8sHXA+5lPfV86LP8VYSEW4HK2l0YNkVq/NsNFGd5f3qymgtC
43rYQoCBFATL5k3FQW4zWl6qqq8cQTeBSCwzevltwGsKsGIWRw1krk+j31FFlGqElMCRkq9KvrB6
cPRIu7NLGNMkdXjflaXA4SFlscO09APaQUdxjyEl2/3SZZrLVBljykeqsl4glbfjjiT82KIhVKk8
OKNdy4kc0HaunBv05PI5lFNYEpUjiRrhtcmaH+mr0uX/+3fv9y8P1XiXvzLirx0nfLkbe+zgEFWa
NgCV1lBF1tyByHyyAgZGQyq1ROCQRwr9BhdAI4zzdIf29QrGHcX0vaTgEH73zf2UPuONE6jIuYXS
RSwiob/LgC+NYtcLriN/lAa2d71BfX/aHSBozV4mNNrbQn8jyBSe4w4R5TgKw0l3iUdmxwEe42X/
DL20WYPLh7Rlhxhy/QUpI980ZSdAp/d2gDGGIjbYX6DjWEApj6XYBlZv035fQJwCXHzVQnHkqUjc
BUHe7llgN9PQeVDgEkLPN1TCTAcPPYaOe2XSjEIxQYurhY/cslt7zcT/o0WG5rjSFcRvt2XjZTI4
OYBwrrHymLuJ1UujPutZMrR2Ffc6lYnZ7daZxTPqvMoJTqevM5yu11Nbpp80/oWhy4SQc28Pzco7
MMIPEDZ7Vm2LxHnMqQYjb7jJPMj/8KuPYkr9UtIeqm2aCl8ZAUCHcjV0+lf1dId1TbnaeC77bMxZ
KtBe0+mpx8qDc4YI1NmrpuUxBA3Syr80RnlAFfwFVcS5wK4YkQnES20u7WmYW6K9CWhOXmDaxFCL
WRZ0HyMUx2o+mBBcNvdmpZ7alrZ7OMUsSwZCP7GSF635wsz6cWHnnvZyNqAaZ2Kf0POAzsmPxM+V
eFxQHKNTEvgz5Bt1Hh07M3Iek1MyiTxbCo2OXc6VxAfyNOSJ1/supgkQizq6vYURNW2arBManqj1
5BnWmx2HOfJ+efaQDTkFDCLnRAh3c+wIN3PUrX71nPG4mV2qEdMIEQ1R6cNNGd39Wj3yPPysvYsB
RJeY//BRoU9B2X958oX/8O0CvUI8b56mAOpheg8oq4pHl5QwpRs9Ed2jL6ClV3FUsiIfYunAs8s+
+Mf3BQ7Tup3p4IU7SXYYgVZ3ZuNxIQRVqBSCxTBoDObmz08H4Gk852BgR63DtribH/LujUKl11Eb
HcnKKWhLhNY8wJ0rwMYE8pNTG/xN24WDqxG8PjL28xEfP8lJWg3pQQwYYCxk2FGRhz7wf336cBTW
WToKhPjTYsCTq0BNl3QlX27Jo/NmIooqBMEOySD+Cf7ei21McBiKjQs+z29H8GQAH3JuZs4mzWd3
EooGAe/AV0aC0yuM+X6m4E/gYIFYVY9Gmu5MIGMJk9+QhmWkjwKYskKKdH6YWM37rfP3rR92Yj2P
QNfyDpF3O7qrWruK83SgSuNGEgxSt1/QDXV5NRaEBEBgVooJ57P8P9pvHABM2Vavc6MePZmG258x
jOKm0N1Y0kqU/MYZxgnn+w8zCXsbT+RdJ7uVAb1VruCseCAC++IcItDkJAVTS4r1hkn1uqpSyZ8V
4+goqFCDlChahYiFWlMtHpJeLlaq1Uvc5s05L1rB5n9YqlIF66CiQmNAKUl5qpshWuWPg7eHlvh3
CImgePWtiuxhWXvgKBM6zZ7NMRvdNuPEMJaJ32kCutYuIXThKRderdFUYlF117X2mdiQr6uhAqaZ
TwVt9Q1Go3UGFHkET1/K2Wds61klnxDL0L4QxYSvsUXUYrSZKbQwbg8KVPfxbxWfs++hcwYBa7t8
HeruvQIQlRrFPxSNGJYz4RXG0w1YCPyoGrwtXe73+djpkROv/e4pvO0dVovQT448exBNQ5v9aH/9
E38oabmeR5hgIuTLxuJCheLvh7Kkf+KvnhFhSEzFfejC+RBa2/lnL0s8baMwOMs+LWkQVIjMgw70
eoH2AkCrRMcWWGoN5XfxpmWwMZG08EXPkJbNrPGbsF2FhYwDzwz0QSfrPJo/Gma+SM8luewwd2DU
jK1i9IrTalrgXC6v3N67em+o0luBc0oe1mZlA0ZllMqL9RJKOYXe37sae2nk1eC1Wen2RQBdbW+C
dnnLES+jU8t0xeiA989SeJQZ6rDGFwjWZ2cPbbhIyL3lBDObIJ0PZawnh9eLHWJtwgBylBMTC8gx
mHy9EuWK1sHT5UFItMLkmxoh1Ac1F3clN2fN2ZT9GdYHnRtZe5Y1SIDngxuRFTYNnWFjQWyRRPZJ
scfxWCGQlXZQ4O9t1j/Y7NMtsiO0FcrP0FFKFOo8W5JI65eIl79SNJxJazOGEazxU4FtdMiTCPdD
1zDkAxsEhTyuBNSiT18mhDrUPublPkKsPqV9r/M2VIwhSBSHi7SCf8LVSqww4kvs1sRlX47SsOS4
eOqFId6a9KuO/v+bSgmQA7Q4FPujhIhLmUq99qKxPjpo2HmXsUfF4+UhmzEiKdEq9V0W0gj6hspn
B8CAO7uuoz2q8UByCzE86ArKaW6uCjaRT6rquOqUEkGSwWWX5u8kgebJK+ghmhKVw0hd0qKD5h9E
KTetKLLuUZvNUq2gCRhx4ubSywiVo81FHLs8JxOJiq0by8hnEWwB2q2XrDqrb0HdpKtmn3NTa5sC
bXgtrcV1kZzIjMXVGayWOqj77sS6fIqTNtys4IgHdaIKBKlrdvD6F17DLUjVea4YQ7OznR9yVAyG
HrZ5W+3Jt9ymOsrnXEBPEUODN6/PORF8wjFqq03e86pfrdsaVA6PSY3v45W3C3Hi2O8//1VTbrou
l5vbDCLSBujhOF3S+NXAu8CtIYf7CjbV43RF54f87Jz8ZPnlzoh1cl53Ss4rY6uy3mF4bmMWKT80
LCEhn/SfQdjRCSI+3SxSrj/GiPR9zShLW3ETNSSWiD3+2TTUUwcsP3LhaBvDS/MRCxRXuwZ3NPyv
AfkH59mw/iBBok7cQBvjatuetqicXNwcF+tYBS9S5tNuEdpRZvJGuq6vyQuAuhZatwecwJR2BmfL
M4u9hhOIvUUcQATBRtc6o/HkfUDy9/kPRcqfoyvCes49XdcofQ72+u2FFSra5LDhpxEg3zbP76um
PIHeZsQ2ibhtuEbceHQUP6A8GqZVfNDi+jb0avsYZs9OmC7vAEregyoYTL24upRJuOPQklBVVHy6
+DwlsK1Ny3/sRzycba+lHwi12kbDJfuWO7jPPSj1OEWGoGGiGoRnJN2tJf8EneukGKAwODYmqF0X
rXtVjYACacEFDYQRWIpdCbAMiz63BGS+01VS7qYZHHuAgFBiBhAGqykkg+e68K9BmgaASaRU84TA
Y1Fo4ruSfKmjArexgbBI3z1rD0vpquNVHqF4EWcnOlOR/0vOqqpkU8wxtXUVmUQEaep8V7zget9i
W49BTHiurWtVLuwuZMOICLnaYNxBULssHeFTp1hpYHZn07iO/azAZszdNcSFD1EnDaYAlvkvOSPC
CoVEmrslQ/l1bygYzEMzSn54Xiescn920NgcwjY6IwZAjHR63Lk6Om4Q/zBw/oulihIFAtMd9kCb
xGW3Mu5/fLopUNqFsi6zkVYgyK6r5ChzYQeEJSSzqALV1meK3zho5Mr6W2u16+4WnEaSUmxFwDrY
Z4TllAJLFf6N9n9EVXZAO/87GcMOFaYUGBCW6MJSjag/nr0fukphl4vyuSLpg7Q2wYn2guitnRO2
qWOw6vbfp70UgIH8mjdU1p0e1I3bVJim3kkoBAr5BCdXtsgS2YW7LkM1tlzOV2qwQuwsaNzHIOhz
MvA8Gzf1WjVlQhphuK0Gh1MANBsxjsrSR72ByYCUKO4CkA2XyiUMMCmWLQlplzO9GL8JnIimQZqT
MoRCyPpWQqQlGUXLc+NkEEIpJ5ulu0kXhEp/RhhbR6phzG8rx7kXkzRLrOTjBhIL+Jdf4Xklggpo
ghUw7kw8Nkl/68YkafjZlk/GXTOQN6MEni4Gn1OyvSJd3Zf8vFUi9kinETH+ELP7ksuAYibNiDXv
GrZKeNo0uaUsCtUe4Aw5HP64fxfp298O1X/D6V6dsFrw7KfCxmJ6w4MCqp9Ywfo3N1xIEbxQNQ0w
F4v8xiCeODYCyyMReGV7/Vwdn2JnOlGlF+C/z79tyeVXrJlJGImmWfRklHSayq0NeeI5N2gyIwIn
Jr2VEsLdn9VumX1eBX9y/ENtT2J+NOTSthfRZvTLiErx7+xj9SbOsY/VFH4DnPspr+X5i0ASzoUM
IvYGM6oPP4gadL06cjXXWkDvrYnrzyjdU2Zb6e/Deq9NEtTT2E/jO398cX4oGw+agma1ZM3F+LZF
WaUHo8M3YZqBIAmhCeS1ngjx5m7/FhurtxniWOMoOgZLbKMxcQbris8mdOGeEdW4IpEnfThK4e1R
rbfm8Ppuq4aLM9dTsSvt/PO9oMwaozn5BNByxw+QZJ5RI556xgNiRuUmobKPAmIkMQ/DEZGXiWdQ
Hq3aZJM9mc0Y89D+LQTTHkp4vlGJ4693Bx7yh+c1oBAUQyc3UHYpG7RSYYEk7hsozI2B8MqfKAhP
Do9AQmvTTpngp2Z1pcmygW81n4l+bYzrQ+cKhsGWx1OcPAr0UhMcdxVMR0AxMBf/QmYy2LKWH2+O
d4NGkIPx9gzuPPOASWiake35WU2wmFmAPmV3yNl4Q1HbeGw5le5sCtVDRnMy4pgjPx+TIes1QROt
gRK3VCltipHp3BjBYedfzBmayhojb7rfL/hT1DrtI4wQrNkqiyfOMG0Y4P14IITF4yBGQ27yxgod
JEJkYyhpHOTX+bVLklUzwPIiDp2GBGnK1MMuQxX7zya3zOprIWgZcmmcqGH5mqcXOyla7z6jC0PK
WZcs1tMYti8OO2xY/6PwI7BTtkM+lRaZwjKeJM+jd5OzyhTZY/jJmGudsobgVELV2EAIgxbcTt6e
1q7f2i6mSd96fSva1JrMwEfF3O69p2TwjLej38GUo5/9Sn3Rt12Gdxa+WXEROthVQxzih+aNJiOx
kee0P87BuF4thA32++1wDOsB5QaGHNSj6Toj33nlkS8FyS7KaV0cQqS07vH5UYWftIHkvHlMK5L/
LeZM/HycqHwRvZK7gGYbqNxhJDZU3z+YQcX7PP36UL5484RetGW/9tcA0cML4qLdWIeT25bY7sq1
CmqIq0w7oF4pS5xOCxFdmKzJc5L5k825qt6uwHgLy+B/bFPoqOGPZr/Tfur2qyb8AypNFBp6OEdk
MRWOKX2Wsc3tB0MnM5IeTyJ1MbKbRbBAKddT9+/zoaR6oqtt+9g8uWSi1rXFqtOBBErSuEPWP+QJ
vaRouRrWQnlmHJZmKmkpgfavcY/zNMTBjxIlrWnQjOK3RRAziI/MQAlvE61imiaYrtlrzIhD1b2j
+gxLQXkBHCqfYzjx8BvdN9oQkOIxRuAgpOUW4TxeQOmkgtnQVR7LqizoHBVH/R0z7a4kdska4k7K
moR5q72DbCLzRHERaWEEHnrCMA4VdeaTynzi7UoBUwoA/kKLAqDPl4Y/p4VNMe7p2d65LxBPtoda
hzjdbCF8UoYtHfIwuJHBlpyVHdGTg2zv/x7Zdk73EeA4JuPEKu5WrS3BCDd6Zv8+qZUBwdd7A0rU
QmRJv6HFFJ/2Iqm/WajsgXvzc1zrXzFeohkwSi7XmayITa7lCgsbHVkBYTn+FEEaMCBd5vI1QA1e
f6/i/wSMl4uunIAmKl9ncuTaWsuEOyebVocDk33bwvzZzgDM1cOZqfcxQZN8nvPQMIQRRwo1N+e6
746NtmMQlRiGESGTBoobnme9jzaEGPEtDOY49BHxteq+gU0LSNHnDyKnnayJmO1q5p8iWW4Ftuiq
/HQizOw05mXoUIHTkt81OWLtsHtaRnqDS3Y3sFYEjGcnAonTb2ZLvxQKXOSXXpOnNukmiZW19vzR
kyjMD1qg6gj3pr83B3pC4qVKsRpCbYr5RAprJV5iTkIHwicMWM2xybacNkRP2tHD4fpgRRLg6brv
owTqtQSVwJ4bTfbJj+CtXLaW0d7s+M6gJLPDIFOD6BGy/a4320V45u3FRmbUNWt3nPxjPs71MO2h
mTBSmf4wf6ih7USq0biFqNlAJCnV8Mc+LUVSH/ZwPCsNbO4zwtxBekk3LxBYQMW8Yk7pqVSIR/85
keNf2m0oN/XLV+aWiRxJOvvNKZ/VQ2NZePUu9B6mJKbwq3Q1IBmLQm/K+rwkd8NHwXkZD0d7I8N0
oDYVq7nFChdsN9qYdtXdimp20VUTdiLCZLDwkoKv7RPsK60ypaF6br020iL0VwQ53/NmT3nB73eg
pmAb7bgG+2/7U0gkatnEOH1l2WrQRyZ2HEO4iTc4pKHpISAGjoory0p2Nii4dma3rJW8DbaXqIg8
DShuAO/yUncwLAFkHSoS9RO1wklx7HvrBq69GZRWs7l90OVjkaE+/heATV74TIRillIZWHGZgTR1
hdeV549JJSLsnTUW5JvnjX758j4QeTryO6LYaquLbcy7axncwpMmocqluQFfswfoof6Tuu1bqP7b
KiJDy7U+WD7o65eMEgiqPuEABiYJyU4+vAOr5uXy3J3u5WuquQd6IMu2GFPEMQ7QUBw0GTEslOU5
aRjUW0ZKYg9rHCJuTI96DfjZe4Yk1bX04PiqVBNsTu7IWXP9woKBuscF9eL+q29SlOcG4AGyJZzq
jsVuN0CGiN1ajHEj2Ey0HWNRam32OdBTb/mg1MTjFwYsVlNIndokypgrRrfh02WIA4U09gM7uFas
aAo9UWth6WPAbovXrW+z0r0it3e3BevTAlxfjZ70qBX/jJegB3/t/bFqFJspgewcfMpREQ+gTC+L
mzG1gy5NtLrG2SmwwEHc+O6ZbT5aLuPJlPp5AU06L2KmZBH08mpMbk1SOrKOmGclhVrRqHIEDwWz
siDs5Ek87Dpc6madFRR/X95TlJIQ6/XEKMatz4bmLWiR8S61DF/096NM9m8IeLCORHgz6Ln/g2s1
GsQ166br6k2tbbPwzXXrZl0zDXOkW+tOZzc8UMyDOUqsOrcC8KXyc2BdBL65JjoyvIyUJmZTBK9Y
4V3gLl8T44+kr9g0Ukgj78wLIX23POgJIUkMPWJYwclH7aBtFV6iTxu/QO2N+7c4/UyZPPXWLdWE
5C6J06GTQFa+5r7ZWc2oqIRRtH3e8yzNwV5Ivksmsq0UbaN6jPAh4XXo8f+FmWq0v3cJhtWOZeWF
X9rIf1ib3Y3dpOXt5qeO0pJoMcbKHLyntFMw9cSsx2FQfepsHLCYcVi1at1kiQS4V3X63E3/U702
z/OdcMcHmou5Rjbnti2u6X7c/6tnrUCRUSjutkdwsLMf6/9ne6XaBo2sKQbMiHbruwhNJJz7Mcxd
5hBHcsLDFgwoiNfzBAGjNXuvOn/aZpAKUolKGk0O4VsXkCzm5Nk3yJvGFwR9fC2Z4aVlJob0rOhT
XWnnYBzOqohrWMX1q0R7q8TsKPwxK3VuWSzXlYDUwVjy/+1VZHZ7PF7Fh3wKUW29XgNYmcP/Z5fc
izbeUgRNc8ENeFp7pHDrgg9QfnsV7TJJ6hjF7y/9IeAvYk1OONNDt3mm30ayXcGMu0bNX7z2fiEn
q3j5QXRq7d4fr0Fv0IdXZE/6t5uUFx88iiTbycln61UjyW0ivgJGrJTfZQn+xz7RB0J28WAQHnKl
FwZWnEAzIdjX+zpSWZLoT03nGgfKt8JupE2fD/Rl2ayunu5WaZuimlD95K3B0BBKYf/ryoeEmWbM
oQim8aJV5+YgAwyETAchGqcWZp5PkycEiC86w0KsVbLKccnOV1ZWwaRnEkq9gYz/1DmNy7ZU6a5Q
rFqqIvNfaW2nN4vCKGs2Ehntxh1Po2xZrn3dhIyVhdT3QA3qc1eZAodybqx3y7ovGrSHvoUbJFca
2u32wmMEw6reKEAIKeNI1nihtt8ienR4eE37ww0/6O47+wUCnrbefsmmN4EsFSYzwBsqyuP9uqE/
mG9tL1Nkq2aBzDVv/lECcBikpGLnEQw/vh0jYivBxb8wxaWJFJ4tylx8zBWtaJTITZHvDs9gtavT
vSuhg9tV4H0pyVik46yQDaaV3Ql3hIyFJDsKK2LelrHtquiOcrydJPwmyor2o0fed6/CKigknjbO
1Qno+rFFtLaFC3o1shiUxyy5t6C4giuK3OTgnzh06rgVG5FqKMrO4BPjj5cqJ0iP5mqPNKRgAZpf
d9g0Oihd5to+fH8XOqW2flxLxkLQv6ZxfTRCrZgM4Jg5zPWYW2IxONv+oLmBZxkyZqGRJl82tX/O
QmoKFEpwbSYh8iaC9HSw6LcS50LA6g5Q4IItD2NBhJ1cT9Qez9P+2TTT/PSTVbDXWg7Vcqnn2uh4
HWPm1qjRYTTmg+Fn/+IykhrkS3Ue7127Mz/I9pjkqg+pQuB4T2m/YWKF6BpsxTRjYhkQxRVsIq11
/M9zCmb5LNKQh4U9HRulIGve5CxFsMiyPGEDGq53bzQE3e/UlJRE6Z5/N7ZLuVD1N6iywiRUbpFK
J6/+DhT8RkfxGPawBE0lPSMKrQRUi1oV+8tCvBTTlWUxZHc5jQhCOAz+PuN23KzFrFLNweos0/BH
s+XX6Ve/YgUidBuHMNXFrIpnZJJaWfo9A88BeT+0PgmFb1TA4UfmZNxxsvskLa1UmYGWmRlesiMp
EjSkPW+w0/53fXnWVZufhS6mqHpySwf0m04NPCT6s0SnB3VnH8BZ1mZ6BgeulJrIqn+OYvVZeS9J
1bSgTnWdJTp67zSsUUSyRepVmLSxL1STAF2oUqvmtU+rse4XsH8FS3LOxB+fD3E36xcdUBoHKyrf
D7WQBYd44msrvnsMs8WGI2SQbClSXaGUHIgP1KMu+FRaUMelZ9N9LI2AYDNsEAykF75K7hl2FWRb
snIzRDPrnumidnCrjgPk7bUSJL7T9ZVm8qw/WUhhcONFHA0JyraC4Hpl97GgPvDGc7aTdLy+T45Z
8KuEUJKELiKTqdzAvgAEi0//93mD7y8tMloj23dDFI8ZI3ZUaY7RLMRhJMZEteCogghHREwd8+dV
rfVFAqCNbajNkMfy6OhviSVUdaX3/vXH9F+rbhgQi/0z86OEwLIRm87nwSAsBjdXAeF+xWNY4l/c
yH0+tlkySvC0Cix+oFhbfEqnMMVTv/QNxHZd7aFHpLHMuI/Bqur+GowaWk9EtvU4kVoojYnW2dtb
7/CHW+k7piXqLbsxmmv0Rrqd6A0hVmPGrL+f7FF3XLO+mq6jup45zIcXUXDkyDt9J9dvoEfmiXz5
w3XlweCD2c5Tq0vP9pzVbFYNYK7saExIfQp8tMrN0DtfiiBRtMIcOFvQc/J+7i5AM/KqTjbCJyKb
JuAoMT1IXcQsTOd2dNHFQLuyznvRqDLPgYvudEX22aQ02/ioqsyZg9LZAFnRY1DM0xuvYrMMGZCZ
q+mb60331SqSj7NszvKw2t/fwJV/E5tNSocUbKiLhNp7owIK7NWnkuIU1HI4CpaiHbI9c9SfqN5z
pRyHVRMYd3bj3pKBZ3CS861HzwQ7o8rJHsDYv8cOjY9/0LBS4wQDzt387Zhbd3lnvpxqNbTXe4LY
iBuYCimNXHd+ZuXDbvDicG0g+WNnKg7kpMKPgjPgLprjR8JgvM3PaHWl8sAxalnNkKKFW2HUjfnK
gw/A2ugDmwWHXNNFyeFUVxGMl2oYTA4GC3VoKeXC6DJZkTBOY7HBFRWzw41amfZU8eDeP/ZRD/JY
VLK5XSfrR2EnB5GwWdcN0gUmocaEzaQkV3/rrBCXo+arCiFTZTFKEHwXVxPemTitNtpRkiR1Y6Kc
7RymkJRMS+gjUjkqWvlNSPEPquGW+39w+tfbWF6TWlMHskfWF4/S/31obZq0Q7aRZ6PWvplxbPwf
5C+3bVYcJhslhz0HHP+RepmXsQmi8b4T7RjFVKBzcM8YhJyw4PvfRC5EbIjfOj76xXKwad4vUr5q
yGYwJycCgwSaeSWFW7NnrWSmWtnmo2c8usYH7zkhcwvgy6aPoTbSu5MkRwTZg5MuUOwyqAY2m62w
b0XGlVlsNsefYKtIcAmHJXtzpunAt+LVB4+eCyHy1WDCVL23fe/hWnfCreuNMT93jDMPLcX8di4G
TAS0KuhdFSvlGzLs+t6RJK9WpUolzrdo8ha6r/L+dUFndRgCZid7tLSk6byC4eB1CksGe6+AI2pb
PQ2yD5ZWYt/XIYEHlafDvZO9a/tZzDOkxLUC2ctGJEsnaaUfPFoZN0t1X5nYSmh9M2G3lzxxB7VI
XXTCw+YZtbeQNh1iW1cbPjEUsd472Dxi2OMmyvIJ8eNZUTNALiGGl8TzRj193e7/EiPKozt8pJxt
6TmyrZ0tDhU+W0i0j/OZnPRs7zR62zhWjcStFGkxGdCibwX8hikx5r/T0E5b2D6ilUB0c1rjaXTW
PcczHDWieZrRvTRisui15Vn1OCcehoslIpUnLoQUbalm8rtmhGS9eGomp+chBGkeTlywZFdyGyux
nkcm9EzSl1WLKj3crTGg76GUjFlRIung2NoLOqZ/bkHU3sfexV930ZDATRvm+4z2L63t0pDLr7KO
Dgbs51hDLBGfNio50gAVPBOmbp1uxPGx4UxwuP8DnqrHC83WgZrUWgv8Fypbn1SOKFdot/lCd8r/
KERnely+FVwtdDa9AytwjwdWfnL3yEG+tkcnkzj0lJ/cwFzB6XBkPEuoNa4XQ1upV6MEg4xteLaF
Xz9h2IgOHmjXX2VYHGcRqiqriIUUuLo/6QEf+kEMvlTzg210Auca+InMqTzKJBf/QgNCM4SZK/eU
1n37jzPtAK5YyJUliXRzE/EvBTmXMEjNwXR8f1xIFgFJqcZQb6rYr3knjnJWdNLc3e1ZyNKjUP8w
PiphSb7drOClrTTCavNLuDqgPllFE1FD7Ystf0a3b4+iLq7YYkDecLcQxHFDd0wQ9A9xOTJWFUmd
LbRKOXJt87iyQd7cFHACzMImyOzYkaOidphdTIz3aAgu1liou4f/TfgtLnzTLSfS+NcjAY/sSfy0
UvwybTS8x3uk5bQIP3BPyCImwd9MAbVmPibo2HqRES350Zt5OLpOTJbyD7gQSPSE08I8CLzZseEH
oX5j+eceGxEY4lIGlQDZEjhufiqK2UsfGLS5Fwo43jWMxbJ7G7PFeYfA/Uu2pcIWRBYUxoCEroCw
vcZ4RP6Ti0E0Ngc8ZPX9r2ZGtuaDkD4PDy788xqnHd8OmrA38JCRUUlyx3eVK1d+ZLvPeLQ1qC4G
tVtMM6hlJ5TEk+06FbM5OVY6TEgNFdeWl00mwhRSRrlLdg95no/n8svnDllLzUhp7f2oEoNRD9PG
OcWzzgzmthjJhpTx6YG61WJ49s9dhCOshLE+L4T3Lir1heGdABxT5uxMxgMcN8IICFTIP+7YP93X
cquzBUq79u5HKiZNPM/XkbgYItCcXThLnwA3W+34OIWgtB9D1zzgb+hj29nehx/zhkd2hC7tUuxT
wDG+KJ6UtwczuMmk13OaIU690ZhDHpsWXnDShZmwH42s2T9XOhs9YFrJ+yMcGa9wYkCg1s4anqmn
9j1FvbZTjHORFdtSZsHlxEa98PLkpg4u62BfdD5ySp88SRe/ZvWihW5yaSloOWhgQp2HcvLJYf0m
cOhXxzozlOvfZhcqIn3BXTZUS3kziSvmul2N+eJcQAyCQIiKRWt1xE5BDmhOcN+LOZKClRi+HyZJ
IdbXoRGA9gpZ5AevEBuFwtoyRC9478S9YC3rvdpj++NTA8db0GEg+hs1XAmrVWOiNjPkt00HwVZC
NrAsm+nVnyNPMbUNKXBdSnaDlOKOLSEF2G5w9vFAIkjT5ieRFLQVjTwui2dZ/5r9duH9fIV51HKj
nhvGgBmTgn2+JNCBxrLm9/0qrgn0MtwlSrsMGAfWwWIg5wahBJnzpoXf5jG7meeQHu7sWbw+aaV0
ep0bSCNMic9PtaC77teb8LthjnYmSZ75ZRrCfazmkfaHjKlo5s+xsEn+AiNKfZaK6UICxpWNAVc0
PGF3t71DMej94PWtm0eugqiOk6RsxrdbKPKKIxyRhvwswhpCHQplAk+aJGefI2wRHP/CVa3FDxkn
+wlcvHUoJXUGogU1GOog2nVmQqgwHY/gL8+EIpTjUQrcQxK3vAYycL7IdbxgDl5O6lSAuwUybaV5
LntBac2sw1egbsq8K9ruGenWrM8xq0EBrQwmEF6OEj+R8Z+DhLAx78T+xDDl46WFLo+a4pwyar/6
eBSf4sXpj1r+3uxpmFuJ28TRH8DqCbo2H2sc6qpqj/fmErPP6XYQHdaEfcrqB98n4tR2WSsmv0K6
bSBjwk0HO7uL2GrmnrHEvgMN4jgjDVHaOuigClRR/w9TJtnveLjctnLtG+s5eIgrLPsSb5e+Z9YQ
vB9s1MQd9bHLu8Fd3mvQmEWB5dD8x/e2Dh4eR7sv2Af21D+z+771+U3/xtEUkulUZf/vl4QBvUJQ
7B8G+rRJsZy6kShw/o/soxei8sSxdrqTqFZkGT8UIeVJxYHQqqPacoOdnUcY7J0xc2USG3ilcNjf
WXmeK7459JG2rowYdNZVInuY/qm90R6zKvv8LQ7dEIBORwr+I8n4PaO0zLfO0isBziWtetdOSKAK
qdxSFz2y3jsQdy1cRMT5yqTU+Fu12yyzd1mC0mLtjUOdJ7G3Yu+zwpd5OKZKgDXnYcGzWPL8CR4Y
UMyFD7Txd+QWV6ZDfXtVje9g49WdfPnaEsVpghSfl48sBHRhTU0T5+NSk1kGmI/H1btXbrnjmFr2
XnghTCo4Fp91+Z4yaFHwWiGBQDaZbwjJPRVgVBbAWdN0Qhw56xiAcUxmzlHO+lrlXuk2Ls3oc1Oo
FKRqJzg3clh1xgLDDwZr3sNxXUXeQSgpCbWIzN5COiQ+q19gWJfPUyQNklO93kxcJk2adEZjYw2T
AEjobDHPIClZ9l4b0ccMXfVYeMtGEwJpuXyJijNY+DpY5Szoa9fZtimDTOIUX5I8ynEYXF0EJq5b
4o7yxx+xZ0blbsIvLHqjhZNwEGCFRwPwE05tFVs5khTQnA0MyydFbUQ6BbWuHQwFYkvbIMYpxUUC
JTQVOJFMN/LXEHtOcmt95o0NO2R/Vr59Y2ZVN27MhFXv7KcSIKlRm1ibj0dy+ctXva0X2V0jLV84
2P/twDGcqor67DDr2xwk0+LuuLqomulZiJ+YedDDfVxKdxd8j7FnKyVr8R0RlgILSpXlnIw0MLRf
pLdwTG4wMu5mO9eC//aeBB2zBAgNx0028IhL62NJQAdFv/VqY3gCgu6/7r3gVNxwW1UV6UHOU+2i
7TtMUn0qqW/aEdckIcMrTrI7UoxslIbUSKNEhaA2qoandxc2vsyHdEPS0vUSwUsz8ll36nUw2/L+
n/xzkEHCIL9z71y8VdJJ0LkooDCx/pK87pnmomHzOxncQ8AUB/o1HCBplL6wf8HNp37FSS+sPiZz
rQA2Bh9pIDftvbaU5uWZ2KvaKyHqWjlFeNI1/WEXbjVxYn0Sy4US3mwavtRAJJq1cFNr9g9bs5MH
q3T7AW1ASpwH4dEbQxqLG+ET/WiMY26s/6R82AuPqVwR6ky6sUz4QAQ+OPFP2Uh9iYrNjdJ/88k2
Rp4FSZwpt/VJido8P3kl/3B+ZTKh+caqu9pVn4zsy6f+lJgJpACRs01WyTK85kZdCB3QUeJ0OMr+
y7SdcZr6HnKEwKbg7A4BHgZH+hbQwLnjDjABBAQEgY8UrGNErJy4f7kl72ngNho78CJgfxgJuyIJ
Bxu+PkAa9gUWfQYuYYbrUQUllBw6XH1RKnJmZ25dMrZ9a3egS5FrrbkijliorgI6YBZYpSiOLlIs
rHtLPCzokmvHhJwvCWGdq/DqROHZokAjzAjIRu1S6xQVB2PY6G6jkiBX+VCins43Fvp7QPZ9f6gW
nabejXawlWVksGCxvz4NF3FjGPzRSmW9NGlqJfO+v/LjGEr2kjUCM49lMWC5PQiEgPxRt5Kkvu09
onbpevwE2N9Raaw7UUdpZqHMXQYiK9aYkX9Gu5tcKJo8QVGu4dMvq6UCF8/wirG677P86jqyL83g
U6RliKnE5UNuZJz87EsePI/SRAaNY9VV6vjsTu+VDCzPtN9Qh8HMdo+NkrZaNXARdRPQ1C+RzbxS
lXbPQnGdgyYPxseJOkJ1NBzi5Vo8SWhpC4wDzp84LaQs84TDuHtwXU/Cl08Gf5rY71NhjaUekMPq
pQMEiSAElLQgMlqMQAnu/yt0acaphSJriKnphy+/zYUfIqfKeg5FRBLfcbXO2HTX24yrrBFDBPW+
fp2II8u/CB6lGWMXUnLJR+Z1PLnLQYUkYAXjvOrpIasY0nP9Doaz5aHwA4lewjzbHUl7Nb61HSWI
DV/FLKJv07bIWMZyFgzi7hF3Z+kIHizZ2l4+DUe2fD7F8yJ5MXGaNUFIlCPatT1FT+ABg3xMrMv5
wyCpH6vbFMabpQpjFo1t7m7fzozvoXaRtiYOn1jXnF88mbxaThF5ZqTpOfgJj435xLmN06VsluoH
zda6cpOi+K41oUwvaWkcF4Prg7gebOh7aTN5kC7/iLsT8yB2jB2S74NBsjdzjrFhisEQDfJGn5mu
Wwvq3zHC2YhJGQeFbXodqWLQVJSOrJ71TARNoHr4TQ+8oDzJcK+/nDwB0VS9a7cj5RVVCLdP7nL6
YzGFuW1xf5P7XfBQw8HqtVpTZo68OIQTYoAibeGcj8OO1u2/dmH+AeO3UVYPbGdxq10BKGer16OU
sWkAof1FBNenf1uAB5bfUCYFEYACAUsv8CgCMniTTFATZJ3ZzmI2/tKaHzlrAA9ZPl2Zpt/dlI1c
ypYZw3c4YnWuVBdh9nNGSlgGDwLrfzDwGH4qckJdpbKg/xnS24L3ymyc0gqdanrLrdffl2hkVlXK
Q8j1MEsKpECu31S6B5aep1hdcrnJTklYmtTOfjKlccUdDsVkgpHlzR0Ky4DvdEgCTEXsPwbUnx28
ycBW47dz11xrNylU3BuJ2hqTrE1xXq9PRxwhYENYylfCcnl/qJuIdxSWUO6pOp3ibttUsORdRgYA
rtMQvo1NhKBZ4rxJNO//zdsDoe5/Q8v/+nI1o/LXdjBwNvitiIq48jbNefw/fA38IoAIvyt5pslq
G1g+wE+peLEZz7fOip6lcf0nEY9NuS9pbGaOmP+ymodB/DxjVLY1Wn6VbEaHoOYxLuPFr2oamiOc
bgLWey9CAMSkaDkMpC+uDeEJZAJjd7Npndrw0x0Hty1icr40cWIl52Mq9dhcKtv5hqCcfL3gUzZU
nomMvbGi1Ze3D0wXv0Pils8BtBg329zjW90F+tH+/A+uE4c58EWyMxXoaU0xkc1hwO6ApWw6TH6w
PgjcUQFSLPcroCrekm+VTlqMZUXO9/SMpU0w8wylHY7e57IZSPVh2FcFFOJW2ubfBgNCYafhiE+D
NIZHjm/6xdja8Th+vauBz3LNMxrDYpjZyVfpPxzN6mDfkc5G46IiMNira4iO16CJC9v4lE2HUd/q
wBCCUuwKbIcM5imMjxBbfiyxjFuU4s+KxbBjL1NhmMbKJNDx1/9j+Vz/9AtOte0p1n3jDtElfLwH
Ap42jreRU7Ny036WJXuos362TgYfT3OAIPkO38tV9fWqeJn8Of6LFzXmJx5OdvYi9kn82VAMgKmP
/6g6otHVAH9vT3T8O9I1mqunw63ytfVjZ5htCcmOAWbmqYokuExFxbPi/gLgoCpPq+/4li5kbyoU
+LcIxTmOCxPaCdFLpzY6+xtsaONUKbqBYXSUpvWIEgoDztm8K+JJTC4bBvGhzyMYT+KKbK5rhAC3
JptthS1dzWYqnF7V7ABiRHEYSs1l0MGDHL70VlGJa8VW3jH3bOmpYr5PfVrZQCaiaCEu+xBiGgum
Vhnj6ka/5wyLWQkJbSuLjOYEvhK1U2haGKI0njQTV1ozWHS2/O/0bIJH2ECdpbJZ14vNNde1w+hm
6mkwbsIJy/Gd8O2al/D43qryb153NZQ2ZgpCbZwJCb19CubZO9rfVvPpO0Mb+e74Br+WLTIB6r08
VUS2tJdyWeM+oXCLPfUBRwyITRCxYkBQwDYc22+h97hMymLzUXbXbnfg1sOjU+zo5Rhmghrf+A4C
AobGLbiBTuCDyvNMO3Jw9cuucZQPi88rMaaMneSVff5KAb7pMfR5RFpu75Y0Tz0yqgsStYFhVKO0
kUVWodH/miki4E865Dxs5XJXUF7aWabUTGMOE+9L2shugteVGeg8Spoy/iKEBmA6Pgvv17+8/EZ2
uhk1wTgxfD/a9j52rOgZ33LpO16BWedLWz6Z4y8nz7bb68FeDIrKxinOg/HDPmZy5xSlsd+wmHfv
nj3ZQI1vFXlPwF3Z2PY50AcgbvdMEBiWShkjqd7ud6t6M9PtyScbWqudcv0qF4BH3fkVoeGDVXLa
97ORyPhIkrGv1bcngLX8ncJM3DvmOBRWaIeFR3csfSkMAxK1TgiTjtBL59selyvyg7rUZ/XAH5C9
mbq1mGz8qpYzgOIm4GbHenz18kcf2An8/sYGMG32eyoItJYdv3M23sK+hD/KGhqr2VQfr1KPeYGh
/aywkXxQdDzosJYanH+TnAZNozI8nG9SSchac7qezbStrqH9w7u/WHS8jVObDPfymMRFIKxn9iiz
tFOwRBmrsSSJkWNSJAv2MWB1kUxI+BTfeKpPBB7hZu095AIc02k5VtYSziBb/LfI8ZgHrvhpEGdT
k3lQNzwzz0QSJ3Tg1advtuiS8sZm570NTAKPLFwjdHHVpJQNDcd48NjGz7SB3bXS8xgm9Viu6MRY
j1yadIluJfjKJucSNNQMb/EJmfGb5+YZSaahKZx2kKPyx5JTkK/ud/EEeZMdSJaJ0idR1q+zPCx/
YUBvszN5ffL7/DXtX9KxyekJYGwbrzpl1L2d9I1RKM8CtAX0k0YRJ6wOpkrVKfhPGiUgg4IoM0Dy
5Rw+3X5b5cbjq7Rqp3jNOXR9XZ1GiV04KFX1OYSSitSlzeG7Ds+/AQjJFwcv08fHiyloepI1KD09
QC4lu2fOP1FxMW6BijL1Rh7vLNgpnGu4xmWA3/mZeoADEfSn8zJQriF121oaUWjSJW4mzGTXz2Xd
JxJ6sC0Bic83Cn+GIqNDSvtMiIfL/bNhY15kaiL1doXd1fiDXjob0c9cjqhJY446vfietbXisBl8
6dnHOzeiRgZOpHPxtHgiJl/BsG2BfLwkoGgpLPDR9GKtooQ6UnvfjWD6aNU0fIyK9a3Xm8JZlsqJ
uHb7jdByoKAjBkg+RMzoRxYOyiym6lf5RfNsIc1RympVhY7c7O3cemw9K7Gbek6rOJVy5a1Jtg4g
Jxq4iIB7bOybKG98S/Pbk1vqeyrEpZ+WOh1pT3qJrHMFjsjAl/euk9vvoBRXg8HoKutgl3NexTkM
T6jsX7lhTW80W/YVzJwmztc8uRVbF7zelLn6ZgseCdi1/NUQhogMD6TlENALY2nkYKleFGVE/QEu
IK1/w15HVpNErEibIrDWd+wgMsGjwheftW6xDezDAxURk6UpX+RZroGtOheSkOCWvDhPesoJL5V9
Q5iSQZflWiddHWpRI9v3EClHDUnLoI59nk7ga/5+kKkVJ9mLKg2lQdxm+jPXR19DREafOCGFQG7y
vNUtEW8DPoT7ORK7lr6qshKx7yuEFzcwtHNh46QPz8BM4qi+G7wkmCZ9AMjz4kj19pfO0S+vdsyE
qII251Sgmoao1kTxlTJSTKo+JLsOjWlocVGnSPURPLzNHIwX8ccYnqWUnHrFbBx3G05uIHP/mmgy
RC6roPYUFYporlHzKLHT2/qZrGjrrIf9dXDwL2t8NbSJ87+WEUbWAyyiG7NVbbQXr2qDBobmNFhQ
WKU4aMD3JR+l7+iP59G5PdQ8Ge4L8KZgjvnf9BKjwbzqgZTgZ8hzaFVrtQpNPeyKnQSqkbqwcv9q
yEAWD7nLi9TOB/Yeqw34y6d8yRbX/XynqX6obSURa47kg0LcUWfhZ0obQJ00TD1JL1MyvVYyi1ct
e6F6zUUv/Q9SFaqxdqjvmw695YvOQ+mROtTeGLzwn06jk7TX+5hL3fVKYrbx/g65McRRO0XWcNUI
X08fqfLhVOfWR4w7SVuW+Qyx73smh+pgGsxxMV/aWOMXKPG/L7Z+aUSywzJUptoncB8+9pjugEVw
qnW5dJ81vBmcEn+opW2tGFwOSC2LEOeKUyMBdYTWtr7ISkz3xXbVu6bKtcGI6a/u78Zn5hug/W0j
Q6ql3ulnddOREXgScChRY29ujRZNVHu94R+lbBP24iJMiYYGAd7lBWZBGxg+AQeXVMlCXXPBSAO+
UtySstUqm0Gx4UFukCKKg1Vg741gxGlTeOOWzuaBz6/pffqYU3wErpJ8hb00CkIkKN51gRfbjvHZ
X/eg9gem7lGDqIuoz5qEP47ixSce5zClW1x04H7TvdMcs6ftsLgjvoDOwxMDy3GW1tF4WQA4DRBk
YaJwtmm7MJrcrJy0fwvWjzVzH2KKycZJbIaGi8+t97SDcKM3snTwvo+oTwIkkXC4Kgw4fAK6h/GX
F97w1conTLR6yHqNKwqr3ztmEyyfOlaz9hdNeFye1cyHd6OED3gP+vQhWJkiehhQlnbvdEBExz16
60B72BLqYPkZfUrLcW1ETRhUG3oZqvMZpHuHKlGf212N+5SoOD3wJhfws3fJq6dco0odm0TLdJ3c
5xC25lZkXGu03hxfXCN2gE6PF3oZVDqnqaCy2+paOWrhPY6g1bO9AV9/q1iWN3Tr+kmo1w6FjufK
dURFNd1pvJNv52CU25Pu/jpnBs6jyVzq8gevPqmc+IyI5Wmqr9NwGvZbfcj8GNAQJcaO7kR16iNE
hEaPxH6hzVJ9noEYkbKH51ET1ELsnzeysIoOVJbHej9NVbp4Qiqxz9qDcIrXCp8WdSz0XC4fv/un
BUH2uT++P8++XHMKPoQHMqRy+Uvuytj2adt267Ie+flu74cn+GBCc1YQqEAdh9Qpgx0k1uG8z6Hf
vZ5zNFTBl2fiNKjBV5KnP/xiAecaXex+nL8wtW8alVzhqI+G6X4DhU/paBHomKOgd0FDTFlEpvBp
YEHo2U4dCMAq0IQh0YOzSSHAEMIkiER+2krb875d4Dx4oJ6UxZuk3k4P5q3OdC9WAOKG4jsDaCUn
sI2d74//QjcQFAzq2KXCcDqV928BLfszk5RAgHAv0GwVUCWg+t4+qp//5fkLoMFMpJBWEYhCjE7e
v72JBaoIfELqR119lh9pGNXG+HyU36WraT00RvMU11ZGsmJGDuYHiApTZ5Hn1+vWNh7SGyopWRRi
3eh3isQZ0135IyyT63LxHj5Ftl3lWMK+ZOUFTVV6rb9IZPi1TgXjX00Q1+1pdPhqPDxVWz2F4acw
raCJtKLkI5e6JdqSGECsJu5aYtAtcwrc1ViqS6D6SMTrh3RjpGODWvC5NYZnMfzhtEYcBuQw9Y1H
toz2+F3VSV5WNu/wDcSMqh7j8kabNDP4kmo2IEEUXvJasGE65YvRTpYyr49PbYKuT+6fHYnWbQh4
buuTsdWC3ZqQx1RFIyShy8DHjR5Ngz9Qy2Rw1ccEs5yfbHdMOq63NOKQ2ZvrR11oAhM4fcRfxQwS
LxJ1mG7xH2Q76vkMUkEYOYwCLvg6Nfrrpr5Ys1iEGF0R+/ByWbJ9kOAVZMDkgk+p4glL5e0q75LA
eUS9m7c1iFRZVVtk5mX9T1isxk01ihlqJaXVO5ZvSbyQpmTu4W3CQ3JxZIOyoyGxoTg6PyMkemqP
c71vZhFJWrDxLY7UfX6V67uJanjMnvFZBTuwJm9HudmJ058jwCWuXWhOO33cY4vSOOqLrgn1jt2h
IjrXyE0jOl93OGu52D4KKSyZ50zmeH6xUs68jKoVtwJGQjg+20ewBN9qwIS8siQx3BIWD7wLmxIy
rCvKdEj5kmpz2jsfFYIdZcUdvT+49uWjUvfbTW5pyY29eXVg9+6hVwySJu5xbYgaiywbu32QYwZ3
ZEFxXVRvw4s83H+ASfOvar2p7yYVQiwFbFMwLVNuxBGjAzVufXJckzs9s2Ors/aBas6RtUbVVnPL
LqU1SiD9i3FBnxSW2/u+W85GAY7VVS3vTZ0g+AIoHzXOvE3nhWjGab94VNqX5X3KtnioyPR0BM8m
IGtre/+KqINFonE8Yq9J8b2/uivy7X6iJi02utXWWNqU03/bdWiazlVNGtm+ElUGW/hY4vyekImd
8XOrlNuicDKphW8dcswCu+adzFOZfuZbc+WlfhKFGqj5OiYzo4TdB86DfIgwkKupHNuTX+R1Qs8v
25RnW5vnEy7ZCVx/deLHmU1HPoDfvofyM9rGlutUBU5GNoj3bLwT+HDEjBePib9kU8OIYQKN+m4Y
BrRNUYrsO330+qUETESGsT2f4jtzMQJnO9xBQTQ/xEYMPTtQ2gqOlKBvArCV1I/JNUxQPK16S9qI
vdBImmMKuWzU5hNjwFozbJKqD5CfxuR9LmBOryqQWckC4MvD2nHUTMqdv9KD/UXKzN1bAdxNPedd
PVtXjmnhArG5WijkvCuRHts05tmF3/gc5Yj5Zdbneoi98pt3vtO0Hcwh5P7skBuUG7OdOFGQ+eui
LVJzBdibfcQp7p2xdxWvqLfkvbTCqfDtNQ/5905fadXAftmu5ejd4UdNxMP/eb/bcc5MKtzAIoKj
lK44VI7dSBkpIGe+o0R2tGoIGJ2GI/ch0BCfrmofcui+U1YEEHdLGbAznQ3AIAPWf6M373Hx0pcm
cFEYFam0ZKttlRRtPVUL77MVCK+2GJ98x+PgJlLgQP88LSz1I+/HFArPmX9vmNisuZqrxuxwBASs
eG+s9mFVVgZXG7WuSLDi7buwxRecdRPVHpA9+7+T5c3OhdWp7VLl/0LImb0M+pNNIbrMpoJKHXM1
eivss5/nblTiFffJCQ11p/UU3L9jxvC/57fb7jfjcvlMJeCfWx6oSP+JizrvqMCBKU67IcZqTq3y
9O/l01U9aqyRJyPYVILdXOTF2eV1bturDz6yCtHyN/4LFdrbpbtsSKLA+A/Lo2upWIlCN3uXtqat
9tehfKRSOQckXCLObL/uj4RmWvdFOBlChp9oO4BNs53E+5AVDao6Z0KmUIEaW2IT5vtppTIbeaht
OrdJyM2oxktc/i9Pae3bXB0UpCwCSHwU+puB8cvxvZVzH5F5+wTnuThqErVUX2bulxSmVtYIyT+d
sW7NgsJF9+CtfJ/L26QRJHKE6EZOoCZidzfnxkYyPT0Xg6/RTdKfU4LigED4TmkkGgy1TkIRGNof
a71IyTm1lNKa4sj8MU/A1DElNNmIFqxPI2NEqaj3RyrElEESD0hg3Ldc8aHo1EfZ6Wl9sbbOqDdP
+iMuUYX+PIlO4DKaMS2AHW22nHk9wGZAEO1CUWtI8UkrE/wN+LJHDBcTnzY+Ke1q47yF7abq633c
IfA/l0ZMzWP7o8kzFqymWeunslfXET642/F0D59Rx8NsrN+4EZnlyMNlbLvubQiQNBXICkLbN4QG
rPlmfW21ecqj4FVP2HPBai//rFsztxzxHfdUGW2bi5x+XSq9SLxLlaq7OM5ZjEf9LWwU6nOJs+Gg
z7LE3JeZn4ARXm8+yazt6Og2nebub6JWGxKfysASKpmtACRM/KG9kwEGQOScNY6HxLXi/lnBBBAL
w8CuFt/J2NN1guafwfW/UIzOXEPgq7sGnCSsBWhN7twU0IB+XFmdNIw2ffAzQYIOTHfvEXr1/8U8
Yo+xjff0Wn/XiXUz3oIee5mV1N76xfj0NXVvpwIT7oTm7xJ0mSo8CVXxTjOwiDt1SeYnMGC+diZE
XTE0U+guwnOq54lh1IVrO8jXpOvkVq/S2ZyIQEP8HMzCO1NuNm+akL/zWqhDm6n684iC414CEHcH
m/IP/pr2KXJdWvVeEN4f/N26tvsiMYYLNR+ZOF6N3EdEmtb1ScggygYSO81ow88KDn8wcogC3bOv
deQLrYZjOl4AoTxhvBYf0/T/AxWNhZoggRIXC5kzQdqgU4X/AFwO5JeQf8YLdpOhCXRyHHPuwxwH
HAjNfFlziieKpEp2gK8MTgsM8W1/X0HGwoHDAlsuhnP77dCKkNcLTkHlyLADpY+jiNi4ET38kqqA
63W93/0vKtQY1ZK6GvhnFBtrjjamIzzxM19Wad+b9a3IhfI7iPkhS+gjsnW/wbab1uzjowp+AXA3
KPUKcUzQwuZfSMRBvc93CGl5qwzb2paGV4xo8Le8GplvG5Q0W7R2z6T2Bvwrkcv/ADhZi7tZcQXR
sBAu8+b43Y17QXbqj54TqRjiP3gRq0bOBEYyN4xMimBrEJ7wii2M2gOzwXNn5JNoGYaBo8F2/woH
1A6oA8NZ9O/5lOSP406xrUds+X+M9TU3S5/3Kx5gSDqvYN2Bwxi5JDx6Wur1l54iTToFxSZkEzMk
Anw/dvbmgMFRjCuUT6PErd4vRkfm7hqI947BRaRODoSnVSnbyFyTCePOF2yRHKBDlebjr78HwAvq
5gBrtrFn/OCpg0gRk2qZy+CUtj8YNY1S89xncJGtQKeuCDUtVAgP7pTEJy3DH+dBykitgryXYkri
4B3UnIgBcVPtZhAeApFgDfJSwV/avz3d7GsX+n93KkQX4l6Mip7cFCs6mE+LNcQFID5mLDD8/UyS
08XWm7nioo1lA41q0DjJJ5MEyZ9l/XPT1x+kR6KPo4NGIwpCVp04q/S14/SNpvyX4DJrGmvBrtG+
emUMl1bGPPoBkYkmGP1seDYNJJes5/tgHQurLzWHB6d44iEMGb/E3jqie4BFt/q/nC9eH9NeqFki
XgQZ9j03HWiily1WVeu0mk8WdLFBl30c1IgdyXJlmisiRzxQT5nNZes+wCnX3GeyldtcYPtPH+v6
O0C5xxwmlJaaKNTFbKpAt8WR0DVkKT7N5Ze4ByQIkWkm7OA5W9lF37b9D7v02RwaXitF2j+XvQwV
l+g3LQ/je5lQxKzuaKi12OKEaHCAFG6KQNHwczLKwt8Hs6huDBuMPiXs3jDatSu1hf5bY9WNFRoZ
HQj2evzdNm4gRRKpeEyDeTMy2jgcgh2uJpql8MwzwmS882sXwR91kK9DvUrpRKRTLRzuuVl5A364
QyA7mQhz0H76gWXcTTRekzb06rzpRKW0g2I5lEMh6zcoALJ5AU6TUFKRvZNg5SyN6Mrw4D0FyhHT
AwWNP8pJZ40gijU9RBwkCSK+0KImuhjRNoOzIDTvXls+oy8Wyuhr1HYxBGTeEcLQjMUBB4cRxFVc
WRsB2zEOHgqZvdMnqoBb0uVIN+elEAkXdnMsbRIw/6jZpJ3b4IVMUoAAXdMnIqS8anVX/H66+Hzx
lToq4ndCM+SvULVAICRmqsIMXjQZn5ZYI7n1gBSV02NIaNBugwH9uqZTWXULbRMl3wDTzqiLJBf2
OedeWTt0DuCoqaUyt6+74hi1yhk4QGg6SdUN5rrAJHmtaBF89hFQlocoj+hPYD6b7RDywgLf624U
RxjQv017177r12GVS5n9oCV7yTwXWRODQ313zxxZRUarlSrkEZ88W1fNvBS4fJ8odePwPNEZDnkF
NTGGZmX/wdG6NWrZO10q5tBZinftKGoGZSspIwVcMb8yql+Kfms/9r/iGPxH8nVr1qd91x8TfDyb
+Z6ZG5THY2D1snVYVdjKutuN1YcM24aIxnMg2js48ABQ6fPDIem40Cqj5/0wNrlCInvbGmd5skUB
gvqQ59v1ihQ/NKGTKhmo3xFD6g9lcDb9m/wz+OkYqN0EKdiRUb45kv+CUWH/BtNFDi0eQKQe83/D
VDYiLX7b7XIDU6VD7+Zvfep5SDmsR+6Qpt6h0apCX1bD8gZU5oU30Mzk+WTG1rKXb9khvPCiU0Mt
n6icpReFG7QfN8Sw1frWK5lE7cC6wncaGjtwq5XRdwjD2tGOdEEg8PmEjSVZQtyQr76hLAj+DVuv
qCaTD3mJqSXvmi2OtxWFQ+AbaMrDHuDiwBRU62VcX9Sae3AggNUW1KGm7NKshwrBL1xi4A3P4qfm
8n5Gu2MwSep09f9tTH2o756Fasq9U5kQWVMA8JqqukorZDX0ys6RBY0E7lVUgxF2cF6Pe/6yl5K0
d0PxrrF/KUKQASnssLHZmfJa7+aIlsPupvdgHXLrpBm9t4jkypA/XU/5/vh29mlGKXXvsXvZo192
Xmq400zyu6bLTM1RXpWBhU2L3n6DtBQcyBhV6yJr4wp/zBJTyJEOA4DwAVXOosCAHUSDpUHHMDsf
22eqVN9DLnBba1yYsjlmWaKYkiO02i5FEy3qbuPzuvvEoU6Uv41sMN71Bw+jzOKXogqVL5D1iBRh
LVyJnAwpgy3B1xZqtOsDE0aNPS6YeGdWa17f5Q2ybhO8fn0NrRqLFUasVrAtkGTu9+iEWctRKSFq
VpIHBvu2c+1Viokdc2012MTtQhitXqzXMUDs4GiP+f8EnQQ0ky2m3zoMcxTBNitP/QNLEaAFr0mS
aTdVVwu/MxoqykBUvsu4jpWdZ7tXgdWNRJ5Y6xTCZS2bBIZb0DQCfEj/aEOZAlrKWWDd4t5GfAxO
UbK8eUBiBtX1+3cP6kfK9BFiTYLYprFjTlvfm30/KlNm038nb69tY8J/NlwLgQfw/PDk4GZTR/9H
46hlV9ubKVccrQGIJA++5KADlE7dlAoW0yEoFed7hkj1mdfmzAc0GmYQAM3U4WxXIid/5oCh6hhX
nVGwupdhOyYtGyM8n3tSshonRQkfHsh9gue0b1cU0jQfmv8A/aTtYFgnQqzih8hwnVaRAefLxSfV
ve4txci0incB2uKadZ0a2w12dwyjjLIUWg/wEIKcf4Mb0O8p4Vi+v4kMFTkiAhTwoOr8Qovo3BAj
N+SY9icVRPJ7pB9XeGSZyh5dRutvyjR7NrwvCRDtajKXZL8gdySfl7hZBAU6EGBnLfkpsRXmLT7M
Ny661qVqj4Z/a52iUZLEIlrws37g1jj1YxHsliHxahMyMcdIkkMVSo5rUi/YxSPnyPMumhTsxvbh
HqFTK71bledxX4GXIlNoxRvgNYzn3gbwBwQFU/SNoPXbswVeaN9IBRGV5UuhIFmHmZMr1ayCghQI
/ynTBYdBNcKedPOSczmhdHplw/VBd2xUNOy8G0DCQATGnLrw3QHlUDbDBqs/wOb8H5Pb/cJ1j2jq
FcnbZ+/4BaqnHoiJKVsbzcCjRQv6xZqJe85WoMa4/aJ8c9teQjRvJpJIQhm6qrPJ8Cjv/NrJOnJ0
+EKa+lQvSe6xMlnBz+vDUBv7lSAVciQbVkIrRmUAIAgVF4awqaq92JN1qSc/dw4wCnx8aSEqpORc
YJygAtfopEiLyx8hskIyOXQx2cTj9Yr95HlyN3G1dBgDJ8QsIAtHZjwziCspn9ilEPl9uxQVT0a0
3BrgaLIfU78/Pf8or5JpbIcuy/RhJk0adRsEjRc70ITWu6HPPlnf819tzTl5H+Mk1iZQboQBdrHK
zSbi+ezeiUmW2BCFQr5BwO6y6WETV3+6FivevjAW/Zlj96jC5FwE7h5gZdEupH/oau3ceSJ3LGm1
yJi/rkrnPOA3dZ6eoHbH+UVrZVAFW1wBpyqaZCCeh17vkLbrXFZcGt1wATsh6xFXA3aenk0VWZuG
aYHOZA8DGakqK7xIvngyu6kzMccgAfVda27BAmKE+f2hT6NlZv0jiGjYY/crBEaLcYuHJm/cpfQr
m72v/kDNsFiwC0k1jHgePOMjscW82JK31KHG9MEy5Oqkio3klciZNJzadCawRdeoj8qwd7rybMRZ
s1C5/UPkiuTVBhQDt9jUV5hgC41Z2QeIkaFY6GeKZnSObrszKFdQ/Us2DRVbVba7aKZ/ObSdZWs1
lN/iNQ7TfCYnhhLoOUiZucE9O8jStbXe7NtQen5qYEqi51g3Fql2ZYjkJu9B03yTUugapqadfYqe
+xC0GhOdJLJQqEj3Kz1LYauyXqvFsp/fw8irZCpx8kbqjVDNkREHlG87K8CBE+DPG2yYetmQjtX9
oVyA1+3TJoGcDkO4kUiJxXq6HgauaGg3QpiDEZueINi4nRk12BPJIUpKfJ4kAWkubAbkjkFugFzX
zpXK4zgMKKAcTTTtoqSGJJSpzjWyrygAu6crav4jN52JCLhGs/WvoqwwW0BApMpo5qN8Ru/5wzvk
m7K/IpHnrkdp14Ey+Sa9N7WTNAJ9nE8/zmQcjqWQUnuT6XZUcOnl3n0UVWx7kmD+vWZpQhaF4DXm
woko0DXHpNoUwfm3uadHOJIMJ3W7+eXobvaGTEduA84t+TbDweT9WrzBqpTglEPrQq+JHNPcPOgg
DtUCaxBbDvBqzfTslnUjPmlEU1Lr63fx2dI9XbF5gPKGf05O8D1PSLLT9qHLYVjtjqyRJdKCf6cG
RLEvC0y6T+9W6sBmAddhbK9UwbCP52KeCPozuciFEzVQ5JXJ9I1sItrJfA6ikWXK6Bqj/lMew6/0
ZPhi67jl9bOa+QyKSV6AIB8mXQlz6cT5WFNlxVVjPx8idaaXrTkR7zfEvd0l/EofqquRrp1C5ss2
4zIW10uQhD65ja47Jr0o0yB8acQtBgR3st1GH1FmZ6Inyx1C1sAlu+hc3sSEMczw/lX78jJ3qbSq
s8kNNBgf+q3ms6xl9/+rubM1kSoyaVW7btp6hEQGAw+0ClbA61JPpkOtNRn5uznZWQaXdVbF4rhP
hHBMt20z/mVxRjBNlQAw2z5yDyPBLf3s1wz6JOWrQiIixUbipyawYRvg7Mn1f0g0sQZIUG+/bs3B
2SnLw6oroelJxUt7VcWpU4ri0Mw5hgbrJlHoFktzFiO6blHIg3KJ1Z386bcLdcu2oQH+tlL7erCs
tTb6fAC7qBJnHr/ztbhFg9A92ptib0iFuEO9p+hSUJLWDaxZmheW46nqLak2C54KOGXKmot9kkQy
WqL3WtOHsC9bsKDz2QXocdTYvxlxyAepQeXFlxWZkvniyflrN5BQYPcko4RmN81mXKzxLZxFLNTV
5X2gs/tX4ssMGTETtivnLDQFEAaVAIP8vMXRrL9ePC0xJbNaWM+X9SL5cjaMR/PEjzaaGksHePJd
bCq+FafKq/HtVlwKon+v9Kscv6u6FFYBV8EpDE86ugoXex5tqp2JxOYYeifkJ6vzvgkcI82zaWdo
bda8c1+owHZ061JYHBLwUbaTkhGTYeCadu7sz6BlFI7PyyJXwxqW2ki7A0SwbSrscnXZluh+oORU
k872JCf04rJWryFumiCksfxsBzjt9Y2Qxj2WV2Zbnb3NFppCmHPRFGfrHIvTIdEBNhdUbNOIvSSQ
DWo3hbJJer+HUNYQOmgANrH9LhVoWpBSBIxMDSoPK9GG3Jrm48FWURiorE+0eYwJr62IcISMTLjt
gR832JNyR0rzHaX6zdURvlfzinzd/mid1ArIkSnbC4Y5/wNHxfkdy6LrKB7VYsGp4x/ZT2+fW1e4
lWnz7Rtqh6zSVDgUc1wFbVn13muGQJMW4W/kD5ANHGlZatTDcWHprj/Y+7BLJBoqZsIJ9V7wX8ZG
cKgw4bXJdNSANus7TYmQYfz4MtXVbD3jPWTaCM5/EHyrgZy6DHpkHPHS+p/j+C5iNHVHrw/90sal
CdWLJK3vb+lz0QVf5hjdNYmHGKRod5/XaJ9t5j5QqTj0bJOFjrQT096VbyOfVrMsK0byU3otbnsF
NNlxDb8PkHOUxKnYX7KuR8Hkt9ZhEZPfbsYf0/J1FilpyGdOqQylnp+UqRt8mukqUrvADiUySDjI
/Wf2rYRmGN427j3Mutzu08CjvWAIxjvpUDDDoM5N2ch2aP1UbUgjrvFQ0ZowQ56LbKDvriKUmHVV
wDUzC8amsokT0lO+zafLybQiQuzZ2iDqiVsozZBUvPM7I1Lv/s0cPfkmlN80MXv0V7uFN51zjRHX
XY8Gpk84/D8wZiGuogWX/DtSj7A23SEAFYg1EnqxjBcYTiU/98Hw0Szaim2wHydik70c0PoIP/Li
cc15LsSil9vADnYU709QNEZaMC0X3qcOzNeDn64V3HGP/At/8/rYfj2P+AjJ+jRHcC7ZDTTwEmVV
mq/S/Yf+HTP2D1sQZgEpqBgIvweb3DQT1eg0HfJgwVg8n1wNG5EmRxTWpd/DQQlxLfuOOILnvU3M
ZIys6sW5Ya7Ms+Qwntizix7d+CHfk6RzhWYbsudiqbvgYwsCtXs1akc3omZ+Aj41j3Z1KmDNrjUQ
tKkZjD4Wsc/vslJahQUKpzdUTDawa9k/gUsGrP8outscyQzROg8Ne9vSpAijOzZVAa2BmDVBpRYn
tTj7ZMN4K3lfFr4NdBw62lqlxlN61H99qtgT/psQriVZXtHyyKBhosRvEyZ4o5BRX0orh6tUdvQy
EJjLA3/LS4cZMPhMd62oPIZQFN1Juqwnsv/K9qLJkcknd+f26iKlduT5a//hjv9WxRGwoPbp/ECX
qIay+2OoNAkXYkek0xXekNMni6VglMHSGwLbRyI5Dw40sfaQV1FNiWrkAFTPBAhiGVsw5lmib5i/
cTlQGcijrpkm0pWSupVmRflHLM0rF4q3L5rU4hqxHiyxHI3Pq6Po0/DCDCIRr11rm+rK3oGAfBYt
Fu7wDB1PhGMQuXJW/XdNS6GLio8BdJU2d0e0P1fC/g8skE12V9Tx+u7+DcI6EvhGEqrjkGMdGe0o
ZFkZ7eRQpDHutV/EI45ERvRZE0OpgPLrBcTIiwyazFzcLQ61i6m/4A0kR8htZLaDa0stnh0Bjzh5
yg/x++ojXaNgoGf8+TKJ4f+4csTVj0n7BbZR2f0eV0cK3Fe3l6iLuoZLx/k4tCXVNEL7gDn35YVA
l7xEAvk5B0i3jMD2s5QLDsYQ5YuQZlq9THte0cvF0Xxr626sWX4wXwXtg9nXFleGax+3FD7tq8zp
Uh2Nb/FWSS2FvKXyvZthP3JPNqUmb6a8jG1irJ1ijjfkw8DRuX1Zbm/fmkjDqTFHdJIERdqsQ+It
ogG8IR3nnX8eOIkNTa/tlmk+j8YJu5Eu1jjT9oBmKnAnpaSUAeNLgWhj9Q8h9x8rByeRDfWrvdQb
hUx6vk/1EnOCyBMLMffy0s6/jxUE90Kyvt8Ov2xoy1lMdZGvoFBErtlOZgcgvq4SHWtsInzNfRwL
hIJIWJRuVy6fXe5KfdaDdMb3h3jHZFvJ37044TbbrA+G00Eft6figFVjfLciMGXj9/aMNhODFjeC
Esk2Vx5qpeD+AN5Cj/6wq1S37cgP2M3EmBfH8iuscBDH+jcVyzFDnp7CI4E92z5e/hq459lrnn+p
RW7BrEsVKSMtc+c/lE6u89lJjQ6h9JOSfkRfPYLo53rnK217TtuH2QIwfpN3of4C3sRrPiuFLHkV
hCmHRz1kQ7C6LrDmej3/BPoEHaNq36//vCpXTOcWnVUCKxC6XcwoW1arkoUzz9Y2JhQhzdQPp5GA
Msh4kw3+mfhiWt06DK144NbMwqJaiQtonzOtds+8mk0rVFVPYNeKLbTL0B340lXJ8ovKl9TVISpK
0T/KefGrdiip/utXL+bfHbVqZDGfp4PXjhTu1++h7Ry6a2qyYF4sdi2z2Mq5LqqI85iC5ZUE9iZl
qN/dM+rb96Q/Uwihk4EEV4ADr/7yBfLsT4hbZ0gZleE4v2I1AjuQ8u3GbieF+gC5EVEV48FSxC4W
8brffzyM3PrbipshjMMvsKx7dxqCqyQJjcGqTbzRt2Iyatv1cfnwbSuHBZo2z9E5nYyTttNkNiAB
oE2k5k/iq7nV+L8MfnKVaYYx25r2ft8TAG7UHOCo/vfc4GLFsAMeS7wXUXAzHpHKQFWEG15MygCM
WUBxg7uWLTh8HbWVVm0SlDOwVDoRnoRy7+Zitf7ASnzwaZVUkpCPeKl7H1F5/ONcYRhJ6TlGjV6/
NTm4zfJOkKYV6vjJxx1Sz5tGNCfw7Olu9LXvjH33IyGJL9rfWRILuRLBwMiMBHjsDymBnJVOgyZh
QISjGtCBFrdDr9CLDCrXsgaUK789j66RJKF38q9LGB7svbF2Tx2acwnZ03luVG2ExlcBZvVGQLFs
rWJWvpAZkxKUb3f4aD6e3W1gM1zGjBvHBU2Ru2lsJx11KnDs3bYef1mg4/ySK8BIV5rWBO6X0DYf
LWtgyXHtI7BHqfyYWf1VPC60zkTGmcgG2An3l3flYMSJ1ObdjE6eaM50wa1kr+h69pDYfA5EGqG4
sc6vifhcg0dG+8gfdNEUItik/UtOLxYR13x5RV8De7nu7wEOCOgDVLtIhxdrZWQHB+aaEtpeNFUT
OcA1NzBFLMgbvv4jiIelak/YNU3s9aUZcsnRTDtfZYjUxDeh2Tx1mnZqEDgYKBXZpAEoLLpwunbk
9428WVv79GX7SqLAAes+bZHDFguMAo4sDpCQSeYRvNgD/yF7t0Qhl34VJvg8OGo8fBngMH8m7rap
ZdyoZcqQqRNQXRJ6wiAuSKN/QmftI1onammNOT7hwTm8ypdksJFGT/RF6YRzAUlyoqd9E2/U0HRi
3rCxV7DDl1KAtPnkxO56kB7Dso+FzotWKbJyGEw52Kb9FKeDLbzJhRAlXb4T5YzcB7nSLKEuZISL
QTekwB59S+WsNi/pFD6/4oFx/QsxExiWluNGzy8PvOq5541AKOTSLRqZ+xVh+kOMBSIAg7bDEDxF
qxj+4Xtkekl0yTUXewLqq34mxa02IsmsCWpZ0c3scOvRbp/0wKvIJeg7J1PS+Fp7dTakqfMrsl5R
dm1ZBvZ7RtuUlyJNQokgJ5Qd1DjUpXNyFM34KI2229rOvvwxTFLSjlP46HQUyi01DLECZJulk5wm
wdWYOMDYFTybg1927fEnnJHIpQEWHWz1zbZhlj51Fr6c9rk/aMCSgVD23uHPvbarRNbJrxHv0JR2
RU51ZyhQXh5uSUMjRCmh24fm/LvuMirZWo2W3w34dlOWhfUVNxaBrRVkGqZwLJXwJg79YYVidxrz
wni+r8Wf9cXNvqMzbUkbz4HEhccHsmah1G3S2GTHLLeExEF4TjWrG4hYI8KknLCK1aWbVORQdn59
ELkb5Lq/hSU/sNQkBUOn+nVtN97PeV39FcZIPWOG/mFohsWIMalvNLOCw/iOTsMfOkotD7p4F8pt
Myglxis77vqtvJlG1+JJmlyEhiSFBteJQY67XYvw3inCE/uv3ubzFJVI5GRXfbb4BhA4HLNhIoUp
n1DvweZE8IjkXDLopfWEB9jmjhXM3rk5s35389ojhikfyJNPEomMbl2n0+FXzEYYO7BwIpk6PTix
3kpXAKuuAklfyXpdO3XPgt6m5g7TtKkBE0oZE5Q9yNKr5Qvd4xQm/KVGgF9hlxUksV6geecZwddh
fypUzfC4kJr5z0ic1gGEX4lZ0PEOXWudPa2uFOkDTLiqy7fAU3/PT1/TCMfnpT3CqSaGEYz8fxit
3knUbsyLb0C8G6Gf6nFfd8vSc7DURIFlHkWR0N7T4G8ISup8qodVLr6Xgd89/OdGwpTytDejKkNQ
zDfanwnMFe6QGupy3KlT7mFt2Ji2LpOxMwpDQNmmPHfGDf3NzTPp/cbexXnQkeYBLBSnL62AAP+J
/lf1aG+P3xsQsrSR9aK5o03s5ylP5GDvkdUwN6H7poK629JkmigM8doPmXiQIIyyY8TQkLFDwgUg
toAyMWXwCVzqN6B1k9dur4vgvKGiv20VXlr6CvpOudOFHKdYTmkEMaBoWedRE7wsCEtFo8AvSdJt
aN23xyKNqZpNVi77yfK1dYXBwe2GCYyggn6OQUx5RPg+IDRLtR8nz9lSUlJZz5Y87FMU5ZGi4IJq
74shqBtIWW4CW558Y3V58rLLqhLV4LJTX6MNhtPBBKYEXzy5VRjHMF/XD6NBu3jXyUcRUdG7WZB9
9Ix2jk/ZrRozOlZhbKIYWuJhXhwSQ0lPTbJd8mPtAe5yyppZJjp4wTpHHFl7OWGQaizSOcEH0EYi
3X2q8nkwm/OqDGXDO8XGdLZoye+9HkUtOYd4T/Om51dve+c6rLvHbUJ1QfxlbSjKEfy4AU35Dgpp
A8OQTiIckpjUtLEvqtKW3iDshv9393HPK6zwmVAiqn+zltaj+BHaIB0Hzuc5UienrK4g27BMV/G2
VnscZ7QjdIHJMiiN0pFf/dlrhlzNTFFCTJpZtbU/dPBihMbfduwKfENfeoFIluc4+wFiGC0cJwe3
T6c/v/b9mqCpQXq9/F5UE5JKhzuBfZ5gEqDfgaxAjkOU2IlN1GstXAsqqxsJARx8g1hb6ODEOp6Z
0a2iAtcfEz+2b2aXDuynyNpJ05EbVEbmsXN3mq58HOIRDLeiYxrAqlMUGcZjb8+F1rMzkqfYrpYX
O7dTKDXlY/nFqxnht4ghh0mClO3WXBx4iRCo6gSZU/HyamBADQ6TqtbfkVx9LosJ2jD94sV6ZJ77
C07pP06LNu1/k8+cTFgUahRpokoJZZMiFfLx0yeE/tSjwxehL3mJVbkii2MxSLZIcHxCSewf8zzJ
gekPU9EMo27p9t7/VSkIRCKrYr4MTkwD6Avrdc2439LaiMbgyuEQd/BVoCRrbCwWQk+3vh/AR3vQ
7f1hv5aXfM/QwE5KzSXO3FMUBGYXb0fAAAKuV8p02TmnqO9uvuxJWyzw1v3MuZ+Cldmv6c60MJ8s
orS2SUqUzo91rgr82yhXsbV8fcYWzJ2cYmfnKo5x58hTVsqMAd9GiROShjS8VxQYrpzwCMhmUmdT
hzewdNA6ONL7h3Tc5kEklMNNwED1xy1+HuDjmtdpmit4SRV3itVLuAyPefVTibN0DuxZqMrIEpgM
4t4ifkrbqT24994LS5x97zZdgefhdbFwe20U7R4G0j5w5iT8/3Wuxa8bqe7/LXfvY5FxS5giR4DE
lL8bcneTSE+1YxTo1nMS3BNGuikdWMOD/lRBEpdy4JZel3qoa4S5KlQXAHq9i7WKa2kasGtdg9FB
rSxDdsGE+2n1CEotCY9Fy0dbCqPXoqYrpdmnVtVtBlMqAz3gfhjpU9uPcrCiYH9Jcg3bAEXZjTlj
s2Dri4Y8T9ipO/ysG9TOMEGjmah6zdlYE8DoIujgKjo/8PHsvweTUxE6IkfiKROkWTjVK5o6H+0u
HbpXHhIu2EJ5PKDE6aNgsKprdmA6/4noaN5LCKiZmbAYNXKr9uG02GM38ZxhMWeVAYDLlTRlPDhM
xCnxfK+aYlqzEwCKhREcAmvLfrHOfguOQnCnmXinGwS03u0W+3Ha2FXAy8YAzWdCueoJEHX68kc0
+BSZ8AzBoLvAxCkecOp6RQl46bVLOA9Edwr9qYHMk9GwnFLlkAa3BN8C1z2UarwVYtDh2LQkyRqu
nzdDwft1P632JS0blZ9M+qBxqQ+5h+7nKIFex6gA90WUO8hwfUTIqxW0a4FirTn6r7Rgz4Ypvc9x
uzb2pQHMeeFObivA2HLGywpZU20bYP5aifMukYIspczzAQd3moEQ72Ny5uNMe7UYJu0FHbXdnJeS
5OwIpvfIq1Evh4ZdGq2awEmbCG5OrCwTamoPfXchJnnPJv20oMcKuihBvHGR+4D5y33y0fb2DTMx
RGOE7nY+Ln88SWriR2IjdqbNIYAC5K1mhmG1g+YA7mgthimLZ5JJMj5lODSLMBR6rI1WLkAse5w7
7V5dyceSKXqjVG0wt4S9V8ZVUuSri9V4a1W0TKkDABRaQ9dG+ssc+G9tE2Bpj0p7gMXrW3VdJT9L
tcv70KlSazlXfJMMy+wBU30FnWsN8chc6UnAYOxks3NJ0Q0ipk+vgOaO/nzdRJhwmx4c77vjIQBW
axH+vwsf1/u10VVmjvf1m7hNDSF3wUIhIRqVdytoZat48ntWPe7sOS+gVMLKONBv8tERn2mLmnGL
TuAoxXacXrgMfYQRTDZMmgIRlVG5P4aS0jK+tsYJNhMFAzY/QJtlX0+3k0MptVzeQdY8JPFed02D
+2AsoDVSTsAllXwdIlQMQzS4QhJwmKOLhFqixrAIzrK2skjmwsuySf0c9ZMhMuYx5kWJ3NvV2Xiq
Qy/ikMuEn4gUrELH0ETALDoS8jb/PaajiIwt8SrvVTUQP4XPXKyqEms8HtPtMq2HquS4r273iyEl
DjeBUe6eN72nL0mGYNq8kHfR4VRseflIUaGiqHqGV2xT3jh5OWVF//uFiLPcBwP3IWgvmnktfDAt
TwRd5ebzNgT3e8yLNy62rY0hm8292/bghOPY2cZa7GWhQnU0uVqaWIyvw8jW9/HUVcPCrdKYG4jq
qCVebLKWxP4utYMVfZGLJ8B/ZB9ZylmDdVvmR1TUr2uuC4LwG6umELSx6Rf45qwhnikyeI9A9SVG
OkbBy5TJqDwA8DJpczbMU/aKZvYkignkJxNn6OARcxuKz8P0uOCx75+fmEQEnKeErSljyHlT8c9+
mjiyAo4fDUJ9T3nTfLR/Nt2YS2fVpH9y0H0m5apnT5k+jRmAueI64XWSxxtJ5Zo6Ub5GVNS/+2my
Ejdd7y6PTTq7GDJo+Yf5ZDkEaSGQuYgG43KwQ3MCzT79++AKz3KPvZoiocO5lSFC2ULZ703GPogR
B9GxvatHGJ81oZ3sTiK1QzwmhOhGvuUksTDAJ6BT5IdwsheFl1Fu2Xec+XxKpttDLTrq/OgcR0nJ
mGWyc0NiJJcZC0fuKcKnL1U0Aerm4XdN3JbhYCoFYMlKVA3CzJtMGrEjdSUjSMgaeijGTNtlm4DB
LlnTHjv6g4WHWgn0N5YDux33BxR413KoyH8RAWjuiS9yp15av5iKy0QIGO56+u+5Ogl9zCnYbIoW
b293LRo+le+UnG0MCuLQ/+23jOoxEpuqMZEFcQHB3/obdRIkgeyqIJ+wrjYN9CWfc6Q2iLQjPMk4
B3ceyU40BX8bim4wD/u2ozAltz1FvhBAqbzzwqiimPvUn/zlatR4L5+W8qfwoHBJdZzYktRa71H8
R4S3y/yVnoqHjA8Q0B1glMVd7vCUw3fqcR86Pn5uIdrG06UcErCHcSU1TDMkmM4AUi8Pk+zApZ6F
Y5eF4h8wgaZHhzgVQ1syY59bfcvmJRUEWvGF0FF2HZ4gsV/fd1Eee1tWmvBsNjqHh26VIfLk3klN
hXQ2SXxmaaNfv08NcNk2l8lOsA/JoTtIenI7x4i/J6lzgFhyzOGlpsPPsN4X6j1SY/RF/fARhwYl
N2OCgoEdK6j8Q0+bul7GdikdBDyJ/+o1qGPa5zviKoSZ9+OcOViaZNUws8jvvuHer0tZn4y6tJe6
H00iKnREHNOc1SP2ZIHVY5VBAZSWMA/M1r3/C2F73ALdxR53P+VcyGPjSsfDSfVYftwZkxt2VUY0
rH+GsbSPUXFCvKPShasWP+0OH7LZ4sQiVLZQc0PhGPkk5cLK/Yr2wssbwCj3+Y3bfs2CPYmUflfN
SnWhmVKiRX8zG82cKscORXmiKs3fqhqfGq4gIuUi+2e/h0S62pxcBBQyy+53Z3zSvTMHf3R/49W8
qz/zf2uEOrmf5Fs52wK0ge+/xcXpCrcu/GrXw7yBkBnDNgOfvuZhE9epQQrHGgUtT2mmhR8r04w7
xzcJd78HexhEYR6tZpzw25dx97wBWs3Yt2hVUOZJagFeB44BvqtFjT41YaaOb+cczH9En08cRgbN
5ghmxj5K7zGKVmrXjdABG8ZPLG1pA0XcQLzJiGGhCWeaOZ8ruiL9V/NR1AI7iGOTlUNgXBgOv0ev
+ig3JHPlPEPeFS6AvV6J3u0So0/ShPwMmRuqpXzndWiXIdj9IBTCOOE1+PJhh6QZQB63l1JpTpoK
YsumU70tfRTL/rlJ46bRHHEzJ+Whpi2ZM7UuPTswrVABSGY8c0hdWrDDfHidRJwVnRlqb229eHLS
kibU1zShbNZAMHsiQvkgZa5Mb3077YsLpUh0UgsQ9E2gHICdrPs2nSwVyfty8frzuS8uqrcly1F3
OLxSSQ9L9fYxkAdCbVbMIygLFOlh6QMsI6JD6e77vpj3ry/9dHDj/urCQl3VQUvLejvpMtZyZIrl
XhY01th8ldIQIQAe2aGFtiXoSQNvB+Vb7qqnwxZ8xRICDQP1R7TOlms88P0YIWLnKrzF9NJPOgwC
J+F9jH5JA4PWkKjskSN/ZX2qIewECbBV5hTyFXwk07CHnm3whlJqjECxrS+E5KtcBvDhF2sfyaT5
EptYIS3LmhvGPDcTI0rlDC304MmCk+/fzRTuLx2XTwzoc/dy/5WYcPHk0tgpTgNMpgV5k7/pts7V
zqGNlLbh8VjwmHjsw3EgUYilVZ7hixPyWY60ZlTB711Turok8OtulhDd5BH0+LzErZ/5baGv81n4
l1Co2nE7qIVJ4hOZ9gsziF2kt6Uzltqn95Bs2Ygtngx99HYkm9p+p+bjx+Vpq2R4GAwAF6zM6gvw
+nDrSCQwnn1HYInWK7Amtvk8mUUsy5VfwKwYOqoIJ/w8eAhC3cznuIqXbdW3C+iDyhHWzwB9pHRF
VjY/iSRX8DGCxbDhtn++Ya6Qwaq25giMGxet/HfKmY/PjJMExHnJ9JMz6VUfGIYWeyRgA9dSlAIA
545vz/EcvzGn0nZfw+fZ7/Oh++VJZVhkGsCSCRjYJiyVKU/zq93lJx1SOnCLmXOuaHIcbaZamC5M
Knk+0ML6pWGhcOV8BP5hI/ryCQ6Suzi0YZoVEmFs9opqQgqeBmRTp8IS2zpk8AWOSin2oat4HPqJ
DdR0dNnAOSw5uOf9yyM6Z8KfbslgnT/+AMmiVgkYD1WV86O2KAS5dxXq//yCJw/nZUYNzjO74dWg
z0uk44im05yabVCfdO7Hmtprzhl+ksQ6ReJiuxgfEmFdtDTaMkby6i6Jm3CgYKiqg+et+lotIYqO
g70P4oyyanTQaVCEDSCHzNBHbcRjiUI/Skk3T0ruoXJ1ugYhQSAygM+xZIdYuo3CEXSYE//cS6H5
Q3V2SLMWCoc2JvvZX/DKtD4llwKiDNliy7VZ5IY07fM0mhFWG5zoVj/feElLQewxNHTeXy71NJLp
0tFFLpKKmD6qhtk3U5W3bq0itdeP9Lwhb2XkUBTfWnlBRDiT3aDauyM916nqbGCh0ZoCotuqke11
afK4uEMgP8oF9TCNqRVdpcjeC6WhpykhtTXaq8H5JvC/WdFdsm07MvFXD0R0VInepIDso9CpUZfa
4aPtkgMMOEzPp4gMhbbfVdYnsvgkNWWSmi5elVzVIOK9X6ii5bbB3++EKX3n2jGa78S4vJ9EgxM8
awI+1Rh65kl6pwIzNj8isp826Qu59XvQcOG5XY8ZmSFLgGbDz71h8lUA2HKsn0bjT55CJoW5kCGi
Apa6xIrjAVhIWhR/FEY0shUOz1ebRX/1y++IKRcOBW3YUDl6A51gwP7hzGfgWJ3mqErRwI58eZrs
7ycBcsVZPll7fomEpM9YTdEwK88IstgFiaGHZOtI8zJvnzDMW68XwpxjAlD6wsrA7HiECxkbFsBe
54llKJoLTq0Muwj0cYBpp8C/AxmWTmiY3rAhXQjWcrVoCvpi6cppX12dhnXLiOh4LEbu6bQPR/te
Jk4CeJ2gz453AWOhIQKOBrTifmCK5MKBBL7HAiTq+UjqS/J/6fmxM6ZDX2Usw0zweaH4FKt1LA4r
gj/caEbe9upza4R3JvJf+67pqe7k7gyptxhjdXHtT+5JyAblw2gV9iL+O3Uedh5TsDQOkqcdwzwO
PL1Oek8k9DyOuk3tJbYxUVDSil1fq5AuWJjPGXFeLd1L4ZnnrYahZoVHUx39Nje1yzzy2vh2icNp
THpZpoh5dZ6aUxHxxxX+NRo8QtgMm/y7xo2F4JMRHYoHHxD9krVQdYZnsD84vNOiDNLrPZeQFg/X
+FImS7iEeVfjA9TvrI97WN9ev2So9wnsIUVeRpZ6cYA6I8vjZEMQ0StPCxtJiLqIwobqkCZ5Ez29
YdwQzmfVTvWGZKUJbxMLb1bLHW7mATJaFE+hAzXdmhKPIMPobPU0RmKINd3G3bkyI5nOGe4wUEoA
RmHG7HEGY6ttRa5k1GQbXk3fwQM5oRh8kJJrNHUBzvV0ZwmYhrtCw6UfrOS1YnofaYUvyS3CSoz6
AZdn0RPKXZO9ECWG/CldBixkeqyCu05Whw==
`protect end_protected
